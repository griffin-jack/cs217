
//------> ./PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ./PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   code@rice-03
//  Generated date: Wed Jan 14 11:37:27 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_core
// ------------------------------------------------------------------


module PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_core
    (
  this_vld, this_rdy, this_dat, data_data_rsc_z, data_addr_rsc_z, data_rw_rsc_z,
      return_rsc_z, ccs_ccore_start_rsc_dat, ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  reg this_rdy;
  input [96:0] this_dat;
  output [63:0] data_data_rsc_z;
  output [23:0] data_addr_rsc_z;
  output data_rw_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations
  wire [63:0] nl_data_data_rsci_d;
  assign nl_data_data_rsci_d = this_dat[63:0];
  wire [23:0] nl_data_addr_rsci_d;
  assign nl_data_addr_rsci_d = this_dat[87:64];
  wire  nl_data_rw_rsci_d;
  assign nl_data_rw_rsci_d = this_dat[96];
  PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd1),
  .width(32'sd64)) data_data_rsci (
      .d(nl_data_data_rsci_d[63:0]),
      .z(data_data_rsc_z)
    );
  PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd2),
  .width(32'sd24)) data_addr_rsci (
      .d(nl_data_addr_rsci_d[23:0]),
      .z(data_addr_rsc_z)
    );
  PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd4),
  .width(32'sd1)) data_rw_rsci (
      .d(nl_data_rw_rsci_d),
      .z(data_rw_rsc_z)
    );
  PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd6),
  .width(32'sd1)) return_rsci (
      .d(this_vld),
      .z(return_rsc_z)
    );
  PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1
      #(.rscid(32'sd153),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_rdy <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB
// ------------------------------------------------------------------


module PECore_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB
    (
  this_vld, this_rdy, this_dat, data_data_rsc_z, data_addr_rsc_z, data_rw_rsc_z,
      return_rsc_z, ccs_ccore_start_rsc_dat, ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  input [96:0] this_dat;
  output [63:0] data_data_rsc_z;
  output [23:0] data_addr_rsc_z;
  output data_rw_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  PECore_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_core
      Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .data_data_rsc_z(data_data_rsc_z),
      .data_addr_rsc_z(data_addr_rsc_z),
      .data_rw_rsc_z(data_rw_rsc_z),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ./PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   code@rice-03
//  Generated date: Wed Jan 14 11:37:22 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_core
// ------------------------------------------------------------------


module PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_core
    (
  this_vld, this_rdy, this_dat, data_data_data_rsc_z, data_logical_addr_rsc_z, return_rsc_z,
      ccs_ccore_start_rsc_dat, ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  reg this_rdy;
  input [73:0] this_dat;
  output [63:0] data_data_data_rsc_z;
  output [7:0] data_logical_addr_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations
  wire [63:0] nl_data_data_data_rsci_d;
  assign nl_data_data_data_rsci_d = this_dat[63:0];
  wire [7:0] nl_data_logical_addr_rsci_d;
  assign nl_data_logical_addr_rsci_d = this_dat[73:66];
  PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd7),
  .width(32'sd64)) data_data_data_rsci (
      .d(nl_data_data_data_rsci_d[63:0]),
      .z(data_data_data_rsc_z)
    );
  PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd9),
  .width(32'sd8)) data_logical_addr_rsci (
      .d(nl_data_logical_addr_rsci_d[7:0]),
      .z(data_logical_addr_rsc_z)
    );
  PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd11),
  .width(32'sd1)) return_rsci (
      .d(this_vld),
      .z(return_rsc_z)
    );
  PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1
      #(.rscid(32'sd152),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_rdy <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB
// ------------------------------------------------------------------


module PECore_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB (
  this_vld, this_rdy, this_dat, data_data_data_rsc_z, data_logical_addr_rsc_z, return_rsc_z,
      ccs_ccore_start_rsc_dat, ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  input [73:0] this_dat;
  output [63:0] data_data_data_rsc_z;
  output [7:0] data_logical_addr_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  PECore_Connections_InBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_core
      Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .data_data_data_rsc_z(data_data_data_rsc_z),
      .data_logical_addr_rsc_z(data_logical_addr_rsc_z),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   code@rice-03
//  Generated date: Wed Jan 14 11:37:19 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_spec_ActVectorType_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_spec_ActVectorType_Connections_SYN_PORT_Push_core
    (
  this_vld, this_rdy, this_dat, m_data_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  reg this_vld;
  input this_rdy;
  output [255:0] this_dat;
  reg [255:0] this_dat;
  input [255:0] m_data_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire [255:0] m_data_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  wire and_dcpl;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_4_cse;
  wire this_vld_mx0c1;


  // Interconnect Declarations for Component Instantiations
  wire  nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd13),
  .width(32'sd256)) m_data_rsci (
      .dat(m_data_rsc_dat),
      .idat(m_data_rsci_idat)
    );
  PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd151),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1
      #(.rscid(32'sd155)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld)
    );
  assign or_4_cse = ccs_ccore_start_rsci_idat | and_dcpl;
  assign and_dcpl = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_rdy);
  assign this_vld_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_vld <= 1'b0;
    end
    else if ( or_4_cse | this_vld_mx0c1 ) begin
      this_vld <= ~ this_vld_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_dat <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~(and_dcpl | (~ ccs_ccore_start_rsci_idat)) ) begin
      this_dat <= m_data_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_4_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_spec_ActVectorType_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module PECore_Connections_OutBlocking_spec_ActVectorType_Connections_SYN_PORT_Push (
  this_vld, this_rdy, this_dat, m_data_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  input this_rdy;
  output [255:0] this_dat;
  input [255:0] m_data_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  PECore_Connections_OutBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_spec_ActVectorType_Connections_SYN_PORT_Push_core
      Connections_OutBlocking_spec_ActVectorType_Connections_SYN_PORT_Push_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .m_data_rsc_dat(m_data_rsc_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ./PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   code@rice-03
//  Generated date: Wed Jan 14 11:37:16 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_core
// ------------------------------------------------------------------


module PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_core
    (
  this_vld, this_rdy, this_dat, data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  reg this_rdy;
  input this_dat;
  output data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations
  PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd15),
  .width(32'sd1)) data_rsci (
      .d(this_dat),
      .z(data_rsc_z)
    );
  PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd17),
  .width(32'sd1)) return_rsci (
      .d(this_vld),
      .z(return_rsc_z)
    );
  PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1
      #(.rscid(32'sd150),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_rdy <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_bool_Connections_SYN_PORT_PopNB
// ------------------------------------------------------------------


module PECore_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB (
  this_vld, this_rdy, this_dat, data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  input this_dat;
  output data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  PECore_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_core
      Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_core_inst (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .data_rsc_z(data_rsc_z),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   code@rice-03
//  Generated date: Wed Jan 14 11:37:24 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push_core
    (
  this_vld, this_rdy, this_dat, m_data_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  reg this_vld;
  input this_rdy;
  output [63:0] this_dat;
  reg [63:0] this_dat;
  input [63:0] m_data_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire [63:0] m_data_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  wire and_dcpl;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_4_cse;
  wire this_vld_mx0c1;


  // Interconnect Declarations for Component Instantiations
  wire  nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd18),
  .width(32'sd64)) m_data_rsci (
      .dat(m_data_rsc_dat),
      .idat(m_data_rsci_idat)
    );
  PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd149),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1
      #(.rscid(32'sd154)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld)
    );
  assign or_4_cse = ccs_ccore_start_rsci_idat | and_dcpl;
  assign and_dcpl = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_rdy);
  assign this_vld_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_vld <= 1'b0;
    end
    else if ( or_4_cse | this_vld_mx0c1 ) begin
      this_vld <= ~ this_vld_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_dat <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~(and_dcpl | (~ ccs_ccore_start_rsci_idat)) ) begin
      this_dat <= m_data_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_4_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module PECore_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push
    (
  this_vld, this_rdy, this_dat, m_data_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  input this_rdy;
  output [63:0] this_dat;
  input [63:0] m_data_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  PECore_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push_core
      Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .m_data_rsc_dat(m_data_rsc_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./PECore_mgc_muladd1_beh.v 
//muladd1
module PECore_mgc_muladd1(a,b,c,cst,d,z);
  // operation is z = a * (b + d) + c + cst
  parameter width_a = 0;
  parameter signd_a = 0;
  parameter width_b = 0;
  parameter signd_b = 0;
  parameter width_c = 0;
  parameter signd_c = 0;
  parameter width_cst = 0;
  parameter signd_cst = 0;
  parameter width_d = 0;
  parameter signd_d = 0;
  parameter width_z = 0;
  parameter add_axb = 1;
  parameter add_c = 1;
  parameter add_d = 1;
  parameter use_const = 1;

  function integer is_square_op;
    input integer alen;
  begin
    if (alen > 1) is_square_op = 0;
    else       is_square_op = 1;
  end endfunction

  input  [width_a-1:0] a;
  input  [width_b-1:0] b;
  input  [width_c-1:0] c;
  input  [width_cst-1:0] cst; // spyglass disable SYNTH_5121,W240
  input  [width_d-1:0] d;
  output [width_z-1:0] z;

  reg [width_a-signd_a:0] aa;
  reg [width_b-signd_b:0] bb;
  reg [width_c-signd_c:0] cc;
  reg [width_d-signd_d:0] dd;
  reg [width_cst-signd_cst:0] cstin;

  localparam width_bd = (width_d) ? 1+ ((width_b-signd_b>width_d-signd_d) ? width_b - signd_b
                                                                          : width_d - signd_d)
                                  : width_b - signd_b;
  localparam is_square = is_square_op(width_a);
  localparam axb_len = (is_square)?width_bd+1+width_bd+1:width_a-signd_a+1+width_bd+1;

  reg [width_bd:0] bd;
  reg [axb_len-1:0] axb;



  // make all inputs signed
  always @(*) aa = signd_a ? a : {1'b0, a};
  always @(*) bb = signd_b ? b : {1'b0, b};
  generate if (width_c != 0) begin
    always @(*) cc = signd_c ? c : {1'b0, c};
  end endgenerate

  generate if (width_d) begin
    if ( !is_square) begin
      (* keep ="true" *) reg [width_d-signd_d:0] d_keep;
      always @(*) d_keep = signd_d ? d : {1'b0, d};
      always @(*) dd = d_keep;
    end else begin
      always @(*) dd = signd_d ? d : {1'b0, d};
    end
  end endgenerate

  always @(*) cstin = signd_cst ? cst : {1'b0, cst};

  // perform pre-adder
  generate
    if (width_d != 0) begin
      if (add_d) begin always @(*)  bd = $signed(bb) + $signed(dd); end
      else       begin always @(*)  bd = $signed(bb) - $signed(dd); end
    end else     begin always @(*)  bd = $signed(bb); end
  endgenerate

  generate
    if (is_square)
      always @(*) axb = $signed(bd) * $signed(bd);
    else
      always @(*) axb = $signed(aa) * $signed(bd);
  endgenerate

  // perform muladd1
  wire [width_z-1:0]  zz;

  generate
    if (use_const) begin
      if ( add_axb &&  add_c && width_c) begin assign zz = $signed(axb) + $signed(cc) + $signed(cstin); end else
      if ( add_axb && !add_c && width_c) begin assign zz = $signed(axb) - $signed(cc) + $signed(cstin); end else
      if (!add_axb &&  add_c && width_c) begin assign zz = $signed(cc) - $signed(axb) + $signed(cstin); end else
      if (!add_axb && !add_c && width_c) begin assign zz = $signed(cstin) - $signed(axb) - $signed(cc); end else
      if ( add_axb )                     begin assign zz = $signed(axb) + $signed(cstin); end else
                                         begin assign zz = $signed(cstin) - $signed(axb); end
    end  else begin
      if ( add_axb &&  add_c && width_c) begin assign zz = $signed(axb) + $signed(cc); end else
      if ( add_axb && !add_c && width_c) begin assign zz = $signed(axb) - $signed(cc); end else
      if (!add_axb &&  add_c && width_c) begin assign zz = $signed(cc) - $signed(axb); end else
      if (!add_axb && !add_c && width_c) begin assign zz = -$signed(axb) - $signed(cc); end else
      if ( add_axb )                     begin assign zz = $signed(axb); end else
                                         begin assign zz = -$signed(axb); end
    end
  endgenerate

  // adjust output
  assign z = zz;
endmodule // mgc_muladd1

//------> ./PECore_mgc_shift_l_beh_v5.v 
module PECore_mgc_shift_l_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> ./PECore_mgc_mulacc_pipe_beh.v 
//mulacc
module PECore_mgc_mulacc_pipe(a,b,c,d,load,datavalid,clk,en,a_rst,s_rst,z);

  parameter width_a = 0;
  parameter signd_a = 0;
  parameter width_b = 0;
  parameter signd_b = 0;
  parameter width_c = 0;
  parameter signd_c = 0;
  parameter width_d = 0;
  parameter signd_d = 0;
  parameter width_z = 0;
  parameter add_d = 1;
  parameter is_square = 0;
  parameter      clock_edge =  1'b0;  // clock polarity (1=posedge, 0=negedge)
  parameter   enable_active =  1'b0;  // enable polarity (1=posedge, 0=negedge)
  parameter    a_rst_active =  1'b1;  // unused
  parameter    s_rst_active =  1'b1;  // unused
  parameter integer  stages = 32'd2;  // number of output registers + 1 (careful!)
  parameter integer n_inreg = 32'd0;  // number of input registers

  function integer max_len;
    input integer a, b;
  begin
    if (a > b) max_len = a;
    else       max_len = b;
  end endfunction

  function integer min_len;
    input integer a, b;
  begin
    if (a > b) min_len = b;
    else       min_len = a;
  end endfunction

  localparam axb_stages = (stages>2) ? 1 : 0;

  localparam preadd_stages = (n_inreg>1) ? 1 : 0;
  localparam bb_stages = n_inreg - preadd_stages;
  localparam cc_stages = n_inreg + axb_stages;
  localparam cc_len = min_len(width_c-signd_c+1, width_z);

  localparam zz_stages = stages - axb_stages;

  localparam width_bd = (width_d>0) ? (1+ ((width_b-signd_b>width_d-signd_d) ? width_b - signd_b : width_d - signd_d)) : width_b - signd_b;
  localparam axb_len = (is_square)?width_bd+1+width_bd+1:width_a-signd_a+1+width_bd+1;

  localparam zz_len = max_len(axb_len, max_len(cc_len, width_z));

  reg [width_bd:0] bd [preadd_stages:0];

  input  [width_a-1:0] a;
  input  [width_b-1:0] b;
  input  [width_c-1:0] c;
  input  [width_d-1:0] d; // spyglass disable SYNTH_5121,W240
  input                load;
  input                datavalid;

  input                clk;    // clock
  input                en;     // enable
  input                a_rst;  // spyglass disable SYNTH_5121,W240
  input                s_rst;  // spyglass disable SYNTH_5121,W240

  output [width_z-1:0] z;

  reg [width_a-signd_a:0] aa [n_inreg:0];
  reg [width_b-signd_b:0] bb [n_inreg:0];
  reg [width_c-signd_c:0] cc [cc_stages:0];
  reg [width_d-signd_d:0] dd [bb_stages:0];
  reg                     accum [cc_stages:0];
  reg                     vl [cc_stages:0];

  genvar i;

  // make all inputs signed
  always @(*) aa[n_inreg]   = signd_a ? a : {1'b0, a};
  always @(*) bb[bb_stages]   = signd_b ? b : {1'b0, b};
  generate if (width_d>0) begin
    always @(*) dd[bb_stages]   = signd_d ? d : {1'b0, d};
  end endgenerate
  always @(*) cc[cc_stages] = (signd_c | width_c >= width_z) ? c : {1'b0, c};
  always @(*) accum[cc_stages] = !load;
  always @(*) vl[cc_stages] = datavalid;

  // input registers
  generate if (n_inreg>0) begin
  for(i = n_inreg-1; i >= 0; i=i-1) begin:ab_pipe
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) aa[i] <= aa[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) aa[i] <= aa[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate
  generate if (bb_stages>0) begin
  for(i = bb_stages-1; i >= 0; i=i-1) begin:in_pipe_bd
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) bb[i] <= bb[i+1];
      if (width_d>0) begin  always @(posedge(clk)) if (en == enable_active) dd[i] <= dd[i+1]; end //spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) bb[i] <= bb[i+1];
      if (width_d>0) begin  always @(negedge(clk)) if (en == enable_active) dd[i] <= dd[i+1]; end //spyglass disable FlopEConst
    end
  end end endgenerate
  generate if (cc_stages>0) begin
  for(i = cc_stages-1; i >= 0; i=i-1) begin:c_pipe
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) cc[i] <= cc[i+1];//spyglass disable FlopEConst
      always @(posedge(clk)) if (en == enable_active) accum[i] <= accum[i+1];//spyglass disable FlopEConst
      always @(posedge(clk)) if (en == enable_active) vl[i] <= vl[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) cc[i] <= cc[i+1];//spyglass disable FlopEConst
      always @(negedge(clk)) if (en == enable_active) accum[i] <= accum[i+1];//spyglass disable FlopEConst
      always @(negedge(clk)) if (en == enable_active) vl[i] <= vl[i+1];
    end
  end end endgenerate

  // perform pre-adder
  generate
    if (width_d>0) begin
      if (add_d != 0) begin always @(*)  bd[preadd_stages] = $signed(bb[0]) + $signed(dd[0]); end
      else            begin always @(*)  bd[preadd_stages] = $signed(bb[0]) - $signed(dd[0]); end
    end else          begin always @(*)  bd[preadd_stages] = $signed(bb[0]); end
  endgenerate
  generate if (preadd_stages>0) begin
  for(i = preadd_stages-1; i >= 0; i=i-1) begin:preadd_pipe
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) bd[i] <= bd[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) bd[i] <= bd[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate

  // perform muladd1
  reg [zz_len-1:0]  zz[zz_stages-1:0];
  wire [zz_len-1:0] z_or_c;
  reg [axb_len-1:0] axb[axb_stages:0];
  generate
    if (is_square>0)
      always @(*) axb[axb_stages] = $signed(bd[0]) * $signed(bd[0]);
    else
      always @(*) axb[axb_stages] = $signed(aa[0]) * $signed(bd[0]);
  endgenerate

  generate if (axb_stages>0) begin
  for(i = axb_stages-1; i >= 0; i=i-1) begin:axb_pipe
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) axb[i] <= axb[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) axb[i] <= axb[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate

  assign z_or_c = accum[0] ? $signed(zz[zz_stages-2]): $signed(cc[0]);
  always @(*) zz[zz_stages-1] = $signed(axb[0]) + $signed(z_or_c);

  // Output registers:
  generate for(i = zz_stages-2; i >= 0; i=i-1) begin:out_pipe
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active && (vl[0] || i != zz_stages-2)) zz[i] <= zz[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active && (vl[0] || i != zz_stages-2)) zz[i] <= zz[i+1];//spyglass disable FlopEConst
    end
  end endgenerate

  // adjust output
  // use a tmp var to satisfy W164a lint violations
  wire [width_z-1:0] z_out_tmp;
  assign z_out_tmp = zz[0][width_z-1:0];
  assign z = z_out_tmp;

endmodule // mgc_mulacc_pipe

//------> ./PECore_mgc_mul4acc_pipe_beh.v 
//mulacc
module PECore_mgc_mul4acc_pipe(a0,a1,b0,b1,c0,c1,d0,d1,e,load,datavalid,clk,en,a_rst,s_rst,z);

  parameter width_a0 = 0;
  parameter signd_a0 = 0;
  parameter width_a1 = 0;
  parameter signd_a1 = 0;
  parameter width_b0 = 0;
  parameter signd_b0 = 0;
  parameter width_b1 = 0;
  parameter signd_b1 = 0;
  parameter width_c0 = 0;
  parameter signd_c0 = 0;
  parameter width_c1 = 0;
  parameter signd_c1 = 0;
  parameter width_d0 = 0;
  parameter signd_d0 = 0;
  parameter width_d1 = 0;
  parameter signd_d1 = 0;
  parameter width_e  = 0;
  parameter signd_e  = 0;
  parameter width_z = 0;
  parameter add_a    = 1;
  parameter add_b    = 1;
  parameter add_c    = 1;
  parameter min_fb_size    = -1;

  parameter      clock_edge =  1'b0;  // clock polarity (1=posedge, 0=negedge)
  parameter   enable_active =  1'b0;  // enable polarity (1=posedge, 0=negedge)
  parameter    a_rst_active =  1'b1;  // unused
  parameter    s_rst_active =  1'b1;  // unused
  parameter integer  stages = 32'd2;  // number of output registers + 1 (careful!)
  parameter integer n_inreg = 32'd0;  // number of input registers

  function integer max_len;
    input integer a, b;
  begin
    if (a > b) max_len = a;
    else       max_len = b;
  end endfunction

  function integer min_len;
    input integer a, b;
  begin
    if (a > b) min_len = b;
    else       min_len = a;
  end endfunction

  localparam nb_prod_reg = 0;
  localparam nb_in_reg = n_inreg - nb_prod_reg;
  localparam nb_sop_reg = (stages>2)?1:0;
  localparam out_stages = stages - nb_sop_reg;

  localparam ee_len = min_len(width_e-signd_e+1, width_z);
  localparam zz_len = (min_fb_size>width_z)?min_fb_size:width_z;
  localparam proda_len = width_a0-signd_a0+width_a1-signd_a1+2;
  localparam prodb_len = width_b0-signd_b0+width_b1-signd_b1+2;
  localparam prodc_len = width_c0-signd_c0+width_c1-signd_c1+2;
  localparam prodd_len = width_d0-signd_d0+width_d1-signd_d1+2;
  localparam sop_len = 2 + max_len(proda_len,max_len(prodb_len,max_len(prodc_len,prodd_len)));

  localparam proda_pol  = (add_a>0)?1:-1;
  localparam prodb_pol  = (add_b>0)?1:-1;
  localparam prodc_pol  = (add_c>0)?1:-1;
  localparam prodd_pol  = 1;

  input  [width_a0-1:0] a0;
  input  [width_a1-1:0] a1;
  input  [width_b0-1:0] b0;
  input  [width_b1-1:0] b1;
  input  [width_c0-1:0] c0;
  input  [width_c1-1:0] c1;
  input  [width_d0-1:0] d0; // spyglass disable SYNTH_5121,W240
  input  [width_d1-1:0] d1; // spyglass disable SYNTH_5121,W240
  input  [width_e-1:0]  e;
  input                load;
  input                datavalid;

  input                clk;    // clock
  input                en;     // enable
  input                a_rst;  // spyglass disable SYNTH_5121,W240
  input                s_rst;  // spyglass disable SYNTH_5121,W240

  output [width_z-1:0] z;



  reg [width_a0-signd_a0:0] aa0 [nb_in_reg:0];
  reg [width_b0-signd_b0:0] bb0 [nb_in_reg:0];
  reg [width_c0-signd_c0:0] cc0 [nb_in_reg:0];
  reg [width_d0-signd_d0:0] dd0 [nb_in_reg:0];
  reg [width_a1-signd_a1:0] aa1 [nb_in_reg:0];
  reg [width_b1-signd_b1:0] bb1 [nb_in_reg:0];
  reg [width_c1-signd_c1:0] cc1 [nb_in_reg:0];
  reg [width_d1-signd_d1:0] dd1 [nb_in_reg:0];
  reg [sop_len-1:0] sop [nb_sop_reg:0];

  reg [width_e-signd_e:0] ee [n_inreg:0];
  reg                     accum [n_inreg:0];
  reg                     vl [n_inreg:0];

  genvar i;

  // make all inputs signed
  always @(*) aa0[nb_in_reg] = signd_a0 ? a0 : {1'b0, a0};
  always @(*) bb0[nb_in_reg] = signd_b0 ? b0 : {1'b0, b0};
  always @(*) cc0[nb_in_reg] = signd_c0 ? c0 : {1'b0, c0};
  generate if (width_d1>0 && width_d0>0) begin
    always @(*) dd0[nb_in_reg] = signd_d0 ? d0 : {1'b0, d0};
  end endgenerate
  always @(*) aa1[nb_in_reg] = signd_a1 ? a1 : {1'b0, a1};
  always @(*) bb1[nb_in_reg] = signd_b1 ? b1 : {1'b0, b1};
  always @(*) cc1[nb_in_reg] = signd_c1 ? c1 : {1'b0, c1};
  generate if (width_d1>0 && width_d0>0) begin
    always @(*) dd1[nb_in_reg] = signd_d1 ? d1 : {1'b0, d1};
  end endgenerate
  always @(*) ee[nb_in_reg] = signd_e ? e : {1'b0, e};
  always @(*) accum[n_inreg] = !load;
  always @(*) vl[n_inreg] = datavalid;

  // input registers
  generate if (n_inreg>0) begin
  for(i = n_inreg-1; i >= 0; i=i-1) begin:in_pipe_prod
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) aa0[i] <= aa0[i+1];//spyglass disable FlopEConst
      always @(posedge(clk)) if (en == enable_active) aa1[i] <= aa1[i+1];//spyglass disable FlopEConst
      always @(posedge(clk)) if (en == enable_active) bb0[i] <= bb0[i+1];//spyglass disable FlopEConst
      always @(posedge(clk)) if (en == enable_active) bb1[i] <= bb1[i+1];//spyglass disable FlopEConst
      always @(posedge(clk)) if (en == enable_active) cc0[i] <= cc0[i+1];//spyglass disable FlopEConst
      always @(posedge(clk)) if (en == enable_active) cc1[i] <= cc1[i+1];//spyglass disable FlopEConst
      if (width_d0>0 && width_d1>0) begin
        always @(posedge(clk)) if (en == enable_active) dd0[i] <= dd0[i+1];//spyglass disable FlopEConst
        always @(posedge(clk)) if (en == enable_active) dd1[i] <= dd1[i+1];//spyglass disable FlopEConst
      end
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) aa0[i] <= aa0[i+1];//spyglass disable FlopEConst
      always @(negedge(clk)) if (en == enable_active) aa1[i] <= aa1[i+1];//spyglass disable FlopEConst
      always @(negedge(clk)) if (en == enable_active) bb0[i] <= bb0[i+1];//spyglass disable FlopEConst
      always @(negedge(clk)) if (en == enable_active) bb1[i] <= bb1[i+1];//spyglass disable FlopEConst
      always @(negedge(clk)) if (en == enable_active) cc0[i] <= cc0[i+1];//spyglass disable FlopEConst
      always @(negedge(clk)) if (en == enable_active) cc1[i] <= cc1[i+1];//spyglass disable FlopEConst
      if (width_d0>0 && width_d1>0) begin
        always @(negedge(clk)) if (en == enable_active) dd0[i] <= dd0[i+1];//spyglass disable FlopEConst
        always @(negedge(clk)) if (en == enable_active) dd1[i] <= dd1[i+1];//spyglass disable FlopEConst
      end
    end
  end end endgenerate

  generate if (n_inreg>0) begin
  for(i = n_inreg-1; i >= 0; i=i-1) begin:in_pipe
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) accum[i] <= accum[i+1];//spyglass disable FlopEConst
      always @(posedge(clk)) if (en == enable_active) vl[i] <= vl[i+1];//spyglass disable FlopEConst
      always @(posedge(clk)) if (en == enable_active) ee[i] <= ee[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) accum[i] <= accum[i+1];//spyglass disable FlopEConst
      always @(negedge(clk)) if (en == enable_active) vl[i] <= vl[i+1];//spyglass disable FlopEConst
      always @(negedge(clk)) if (en == enable_active) ee[i] <= ee[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate

  // perform products
  reg  [width_a0-signd_a0+1+width_a1-signd_a1+1-1:0] xa[nb_prod_reg:0];
  reg  [width_b0-signd_b0+1+width_b1-signd_b1+1-1:0] xb[nb_prod_reg:0];
  reg  [width_c0-signd_c0+1+width_c1-signd_c1+1-1:0] xc[nb_prod_reg:0];
  reg  [width_d0-signd_d0+1+width_d1-signd_d1+1-1:0] xd[nb_prod_reg:0];
  always @(*) xa[nb_prod_reg] = $signed(aa0[0]) * $signed(aa1[0]);
  always @(*) xb[nb_prod_reg] = $signed(bb0[0]) * $signed(bb1[0]);
  always @(*) xc[nb_prod_reg] = $signed(cc0[0]) * $signed(cc1[0]);
  generate if (nb_prod_reg>0) begin
  for(i = nb_prod_reg-1; i >= 0; i=i-1) begin:prod_pipe1
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) xa[i] <= xa[i+1];//spyglass disable FlopEConst
      always @(posedge(clk)) if (en == enable_active) xb[i] <= xb[i+1];//spyglass disable FlopEConst
      always @(posedge(clk)) if (en == enable_active) xc[i] <= xc[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) xa[i] <= xa[i+1];//spyglass disable FlopEConst
      always @(negedge(clk)) if (en == enable_active) xb[i] <= xb[i+1];//spyglass disable FlopEConst
      always @(negedge(clk)) if (en == enable_active) xc[i] <= xc[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate

  generate if (width_d0>0 && width_d1>0) begin:prod_pipe2
    always @(*) xd[nb_prod_reg] = $signed(dd0[0]) * $signed(dd1[0]);
    if (nb_prod_reg>0) begin
    for(i = nb_prod_reg-1; i >= 0; i=i-1) begin:prod_pipe3
      if (clock_edge == 1'b1) begin:pos
        always @(posedge(clk)) if (en == enable_active) xd[i] <= xd[i+1];//spyglass disable FlopEConst
      end else begin:neg
        always @(negedge(clk)) if (en == enable_active) xd[i] <= xd[i+1];//spyglass disable FlopEConst
      end
    end end
  end endgenerate


  generate
    if ( width_d0>0 && width_d1>0)       always @(*) sop[nb_sop_reg] = proda_pol*$signed(xa[0]) + prodb_pol*$signed(xb[0]) + prodc_pol*$signed(xc[0]) + prodd_pol*$signed(xd[0]);
    if ( width_d0==0 && width_d1==0) begin
      // Not supported by Vivado2020.2 : always @(*) sop[sumofprod_stages] = proda_pol*$signed(xa[0]) + prodb_pol*$signed(xb[0]) + prodc_pol*$signed(c1xc2[0]);
      if ( add_a==1 && add_b==1 && add_c==1) always @(*) sop[nb_sop_reg] = $signed(xa[0]) + $signed(xb[0]) + $signed(xc[0]);
      if ( add_a==1 && add_b==1 && add_c==0) always @(*) sop[nb_sop_reg] = $signed(xa[0]) + $signed(xb[0]) - $signed(xc[0]);
      if ( add_a==1 && add_b==0 && add_c==1) always @(*) sop[nb_sop_reg] = $signed(xa[0]) - $signed(xb[0]) + $signed(xc[0]);
      if ( add_a==1 && add_b==0 && add_c==0) always @(*) sop[nb_sop_reg] = $signed(xa[0]) - $signed(xb[0]) - $signed(xc[0]);
      if ( add_a==0 && add_b==1 && add_c==1) always @(*) sop[nb_sop_reg] = -$signed(xa[0]) + $signed(xb[0]) + $signed(xc[0]);
      if ( add_a==0 && add_b==1 && add_c==0) always @(*) sop[nb_sop_reg] = -$signed(xa[0]) + $signed(xb[0]) - $signed(xc[0]);
      if ( add_a==0 && add_b==0 && add_c==1) always @(*) sop[nb_sop_reg] = -$signed(xa[0]) - $signed(xb[0]) + $signed(xc[0]);
      if ( add_a==0 && add_b==0 && add_c==0) always @(*) sop[nb_sop_reg] = -$signed(xa[0]) - $signed(xb[0]) - $signed(xc[0]);
    end
  endgenerate
  generate if (nb_sop_reg>0) begin
  for(i = nb_sop_reg-1; i >= 0; i=i-1) begin:sop_pipe1
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active) sop[i] <= sop[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active) sop[i] <= sop[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate

  reg  [zz_len-1:0]  zz[out_stages-1:0];
  wire [zz_len-1:0]  z_or_e;
  assign z_or_e = accum[0] ? $signed(zz[out_stages-2]) : $signed(ee[0]);
  always @(*) zz[out_stages-1] = $signed(z_or_e) + $signed(sop[0]);

  // Output registers:
  generate if (out_stages>1) begin
  for(i = out_stages-2; i >= 0; i=i-1) begin:out_pipe
    if (clock_edge == 1'b1) begin:pos
      always @(posedge(clk)) if (en == enable_active && (vl[0] || i != out_stages-2)) zz[i] <= zz[i+1];//spyglass disable FlopEConst
    end else begin:neg
      always @(negedge(clk)) if (en == enable_active && (vl[0] || i != out_stages-2)) zz[i] <= zz[i+1];//spyglass disable FlopEConst
    end
  end end endgenerate

  // adjust output
  assign z = zz[0];

endmodule // mgc_mul4acc_pipe

//------> /cad/mentor/2024.2_1/Mgc_home/pkgs/ccs_xilinx/hdl/BLOCK_1R1W_RBW.v 
// Memory Type:            BLOCK
// Operating Mode:         Simple Dual Port (2-Port)
// Clock Mode:             Single Clock
// 
// RTL Code RW Resolution: RBW
// Catapult RW Resolution: RBW
// 
// HDL Work Library:       Xilinx_RAMS_lib
// Component Name:         BLOCK_1R1W_RBW
// Latency = 1:            RAM with no registers on inputs or outputs
//         = 2:            adds embedded register on RAM output
//         = 3:            adds fabric registers to non-clock input RAM pins
//         = 4:            adds fabric register to output (driven by embedded register from latency=2)
// suppress_sim_read_addr_range_errs:  0 - report errors  1 - suppress errors

module BLOCK_1R1W_RBW #(
  parameter addr_width = 8 ,
  parameter data_width = 7 ,
  parameter depth = 256 ,
  parameter latency = 1 ,
  parameter suppress_sim_read_addr_range_errs = 1 
  
)( clk,clken,d,q,radr,re,wadr,we);

  input  clk;
  input  clken;
  input [data_width-1:0] d;
  output [data_width-1:0] q;
  input [addr_width-1:0] radr;
  input  re;
  input [addr_width-1:0] wadr;
  input  we;
  
  (* ram_style = "block" , syn_ramstyle = "block" *)
  reg [data_width-1:0] mem [depth-1:0];
  integer j;
  initial for (j = 0; j < depth; j = j + 1) mem[j] = 0;
  
  reg [data_width-1:0] ramq;
  
  // Port Map
  // readA :: CLOCK clk ENABLE clken DATA_OUT q ADDRESS radr READ_ENABLE re
  // writeA :: CLOCK clk ENABLE clken DATA_IN d ADDRESS wadr WRITE_ENABLE we

  generate
    // Register all non-clock inputs (latency < 3)
    if (latency > 2 ) begin
      reg [addr_width-1:0] radr_reg;
      reg re_reg;
      reg [data_width-1:0] d_reg;
      reg [addr_width-1:0] wadr_reg;
      reg we_reg;
      
      always @(posedge clk) begin
        if (clken) begin
          radr_reg <= radr;
          re_reg <= re;
        end
      end
      always @(posedge clk) begin
        if (clken) begin
          d_reg <= d;
          wadr_reg <= wadr;
          we_reg <= we;
        end
      end
      
    // Access memory with registered inputs
      always @(posedge clk) begin
        if (clken) begin
            ramq <= mem[radr_reg];
            if (we_reg) begin
              mem[wadr_reg] <= d_reg;
            end
        end
      end
      
    end // END register inputs

    else begin
    // latency = 1||2: Access memory with non-registered inputs
      always @(posedge clk) begin
        if (clken) begin
            ramq <= mem[radr];
            if (we) begin
              mem[wadr] <= d;
            end
        end
      end
      
    end
  endgenerate //END input port generate 

  generate
    // latency=1: sequential RAM outputs drive module outputs
    if (latency == 1) begin
      assign q = ramq;
      
    end

    else if (latency == 2 || latency == 3) begin
    // latency=2: sequential (RAM output => tmp register => module output)
      reg [data_width-1:0] tmpq;
      
      always @(posedge clk) begin
        if (clken) begin
          tmpq <= ramq;
        end
      end
      
      assign q = tmpq;
      
    end
    else if (latency == 4) begin
    // latency=4: (RAM => tmp1 register => tmp2 fabric register => module output)
      reg [data_width-1:0] tmp1q;
      
      reg [data_width-1:0] tmp2q;
      
      always @(posedge clk) begin
        if (clken) begin
          tmp1q <= ramq;
        end
      end
      
      always @(posedge clk) begin
        if (clken) begin
          tmp2q <= tmp1q;
        end
      end
      
      assign q = tmp2q;
      
    end
    else begin
      //Add error check if latency > 4 or add N-pipeline regs
    end
  endgenerate //END output port generate

endmodule

//------> ./PECore.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
// 
//  Generated by:   code@iron-06
//  Generated date: Thu Jan 15 13:41:12 2026
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_146_12_64_4096_1_4096_64_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_146_12_64_4096_1_4096_64_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [63:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [63:0] d;
  output [11:0] wadr;
  input clken_d;
  input [63:0] d_d;
  output [63:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_145_12_64_4096_1_4096_64_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_145_12_64_4096_1_4096_64_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [63:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [63:0] d;
  output [11:0] wadr;
  input clken_d;
  input [63:0] d_d;
  output [63:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_144_12_64_4096_1_4096_64_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_144_12_64_4096_1_4096_64_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [63:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [63:0] d;
  output [11:0] wadr;
  input clken_d;
  input [63:0] d_d;
  output [63:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_143_12_64_4096_1_4096_64_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_143_12_64_4096_1_4096_64_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [63:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [63:0] d;
  output [11:0] wadr;
  input clken_d;
  input [63:0] d_d;
  output [63:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_142_12_64_4096_1_4096_64_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_142_12_64_4096_1_4096_64_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [63:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [63:0] d;
  output [11:0] wadr;
  input clken_d;
  input [63:0] d_d;
  output [63:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_141_12_64_4096_1_4096_64_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_141_12_64_4096_1_4096_64_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [63:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [63:0] d;
  output [11:0] wadr;
  input clken_d;
  input [63:0] d_d;
  output [63:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_140_12_64_4096_1_4096_64_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_140_12_64_4096_1_4096_64_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [63:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [63:0] d;
  output [11:0] wadr;
  input clken_d;
  input [63:0] d_d;
  output [63:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_139_12_64_4096_1_4096_64_1_gen
// ------------------------------------------------------------------


module PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_139_12_64_4096_1_4096_64_1_gen
    (
  clken, q, re, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, re_d, wadr_d, we_d,
      writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [63:0] q;
  output re;
  output [11:0] radr;
  output we;
  output [63:0] d;
  output [11:0] wadr;
  input clken_d;
  input [63:0] d_d;
  output [63:0] q_d;
  input [11:0] radr_d;
  input re_d;
  input [11:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_PECoreRun_fsm
//  FSM Module
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_PECoreRun_fsm (
  clk, rst, PECoreRun_wen, fsm_output
);
  input clk;
  input rst;
  input PECoreRun_wen;
  output fsm_output;
  reg fsm_output;


  // FSM State Type Declaration for PECore_PECore_PECoreRun_PECoreRun_fsm_1
  parameter
    PECoreRun_rlp_C_0 = 1'd0,
    while_C_0 = 1'd1;

  reg  state_var;
  reg  state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : PECore_PECore_PECoreRun_PECoreRun_fsm_1
    case (state_var)
      while_C_0 : begin
        fsm_output = 1'b1;
        state_var_NS = while_C_0;
      end
      // PECoreRun_rlp_C_0
      default : begin
        fsm_output = 1'b0;
        state_var_NS = while_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      state_var <= PECoreRun_rlp_C_0;
    end
    else if ( PECoreRun_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_staller
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_staller (
  clk, rst, PECoreRun_wen, PECoreRun_wten, act_port_Push_mioi_wen_comp, rva_out_Push_mioi_wen_comp
);
  input clk;
  input rst;
  output PECoreRun_wen;
  output PECoreRun_wten;
  input act_port_Push_mioi_wen_comp;
  input rva_out_Push_mioi_wen_comp;


  // Interconnect Declarations
  reg PECoreRun_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign PECoreRun_wen = act_port_Push_mioi_wen_comp & rva_out_Push_mioi_wen_comp;
  assign PECoreRun_wten = PECoreRun_wten_reg;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECoreRun_wten_reg <= 1'b0;
    end
    else begin
      PECoreRun_wten_reg <= ~ PECoreRun_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_wait_dp
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_wait_dp (
  weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d, weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d,
      weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d, weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d,
      weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d, weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d,
      weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d, weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d,
      ProductSum_for_acc_11_cmp_en, ProductSum_for_acc_9_cmp_en, PECoreRun_wen, weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo,
      weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_unreg, weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo,
      weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_unreg, weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo,
      weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_unreg, weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo,
      weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_unreg, weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo,
      weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_unreg, weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo,
      weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_unreg, weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo,
      weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_unreg, weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo,
      weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_unreg, ProductSum_for_acc_11_cmp_cgo,
      ProductSum_for_acc_11_cmp_cgo_ir_unreg, ProductSum_for_acc_9_cmp_cgo, ProductSum_for_acc_9_cmp_cgo_ir_unreg
);
  output weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d;
  output weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d;
  output weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d;
  output weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d;
  output weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d;
  output weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d;
  output weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d;
  output weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d;
  output ProductSum_for_acc_11_cmp_en;
  output ProductSum_for_acc_9_cmp_en;
  input PECoreRun_wen;
  input weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo;
  input weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo;
  input weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo;
  input weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo;
  input weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo;
  input weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo;
  input weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo;
  input weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_unreg;
  input weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo;
  input weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_unreg;
  input ProductSum_for_acc_11_cmp_cgo;
  input ProductSum_for_acc_11_cmp_cgo_ir_unreg;
  input ProductSum_for_acc_9_cmp_cgo;
  input ProductSum_for_acc_9_cmp_cgo_ir_unreg;



  // Interconnect Declarations for Component Instantiations 
  assign weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo
      | weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo
      | weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo
      | weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo
      | weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo
      | weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo
      | weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo
      | weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_unreg);
  assign weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d = PECoreRun_wen & (weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo
      | weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_unreg);
  assign ProductSum_for_acc_11_cmp_en = ~(PECoreRun_wen & (ProductSum_for_acc_11_cmp_cgo
      | ProductSum_for_acc_11_cmp_cgo_ir_unreg));
  assign ProductSum_for_acc_9_cmp_en = ~(PECoreRun_wen & (ProductSum_for_acc_9_cmp_cgo
      | ProductSum_for_acc_9_cmp_cgo_ir_unreg));
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_dp
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_dp (
  clk, rst, rva_out_Push_mioi_oswt, rva_out_Push_mioi_wen_comp, rva_out_Push_mioi_biwt,
      rva_out_Push_mioi_bdwt, rva_out_Push_mioi_bcwt
);
  input clk;
  input rst;
  input rva_out_Push_mioi_oswt;
  output rva_out_Push_mioi_wen_comp;
  input rva_out_Push_mioi_biwt;
  input rva_out_Push_mioi_bdwt;
  output rva_out_Push_mioi_bcwt;
  reg rva_out_Push_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign rva_out_Push_mioi_wen_comp = (~ rva_out_Push_mioi_oswt) | rva_out_Push_mioi_biwt
      | rva_out_Push_mioi_bcwt;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      rva_out_Push_mioi_bcwt <= ~((~(rva_out_Push_mioi_bcwt | rva_out_Push_mioi_biwt))
          | rva_out_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl (
  PECoreRun_wen, rva_out_Push_mioi_oswt, rva_out_Push_mioi_biwt, rva_out_Push_mioi_bdwt,
      rva_out_Push_mioi_bcwt, rva_out_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct,
      rva_out_Push_mioi_ccs_ccore_done_sync_vld, rva_out_Push_mioi_oswt_pff
);
  input PECoreRun_wen;
  input rva_out_Push_mioi_oswt;
  output rva_out_Push_mioi_biwt;
  output rva_out_Push_mioi_bdwt;
  input rva_out_Push_mioi_bcwt;
  output rva_out_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct;
  input rva_out_Push_mioi_ccs_ccore_done_sync_vld;
  input rva_out_Push_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign rva_out_Push_mioi_bdwt = rva_out_Push_mioi_oswt & PECoreRun_wen;
  assign rva_out_Push_mioi_biwt = rva_out_Push_mioi_oswt & (~ rva_out_Push_mioi_bcwt)
      & rva_out_Push_mioi_ccs_ccore_done_sync_vld;
  assign rva_out_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct = PECoreRun_wen
      & rva_out_Push_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_dp (
  clk, rst, start_PopNB_mioi_data_rsc_z_mxwt, start_PopNB_mioi_return_rsc_z_mxwt,
      start_PopNB_mioi_biwt, start_PopNB_mioi_bdwt, start_PopNB_mioi_data_rsc_z,
      start_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output start_PopNB_mioi_data_rsc_z_mxwt;
  output start_PopNB_mioi_return_rsc_z_mxwt;
  input start_PopNB_mioi_biwt;
  input start_PopNB_mioi_bdwt;
  input start_PopNB_mioi_data_rsc_z;
  input start_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg start_PopNB_mioi_bcwt;
  reg start_PopNB_mioi_data_rsc_z_bfwt;
  reg start_PopNB_mioi_return_rsc_z_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign start_PopNB_mioi_data_rsc_z_mxwt = MUX_s_1_2_2(start_PopNB_mioi_data_rsc_z,
      start_PopNB_mioi_data_rsc_z_bfwt, start_PopNB_mioi_bcwt);
  assign start_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(start_PopNB_mioi_return_rsc_z,
      start_PopNB_mioi_return_rsc_z_bfwt, start_PopNB_mioi_bcwt);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      start_PopNB_mioi_bcwt <= 1'b0;
    end
    else begin
      start_PopNB_mioi_bcwt <= ~((~(start_PopNB_mioi_bcwt | start_PopNB_mioi_biwt))
          | start_PopNB_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      start_PopNB_mioi_data_rsc_z_bfwt <= 1'b0;
      start_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else if ( start_PopNB_mioi_biwt ) begin
      start_PopNB_mioi_data_rsc_z_bfwt <= start_PopNB_mioi_data_rsc_z;
      start_PopNB_mioi_return_rsc_z_bfwt <= start_PopNB_mioi_return_rsc_z;
    end
  end

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_ctrl (
  PECoreRun_wen, PECoreRun_wten, start_PopNB_mioi_oswt, start_PopNB_mioi_biwt, start_PopNB_mioi_bdwt,
      start_PopNB_mioi_biwt_pff, start_PopNB_mioi_oswt_pff
);
  input PECoreRun_wen;
  input PECoreRun_wten;
  input start_PopNB_mioi_oswt;
  output start_PopNB_mioi_biwt;
  output start_PopNB_mioi_bdwt;
  output start_PopNB_mioi_biwt_pff;
  input start_PopNB_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign start_PopNB_mioi_bdwt = start_PopNB_mioi_oswt & PECoreRun_wen;
  assign start_PopNB_mioi_biwt = (~ PECoreRun_wten) & start_PopNB_mioi_oswt;
  assign start_PopNB_mioi_biwt_pff = PECoreRun_wen & start_PopNB_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_dp
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_dp (
  clk, rst, act_port_Push_mioi_oswt, act_port_Push_mioi_wen_comp, act_port_Push_mioi_biwt,
      act_port_Push_mioi_bdwt, act_port_Push_mioi_bcwt
);
  input clk;
  input rst;
  input act_port_Push_mioi_oswt;
  output act_port_Push_mioi_wen_comp;
  input act_port_Push_mioi_biwt;
  input act_port_Push_mioi_bdwt;
  output act_port_Push_mioi_bcwt;
  reg act_port_Push_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign act_port_Push_mioi_wen_comp = (~ act_port_Push_mioi_oswt) | act_port_Push_mioi_biwt
      | act_port_Push_mioi_bcwt;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      act_port_Push_mioi_bcwt <= ~((~(act_port_Push_mioi_bcwt | act_port_Push_mioi_biwt))
          | act_port_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_ctrl (
  PECoreRun_wen, act_port_Push_mioi_oswt, act_port_Push_mioi_biwt, act_port_Push_mioi_bdwt,
      act_port_Push_mioi_bcwt, act_port_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct,
      act_port_Push_mioi_ccs_ccore_done_sync_vld, act_port_Push_mioi_oswt_pff
);
  input PECoreRun_wen;
  input act_port_Push_mioi_oswt;
  output act_port_Push_mioi_biwt;
  output act_port_Push_mioi_bdwt;
  input act_port_Push_mioi_bcwt;
  output act_port_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct;
  input act_port_Push_mioi_ccs_ccore_done_sync_vld;
  input act_port_Push_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign act_port_Push_mioi_bdwt = act_port_Push_mioi_oswt & PECoreRun_wen;
  assign act_port_Push_mioi_biwt = act_port_Push_mioi_oswt & (~ act_port_Push_mioi_bcwt)
      & act_port_Push_mioi_ccs_ccore_done_sync_vld;
  assign act_port_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct = PECoreRun_wen
      & act_port_Push_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_dp
    (
  clk, rst, input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt,
      input_port_PopNB_mioi_return_rsc_z_mxwt, input_port_PopNB_mioi_biwt, input_port_PopNB_mioi_bdwt,
      input_port_PopNB_mioi_data_data_data_rsc_z, input_port_PopNB_mioi_data_logical_addr_rsc_z,
      input_port_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output [63:0] input_port_PopNB_mioi_data_data_data_rsc_z_mxwt;
  output [7:0] input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt;
  output input_port_PopNB_mioi_return_rsc_z_mxwt;
  input input_port_PopNB_mioi_biwt;
  input input_port_PopNB_mioi_bdwt;
  input [63:0] input_port_PopNB_mioi_data_data_data_rsc_z;
  input [7:0] input_port_PopNB_mioi_data_logical_addr_rsc_z;
  input input_port_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg input_port_PopNB_mioi_bcwt;
  reg [63:0] input_port_PopNB_mioi_data_data_data_rsc_z_bfwt;
  reg [7:0] input_port_PopNB_mioi_data_logical_addr_rsc_z_bfwt;
  reg input_port_PopNB_mioi_return_rsc_z_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign input_port_PopNB_mioi_data_data_data_rsc_z_mxwt = MUX_v_64_2_2(input_port_PopNB_mioi_data_data_data_rsc_z,
      input_port_PopNB_mioi_data_data_data_rsc_z_bfwt, input_port_PopNB_mioi_bcwt);
  assign input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt = MUX_v_8_2_2(input_port_PopNB_mioi_data_logical_addr_rsc_z,
      input_port_PopNB_mioi_data_logical_addr_rsc_z_bfwt, input_port_PopNB_mioi_bcwt);
  assign input_port_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(input_port_PopNB_mioi_return_rsc_z,
      input_port_PopNB_mioi_return_rsc_z_bfwt, input_port_PopNB_mioi_bcwt);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_port_PopNB_mioi_bcwt <= 1'b0;
    end
    else begin
      input_port_PopNB_mioi_bcwt <= ~((~(input_port_PopNB_mioi_bcwt | input_port_PopNB_mioi_biwt))
          | input_port_PopNB_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_port_PopNB_mioi_data_data_data_rsc_z_bfwt <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      input_port_PopNB_mioi_data_logical_addr_rsc_z_bfwt <= 8'b00000000;
      input_port_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else if ( input_port_PopNB_mioi_biwt ) begin
      input_port_PopNB_mioi_data_data_data_rsc_z_bfwt <= input_port_PopNB_mioi_data_data_data_rsc_z;
      input_port_PopNB_mioi_data_logical_addr_rsc_z_bfwt <= input_port_PopNB_mioi_data_logical_addr_rsc_z;
      input_port_PopNB_mioi_return_rsc_z_bfwt <= input_port_PopNB_mioi_return_rsc_z;
    end
  end

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input  sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_ctrl
    (
  PECoreRun_wen, PECoreRun_wten, input_port_PopNB_mioi_oswt, input_port_PopNB_mioi_biwt,
      input_port_PopNB_mioi_bdwt, input_port_PopNB_mioi_biwt_pff, input_port_PopNB_mioi_oswt_pff
);
  input PECoreRun_wen;
  input PECoreRun_wten;
  input input_port_PopNB_mioi_oswt;
  output input_port_PopNB_mioi_biwt;
  output input_port_PopNB_mioi_bdwt;
  output input_port_PopNB_mioi_biwt_pff;
  input input_port_PopNB_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign input_port_PopNB_mioi_bdwt = input_port_PopNB_mioi_oswt & PECoreRun_wen;
  assign input_port_PopNB_mioi_biwt = (~ PECoreRun_wten) & input_port_PopNB_mioi_oswt;
  assign input_port_PopNB_mioi_biwt_pff = PECoreRun_wen & input_port_PopNB_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp (
  clk, rst, rva_in_PopNB_mioi_data_data_rsc_z_mxwt, rva_in_PopNB_mioi_data_addr_rsc_z_mxwt,
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt, rva_in_PopNB_mioi_return_rsc_z_mxwt,
      rva_in_PopNB_mioi_biwt, rva_in_PopNB_mioi_bdwt, rva_in_PopNB_mioi_data_data_rsc_z,
      rva_in_PopNB_mioi_data_addr_rsc_z, rva_in_PopNB_mioi_data_rw_rsc_z, rva_in_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output [63:0] rva_in_PopNB_mioi_data_data_rsc_z_mxwt;
  output [19:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt;
  output rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  output rva_in_PopNB_mioi_return_rsc_z_mxwt;
  input rva_in_PopNB_mioi_biwt;
  input rva_in_PopNB_mioi_bdwt;
  input [63:0] rva_in_PopNB_mioi_data_data_rsc_z;
  input [23:0] rva_in_PopNB_mioi_data_addr_rsc_z;
  input rva_in_PopNB_mioi_data_rw_rsc_z;
  input rva_in_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg rva_in_PopNB_mioi_bcwt;
  reg [63:0] rva_in_PopNB_mioi_data_data_rsc_z_bfwt;
  reg rva_in_PopNB_mioi_data_rw_rsc_z_bfwt;
  reg rva_in_PopNB_mioi_return_rsc_z_bfwt;
  reg [19:0] rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_23_4;


  // Interconnect Declarations for Component Instantiations 
  assign rva_in_PopNB_mioi_data_data_rsc_z_mxwt = MUX_v_64_2_2(rva_in_PopNB_mioi_data_data_rsc_z,
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt, rva_in_PopNB_mioi_bcwt);
  assign rva_in_PopNB_mioi_data_rw_rsc_z_mxwt = MUX_s_1_2_2(rva_in_PopNB_mioi_data_rw_rsc_z,
      rva_in_PopNB_mioi_data_rw_rsc_z_bfwt, rva_in_PopNB_mioi_bcwt);
  assign rva_in_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(rva_in_PopNB_mioi_return_rsc_z,
      rva_in_PopNB_mioi_return_rsc_z_bfwt, rva_in_PopNB_mioi_bcwt);
  assign rva_in_PopNB_mioi_data_addr_rsc_z_mxwt = MUX_v_20_2_2((rva_in_PopNB_mioi_data_addr_rsc_z[23:4]),
      rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_23_4, rva_in_PopNB_mioi_bcwt);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_PopNB_mioi_bcwt <= 1'b0;
    end
    else begin
      rva_in_PopNB_mioi_bcwt <= ~((~(rva_in_PopNB_mioi_bcwt | rva_in_PopNB_mioi_biwt))
          | rva_in_PopNB_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_23_4 <= 20'b00000000000000000000;
      rva_in_PopNB_mioi_data_rw_rsc_z_bfwt <= 1'b0;
      rva_in_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else if ( rva_in_PopNB_mioi_biwt ) begin
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt <= rva_in_PopNB_mioi_data_data_rsc_z;
      rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_23_4 <= rva_in_PopNB_mioi_data_addr_rsc_z[23:4];
      rva_in_PopNB_mioi_data_rw_rsc_z_bfwt <= rva_in_PopNB_mioi_data_rw_rsc_z;
      rva_in_PopNB_mioi_return_rsc_z_bfwt <= rva_in_PopNB_mioi_return_rsc_z;
    end
  end

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [19:0] MUX_v_20_2_2;
    input [19:0] input_0;
    input [19:0] input_1;
    input  sel;
    reg [19:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_20_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input  sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl (
  PECoreRun_wen, PECoreRun_wten, rva_in_PopNB_mioi_oswt, rva_in_PopNB_mioi_biwt,
      rva_in_PopNB_mioi_bdwt, rva_in_PopNB_mioi_biwt_pff, rva_in_PopNB_mioi_oswt_pff
);
  input PECoreRun_wen;
  input PECoreRun_wten;
  input rva_in_PopNB_mioi_oswt;
  output rva_in_PopNB_mioi_biwt;
  output rva_in_PopNB_mioi_bdwt;
  output rva_in_PopNB_mioi_biwt_pff;
  input rva_in_PopNB_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign rva_in_PopNB_mioi_bdwt = rva_in_PopNB_mioi_oswt & PECoreRun_wen;
  assign rva_in_PopNB_mioi_biwt = (~ PECoreRun_wten) & rva_in_PopNB_mioi_oswt;
  assign rva_in_PopNB_mioi_biwt_pff = PECoreRun_wen & rva_in_PopNB_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_rva_out_Push_mioi
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_rva_out_Push_mioi (
  clk, rst, rva_out_vld, rva_out_rdy, rva_out_dat, PECoreRun_wen, rva_out_Push_mioi_oswt,
      rva_out_Push_mioi_wen_comp, rva_out_Push_mioi_m_data_rsc_dat_PECoreRun, rva_out_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output rva_out_vld;
  input rva_out_rdy;
  output [63:0] rva_out_dat;
  input PECoreRun_wen;
  input rva_out_Push_mioi_oswt;
  output rva_out_Push_mioi_wen_comp;
  input [63:0] rva_out_Push_mioi_m_data_rsc_dat_PECoreRun;
  input rva_out_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire rva_out_Push_mioi_biwt;
  wire rva_out_Push_mioi_bdwt;
  wire rva_out_Push_mioi_bcwt;
  wire rva_out_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct;
  wire rva_out_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  PECore_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push
      rva_out_Push_mioi (
      .this_vld(rva_out_vld),
      .this_rdy(rva_out_rdy),
      .this_dat(rva_out_dat),
      .m_data_rsc_dat(rva_out_Push_mioi_m_data_rsc_dat_PECoreRun),
      .ccs_ccore_start_rsc_dat(rva_out_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct),
      .ccs_ccore_done_sync_vld(rva_out_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  PECore_PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl_inst
      (
      .PECoreRun_wen(PECoreRun_wen),
      .rva_out_Push_mioi_oswt(rva_out_Push_mioi_oswt),
      .rva_out_Push_mioi_biwt(rva_out_Push_mioi_biwt),
      .rva_out_Push_mioi_bdwt(rva_out_Push_mioi_bdwt),
      .rva_out_Push_mioi_bcwt(rva_out_Push_mioi_bcwt),
      .rva_out_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct(rva_out_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct),
      .rva_out_Push_mioi_ccs_ccore_done_sync_vld(rva_out_Push_mioi_ccs_ccore_done_sync_vld),
      .rva_out_Push_mioi_oswt_pff(rva_out_Push_mioi_oswt_pff)
    );
  PECore_PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_dp PECore_PECoreRun_rva_out_Push_mioi_rva_out_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_out_Push_mioi_oswt(rva_out_Push_mioi_oswt),
      .rva_out_Push_mioi_wen_comp(rva_out_Push_mioi_wen_comp),
      .rva_out_Push_mioi_biwt(rva_out_Push_mioi_biwt),
      .rva_out_Push_mioi_bdwt(rva_out_Push_mioi_bdwt),
      .rva_out_Push_mioi_bcwt(rva_out_Push_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_start_PopNB_mioi
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_start_PopNB_mioi (
  clk, rst, start_vld, start_rdy, start_dat, PECoreRun_wen, PECoreRun_wten, start_PopNB_mioi_oswt,
      start_PopNB_mioi_data_rsc_z_mxwt, start_PopNB_mioi_return_rsc_z_mxwt, start_PopNB_mioi_oswt_pff
);
  input clk;
  input rst;
  input start_vld;
  output start_rdy;
  input start_dat;
  input PECoreRun_wen;
  input PECoreRun_wten;
  input start_PopNB_mioi_oswt;
  output start_PopNB_mioi_data_rsc_z_mxwt;
  output start_PopNB_mioi_return_rsc_z_mxwt;
  input start_PopNB_mioi_oswt_pff;


  // Interconnect Declarations
  wire start_PopNB_mioi_biwt;
  wire start_PopNB_mioi_bdwt;
  wire start_PopNB_mioi_data_rsc_z;
  wire start_PopNB_mioi_return_rsc_z;
  wire start_PopNB_mioi_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  PECore_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB  start_PopNB_mioi
      (
      .this_vld(start_vld),
      .this_rdy(start_rdy),
      .this_dat(start_dat),
      .data_rsc_z(start_PopNB_mioi_data_rsc_z),
      .return_rsc_z(start_PopNB_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(start_PopNB_mioi_biwt_iff),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  PECore_PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_ctrl PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_ctrl_inst
      (
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .start_PopNB_mioi_oswt(start_PopNB_mioi_oswt),
      .start_PopNB_mioi_biwt(start_PopNB_mioi_biwt),
      .start_PopNB_mioi_bdwt(start_PopNB_mioi_bdwt),
      .start_PopNB_mioi_biwt_pff(start_PopNB_mioi_biwt_iff),
      .start_PopNB_mioi_oswt_pff(start_PopNB_mioi_oswt_pff)
    );
  PECore_PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_dp PECore_PECoreRun_start_PopNB_mioi_start_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .start_PopNB_mioi_data_rsc_z_mxwt(start_PopNB_mioi_data_rsc_z_mxwt),
      .start_PopNB_mioi_return_rsc_z_mxwt(start_PopNB_mioi_return_rsc_z_mxwt),
      .start_PopNB_mioi_biwt(start_PopNB_mioi_biwt),
      .start_PopNB_mioi_bdwt(start_PopNB_mioi_bdwt),
      .start_PopNB_mioi_data_rsc_z(start_PopNB_mioi_data_rsc_z),
      .start_PopNB_mioi_return_rsc_z(start_PopNB_mioi_return_rsc_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_act_port_Push_mioi
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_act_port_Push_mioi (
  clk, rst, act_port_vld, act_port_rdy, act_port_dat, PECoreRun_wen, act_port_Push_mioi_oswt,
      act_port_Push_mioi_wen_comp, act_port_Push_mioi_m_data_rsc_dat_PECoreRun, act_port_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output act_port_vld;
  input act_port_rdy;
  output [255:0] act_port_dat;
  input PECoreRun_wen;
  input act_port_Push_mioi_oswt;
  output act_port_Push_mioi_wen_comp;
  input [255:0] act_port_Push_mioi_m_data_rsc_dat_PECoreRun;
  input act_port_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire act_port_Push_mioi_biwt;
  wire act_port_Push_mioi_bdwt;
  wire act_port_Push_mioi_bcwt;
  wire act_port_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct;
  wire act_port_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  PECore_Connections_OutBlocking_spec_ActVectorType_Connections_SYN_PORT_Push  act_port_Push_mioi
      (
      .this_vld(act_port_vld),
      .this_rdy(act_port_rdy),
      .this_dat(act_port_dat),
      .m_data_rsc_dat(act_port_Push_mioi_m_data_rsc_dat_PECoreRun),
      .ccs_ccore_start_rsc_dat(act_port_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct),
      .ccs_ccore_done_sync_vld(act_port_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  PECore_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_ctrl PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_ctrl_inst
      (
      .PECoreRun_wen(PECoreRun_wen),
      .act_port_Push_mioi_oswt(act_port_Push_mioi_oswt),
      .act_port_Push_mioi_biwt(act_port_Push_mioi_biwt),
      .act_port_Push_mioi_bdwt(act_port_Push_mioi_bdwt),
      .act_port_Push_mioi_bcwt(act_port_Push_mioi_bcwt),
      .act_port_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct(act_port_Push_mioi_ccs_ccore_start_rsc_dat_PECoreRun_sct),
      .act_port_Push_mioi_ccs_ccore_done_sync_vld(act_port_Push_mioi_ccs_ccore_done_sync_vld),
      .act_port_Push_mioi_oswt_pff(act_port_Push_mioi_oswt_pff)
    );
  PECore_PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_dp PECore_PECoreRun_act_port_Push_mioi_act_port_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .act_port_Push_mioi_oswt(act_port_Push_mioi_oswt),
      .act_port_Push_mioi_wen_comp(act_port_Push_mioi_wen_comp),
      .act_port_Push_mioi_biwt(act_port_Push_mioi_biwt),
      .act_port_Push_mioi_bdwt(act_port_Push_mioi_bdwt),
      .act_port_Push_mioi_bcwt(act_port_Push_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_input_port_PopNB_mioi
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_input_port_PopNB_mioi (
  clk, rst, input_port_vld, input_port_rdy, input_port_dat, PECoreRun_wen, PECoreRun_wten,
      input_port_PopNB_mioi_oswt, input_port_PopNB_mioi_data_data_data_rsc_z_mxwt,
      input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt, input_port_PopNB_mioi_return_rsc_z_mxwt,
      input_port_PopNB_mioi_oswt_pff
);
  input clk;
  input rst;
  input input_port_vld;
  output input_port_rdy;
  input [73:0] input_port_dat;
  input PECoreRun_wen;
  input PECoreRun_wten;
  input input_port_PopNB_mioi_oswt;
  output [63:0] input_port_PopNB_mioi_data_data_data_rsc_z_mxwt;
  output [7:0] input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt;
  output input_port_PopNB_mioi_return_rsc_z_mxwt;
  input input_port_PopNB_mioi_oswt_pff;


  // Interconnect Declarations
  wire input_port_PopNB_mioi_biwt;
  wire input_port_PopNB_mioi_bdwt;
  wire [63:0] input_port_PopNB_mioi_data_data_data_rsc_z;
  wire [7:0] input_port_PopNB_mioi_data_logical_addr_rsc_z;
  wire input_port_PopNB_mioi_return_rsc_z;
  wire input_port_PopNB_mioi_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  PECore_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB  input_port_PopNB_mioi
      (
      .this_vld(input_port_vld),
      .this_rdy(input_port_rdy),
      .this_dat(input_port_dat),
      .data_data_data_rsc_z(input_port_PopNB_mioi_data_data_data_rsc_z),
      .data_logical_addr_rsc_z(input_port_PopNB_mioi_data_logical_addr_rsc_z),
      .return_rsc_z(input_port_PopNB_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(input_port_PopNB_mioi_biwt_iff),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  PECore_PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_ctrl PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_ctrl_inst
      (
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .input_port_PopNB_mioi_oswt(input_port_PopNB_mioi_oswt),
      .input_port_PopNB_mioi_biwt(input_port_PopNB_mioi_biwt),
      .input_port_PopNB_mioi_bdwt(input_port_PopNB_mioi_bdwt),
      .input_port_PopNB_mioi_biwt_pff(input_port_PopNB_mioi_biwt_iff),
      .input_port_PopNB_mioi_oswt_pff(input_port_PopNB_mioi_oswt_pff)
    );
  PECore_PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_dp PECore_PECoreRun_input_port_PopNB_mioi_input_port_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .input_port_PopNB_mioi_data_data_data_rsc_z_mxwt(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt),
      .input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt(input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt),
      .input_port_PopNB_mioi_return_rsc_z_mxwt(input_port_PopNB_mioi_return_rsc_z_mxwt),
      .input_port_PopNB_mioi_biwt(input_port_PopNB_mioi_biwt),
      .input_port_PopNB_mioi_bdwt(input_port_PopNB_mioi_bdwt),
      .input_port_PopNB_mioi_data_data_data_rsc_z(input_port_PopNB_mioi_data_data_data_rsc_z),
      .input_port_PopNB_mioi_data_logical_addr_rsc_z(input_port_PopNB_mioi_data_logical_addr_rsc_z),
      .input_port_PopNB_mioi_return_rsc_z(input_port_PopNB_mioi_return_rsc_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun_rva_in_PopNB_mioi
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun_rva_in_PopNB_mioi (
  clk, rst, rva_in_vld, rva_in_rdy, rva_in_dat, PECoreRun_wen, PECoreRun_wten, rva_in_PopNB_mioi_oswt,
      rva_in_PopNB_mioi_data_data_rsc_z_mxwt, rva_in_PopNB_mioi_data_addr_rsc_z_mxwt,
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt, rva_in_PopNB_mioi_return_rsc_z_mxwt,
      rva_in_PopNB_mioi_oswt_pff
);
  input clk;
  input rst;
  input rva_in_vld;
  output rva_in_rdy;
  input [96:0] rva_in_dat;
  input PECoreRun_wen;
  input PECoreRun_wten;
  input rva_in_PopNB_mioi_oswt;
  output [63:0] rva_in_PopNB_mioi_data_data_rsc_z_mxwt;
  output [19:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt;
  output rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  output rva_in_PopNB_mioi_return_rsc_z_mxwt;
  input rva_in_PopNB_mioi_oswt_pff;


  // Interconnect Declarations
  wire rva_in_PopNB_mioi_biwt;
  wire rva_in_PopNB_mioi_bdwt;
  wire [63:0] rva_in_PopNB_mioi_data_data_rsc_z;
  wire [23:0] rva_in_PopNB_mioi_data_addr_rsc_z;
  wire rva_in_PopNB_mioi_data_rw_rsc_z;
  wire rva_in_PopNB_mioi_return_rsc_z;
  wire [19:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt_pconst;
  wire rva_in_PopNB_mioi_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  PECore_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB
      rva_in_PopNB_mioi (
      .this_vld(rva_in_vld),
      .this_rdy(rva_in_rdy),
      .this_dat(rva_in_dat),
      .data_data_rsc_z(rva_in_PopNB_mioi_data_data_rsc_z),
      .data_addr_rsc_z(rva_in_PopNB_mioi_data_addr_rsc_z),
      .data_rw_rsc_z(rva_in_PopNB_mioi_data_rw_rsc_z),
      .return_rsc_z(rva_in_PopNB_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(rva_in_PopNB_mioi_biwt_iff),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  PECore_PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl_inst
      (
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .rva_in_PopNB_mioi_oswt(rva_in_PopNB_mioi_oswt),
      .rva_in_PopNB_mioi_biwt(rva_in_PopNB_mioi_biwt),
      .rva_in_PopNB_mioi_bdwt(rva_in_PopNB_mioi_bdwt),
      .rva_in_PopNB_mioi_biwt_pff(rva_in_PopNB_mioi_biwt_iff),
      .rva_in_PopNB_mioi_oswt_pff(rva_in_PopNB_mioi_oswt_pff)
    );
  PECore_PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp PECore_PECoreRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_in_PopNB_mioi_data_data_rsc_z_mxwt(rva_in_PopNB_mioi_data_data_rsc_z_mxwt),
      .rva_in_PopNB_mioi_data_addr_rsc_z_mxwt(rva_in_PopNB_mioi_data_addr_rsc_z_mxwt_pconst),
      .rva_in_PopNB_mioi_data_rw_rsc_z_mxwt(rva_in_PopNB_mioi_data_rw_rsc_z_mxwt),
      .rva_in_PopNB_mioi_return_rsc_z_mxwt(rva_in_PopNB_mioi_return_rsc_z_mxwt),
      .rva_in_PopNB_mioi_biwt(rva_in_PopNB_mioi_biwt),
      .rva_in_PopNB_mioi_bdwt(rva_in_PopNB_mioi_bdwt),
      .rva_in_PopNB_mioi_data_data_rsc_z(rva_in_PopNB_mioi_data_data_rsc_z),
      .rva_in_PopNB_mioi_data_addr_rsc_z(rva_in_PopNB_mioi_data_addr_rsc_z),
      .rva_in_PopNB_mioi_data_rw_rsc_z(rva_in_PopNB_mioi_data_rw_rsc_z),
      .rva_in_PopNB_mioi_return_rsc_z(rva_in_PopNB_mioi_return_rsc_z)
    );
  assign rva_in_PopNB_mioi_data_addr_rsc_z_mxwt = rva_in_PopNB_mioi_data_addr_rsc_z_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore_PECore_PECoreRun
// ------------------------------------------------------------------


module PECore_PECore_PECoreRun (
  clk, rst, start_vld, start_rdy, start_dat, input_port_vld, input_port_rdy, input_port_dat,
      rva_in_vld, rva_in_rdy, rva_in_dat, rva_out_vld, rva_out_rdy, rva_out_dat,
      act_port_vld, act_port_rdy, act_port_dat, SC_SRAM_CONFIG, weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d,
      weight_mem_banks_bank_a0_a0_a0_a_rsci_d_d, weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d,
      weight_mem_banks_bank_a0_a0_a0_a_rsci_radr_d, weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d,
      weight_mem_banks_bank_a0_a0_a1_a_rsci_d_d, weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d,
      weight_mem_banks_bank_a0_a0_a1_a_rsci_radr_d, weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d,
      weight_mem_banks_bank_a0_a1_a0_a_rsci_d_d, weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d,
      weight_mem_banks_bank_a0_a1_a0_a_rsci_radr_d, weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d,
      weight_mem_banks_bank_a0_a1_a1_a_rsci_d_d, weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d,
      weight_mem_banks_bank_a0_a1_a1_a_rsci_radr_d, weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d,
      weight_mem_banks_bank_a1_a0_a0_a_rsci_d_d, weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d,
      weight_mem_banks_bank_a1_a0_a0_a_rsci_radr_d, weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d,
      weight_mem_banks_bank_a1_a0_a1_a_rsci_d_d, weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d,
      weight_mem_banks_bank_a1_a0_a1_a_rsci_radr_d, weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d,
      weight_mem_banks_bank_a1_a1_a0_a_rsci_d_d, weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d,
      weight_mem_banks_bank_a1_a1_a0_a_rsci_radr_d, weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d,
      weight_mem_banks_bank_a1_a1_a1_a_rsci_d_d, weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d,
      weight_mem_banks_bank_a1_a1_a1_a_rsci_radr_d, ProductSum_for_acc_11_cmp_a,
      ProductSum_for_acc_11_cmp_en, ProductSum_for_acc_11_cmp_z, ProductSum_for_acc_10_cmp_a,
      ProductSum_for_acc_10_cmp_z, ProductSum_for_acc_9_cmp_a0, ProductSum_for_acc_9_cmp_b0,
      ProductSum_for_acc_9_cmp_c0, ProductSum_for_acc_9_cmp_en, ProductSum_for_acc_9_cmp_z,
      ProductSum_for_acc_8_cmp_a0, ProductSum_for_acc_8_cmp_b0, ProductSum_for_acc_8_cmp_c0,
      ProductSum_for_acc_8_cmp_z, PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_a,
      PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_z, PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_4_cmp_a,
      PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_4_cmp_z, PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_a0,
      PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_b0, PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_c0,
      PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_z, PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_a0,
      PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_b0, PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_c0,
      PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_z, PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_a,
      PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_z, PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_4_cmp_a,
      PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_4_cmp_z, PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_a0,
      PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_b0, PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_c0,
      PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_z, PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_a0,
      PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_b0, PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_c0,
      PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_z, PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_a,
      PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_z, PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_4_cmp_a,
      PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_4_cmp_z, PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_a0,
      PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_b0, PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_c0,
      PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_z, PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_a0,
      PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_b0, PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_c0,
      PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_z, PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_a,
      PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_z, PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_4_cmp_a,
      PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_4_cmp_z, PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_a0,
      PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_b0, PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_c0,
      PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_z, PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_a0,
      PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_b0, PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_c0,
      PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_z, PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_a,
      PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_load, PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_z,
      PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_a, PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_b,
      PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_z, PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_a0,
      PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_b0, PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_c0,
      PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_z, PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_a0,
      PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_b0, PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_c0,
      PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_z, PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_a,
      PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_z, PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_4_cmp_a,
      PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_4_cmp_z, PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_a0,
      PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_b0, PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_c0,
      PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_z, PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_a0,
      PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_b0, PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_c0,
      PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_z, PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_a,
      PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_z, PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_a,
      PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_z, PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_a0,
      PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_b0, PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_c0,
      PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_z, PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_a0,
      PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_b0, PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_c0,
      PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_z, ProductSum_for_acc_11_cmp_b_pff,
      ProductSum_for_acc_11_cmp_load_pff, ProductSum_for_acc_11_cmp_datavalid_pff,
      ProductSum_for_acc_10_cmp_b_pff, ProductSum_for_acc_9_cmp_a1_pff, ProductSum_for_acc_9_cmp_b1_pff,
      ProductSum_for_acc_9_cmp_c1_pff, ProductSum_for_acc_9_cmp_load_pff, ProductSum_for_acc_9_cmp_datavalid_pff,
      ProductSum_for_acc_8_cmp_a1_pff, ProductSum_for_acc_8_cmp_b1_pff, ProductSum_for_acc_8_cmp_c1_pff,
      PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_load_pff, PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_load_pff,
      PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_load_pff, PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_load_pff,
      PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_load_pff, PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_load_pff,
      PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_load_pff, PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_load_pff,
      PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_load_pff, PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_load_pff,
      PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_load_pff, PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_load_pff,
      PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_load_pff, weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_pff,
      weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_pff, weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_pff,
      weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_pff, weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_pff,
      weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_pff, weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_pff,
      weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_pff, weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_pff,
      weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_pff, weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_pff,
      weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_pff, weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_pff,
      weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_pff, weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_pff,
      weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_pff, weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_pff,
      weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_pff
);
  input clk;
  input rst;
  input start_vld;
  output start_rdy;
  input start_dat;
  input input_port_vld;
  output input_port_rdy;
  input [73:0] input_port_dat;
  input rva_in_vld;
  output rva_in_rdy;
  input [96:0] rva_in_dat;
  output rva_out_vld;
  input rva_out_rdy;
  output [63:0] rva_out_dat;
  output act_port_vld;
  input act_port_rdy;
  output [255:0] act_port_dat;
  input [31:0] SC_SRAM_CONFIG;
  output weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d;
  output [63:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_d_d;
  input [63:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_radr_d;
  output weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d;
  output [63:0] weight_mem_banks_bank_a0_a0_a1_a_rsci_d_d;
  input [63:0] weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a0_a0_a1_a_rsci_radr_d;
  output weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d;
  output [63:0] weight_mem_banks_bank_a0_a1_a0_a_rsci_d_d;
  input [63:0] weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a0_a1_a0_a_rsci_radr_d;
  output weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d;
  output [63:0] weight_mem_banks_bank_a0_a1_a1_a_rsci_d_d;
  input [63:0] weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a0_a1_a1_a_rsci_radr_d;
  output weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d;
  output [63:0] weight_mem_banks_bank_a1_a0_a0_a_rsci_d_d;
  input [63:0] weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a1_a0_a0_a_rsci_radr_d;
  output weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d;
  output [63:0] weight_mem_banks_bank_a1_a0_a1_a_rsci_d_d;
  input [63:0] weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a1_a0_a1_a_rsci_radr_d;
  output weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d;
  output [63:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_d_d;
  input [63:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_radr_d;
  output weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d;
  output [63:0] weight_mem_banks_bank_a1_a1_a1_a_rsci_d_d;
  input [63:0] weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d;
  output [11:0] weight_mem_banks_bank_a1_a1_a1_a_rsci_radr_d;
  output [7:0] ProductSum_for_acc_11_cmp_a;
  output ProductSum_for_acc_11_cmp_en;
  input [22:0] ProductSum_for_acc_11_cmp_z;
  output [7:0] ProductSum_for_acc_10_cmp_a;
  input [22:0] ProductSum_for_acc_10_cmp_z;
  output [7:0] ProductSum_for_acc_9_cmp_a0;
  output [7:0] ProductSum_for_acc_9_cmp_b0;
  output [7:0] ProductSum_for_acc_9_cmp_c0;
  output ProductSum_for_acc_9_cmp_en;
  input [22:0] ProductSum_for_acc_9_cmp_z;
  output [7:0] ProductSum_for_acc_8_cmp_a0;
  output [7:0] ProductSum_for_acc_8_cmp_b0;
  output [7:0] ProductSum_for_acc_8_cmp_c0;
  input [22:0] ProductSum_for_acc_8_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_a;
  input [22:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_4_cmp_a;
  input [22:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_4_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_c0;
  input [22:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_c0;
  input [22:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_a;
  input [22:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_4_cmp_a;
  input [22:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_4_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_c0;
  input [22:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_c0;
  input [22:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_a;
  input [22:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_4_cmp_a;
  input [22:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_4_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_c0;
  input [22:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_c0;
  input [22:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_a;
  input [22:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_4_cmp_a;
  input [22:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_4_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_c0;
  input [22:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_c0;
  input [22:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_a;
  output PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_load;
  input [22:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_a;
  output [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_b;
  input [22:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_c0;
  input [22:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_c0;
  input [22:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_a;
  input [22:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_4_cmp_a;
  input [22:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_4_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_c0;
  input [22:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_c0;
  input [22:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_a;
  input [22:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_a;
  input [22:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_c0;
  input [22:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_z;
  output [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_a0;
  output [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_b0;
  output [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_c0;
  input [22:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_z;
  output [7:0] ProductSum_for_acc_11_cmp_b_pff;
  output ProductSum_for_acc_11_cmp_load_pff;
  output ProductSum_for_acc_11_cmp_datavalid_pff;
  output [7:0] ProductSum_for_acc_10_cmp_b_pff;
  output [7:0] ProductSum_for_acc_9_cmp_a1_pff;
  output [7:0] ProductSum_for_acc_9_cmp_b1_pff;
  output [7:0] ProductSum_for_acc_9_cmp_c1_pff;
  output ProductSum_for_acc_9_cmp_load_pff;
  output ProductSum_for_acc_9_cmp_datavalid_pff;
  output [7:0] ProductSum_for_acc_8_cmp_a1_pff;
  output [7:0] ProductSum_for_acc_8_cmp_b1_pff;
  output [7:0] ProductSum_for_acc_8_cmp_c1_pff;
  output PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_load_pff;
  output PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_load_pff;
  output PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_load_pff;
  output PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_load_pff;
  output PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_load_pff;
  output PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_load_pff;
  output PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_load_pff;
  output PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_load_pff;
  output PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_load_pff;
  output PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_load_pff;
  output PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_load_pff;
  output PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_load_pff;
  output PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_load_pff;
  output weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_pff;
  output [11:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_pff;
  output weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_pff;
  output weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_pff;
  output weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_pff;
  output weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_pff;
  output weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_pff;
  output weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_pff;
  output weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_pff;
  output weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_pff;
  output weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_pff;
  output weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_pff;
  output weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_pff;
  output weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_pff;
  output [11:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_pff;
  output weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_pff;
  output weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_pff;
  output weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_pff;


  // Interconnect Declarations
  wire PECoreRun_wen;
  wire PECoreRun_wten;
  wire [63:0] rva_in_PopNB_mioi_data_data_rsc_z_mxwt;
  wire [19:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt;
  wire rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  wire rva_in_PopNB_mioi_return_rsc_z_mxwt;
  wire [63:0] input_port_PopNB_mioi_data_data_data_rsc_z_mxwt;
  wire [7:0] input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt;
  wire input_port_PopNB_mioi_return_rsc_z_mxwt;
  wire act_port_Push_mioi_wen_comp;
  wire start_PopNB_mioi_data_rsc_z_mxwt;
  wire start_PopNB_mioi_return_rsc_z_mxwt;
  wire rva_out_Push_mioi_wen_comp;
  wire [10:0] PEManager_15U_GetWeightAddr_else_acc_4_cmp_z;
  wire fsm_output;
  wire pe_config_UpdateManagerCounter_if_if_unequal_tmp;
  wire [7:0] weight_mem_write_arbxbar_xbar_for_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_for_1_lshift_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_3_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_1_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp;
  wire [7:0] weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp;
  wire while_mux_1298_tmp;
  wire while_mux_1285_tmp;
  wire while_mux_1283_tmp;
  wire while_mux_1282_tmp;
  wire while_mux_1281_tmp;
  wire while_mux_1280_tmp;
  wire while_mux_1279_tmp;
  wire while_mux_1278_tmp;
  wire while_mux_1277_tmp;
  wire while_mux_1276_tmp;
  wire while_mux_1275_tmp;
  wire while_mux_1274_tmp;
  wire while_mux_1273_tmp;
  wire while_mux_1272_tmp;
  wire while_mux_1271_tmp;
  wire while_mux_1270_tmp;
  wire while_mux_1269_tmp;
  wire while_mux_1268_tmp;
  wire while_mux_1267_tmp;
  wire while_mux_1266_tmp;
  wire while_mux_1265_tmp;
  wire while_mux_1264_tmp;
  wire while_mux_1263_tmp;
  wire while_mux_1262_tmp;
  wire while_mux_1261_tmp;
  wire while_mux_1260_tmp;
  wire while_mux_1259_tmp;
  wire while_mux_1258_tmp;
  wire while_mux_1257_tmp;
  wire while_mux_1256_tmp;
  wire while_mux_1251_tmp;
  wire while_mux_1250_tmp;
  wire while_mux_1249_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_124_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_30_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_113_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_112_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_26_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_101_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_100_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_22_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_89_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_88_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_18_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_77_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_76_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_14_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_65_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_64_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_10_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_53_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_52_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_6_tmp;
  wire weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_2_tmp;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_mux_1_tmp;
  wire weight_mem_run_1_if_for_weight_mem_run_1_if_for_weight_mem_run_1_if_for_nor_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_126_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_122_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_114_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_110_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_102_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_98_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_90_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_86_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_78_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_74_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_66_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_62_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_54_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_50_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_42_tmp;
  wire Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_38_tmp;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_tmp;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_and_49_tmp;
  wire PECore_DecodeAxiRead_case_4_switch_lp_nor_6_tmp;
  wire PECore_DecodeAxiRead_case_4_switch_lp_nor_8_tmp;
  wire and_dcpl_4;
  wire and_dcpl_5;
  wire and_dcpl_6;
  wire and_dcpl_27;
  wire and_dcpl_31;
  wire and_dcpl_32;
  wire or_tmp_2;
  wire or_tmp_3;
  wire and_dcpl_40;
  wire and_dcpl_41;
  wire or_tmp_4;
  wire and_tmp;
  wire or_tmp_5;
  wire nor_tmp_1;
  wire and_dcpl_69;
  wire and_dcpl_78;
  wire and_dcpl_79;
  wire and_dcpl_80;
  wire and_dcpl_82;
  wire and_dcpl_84;
  wire and_dcpl_86;
  wire and_dcpl_88;
  wire and_dcpl_90;
  wire and_dcpl_92;
  wire or_dcpl_13;
  wire or_dcpl_16;
  wire or_dcpl_21;
  wire and_dcpl_149;
  wire and_dcpl_150;
  wire and_dcpl_151;
  wire and_dcpl_152;
  wire and_dcpl_153;
  wire and_dcpl_154;
  wire and_dcpl_155;
  wire and_dcpl_156;
  wire and_dcpl_162;
  wire and_dcpl_168;
  wire and_dcpl_178;
  wire and_dcpl_179;
  wire and_dcpl_181;
  wire and_dcpl_182;
  wire and_dcpl_184;
  wire and_dcpl_185;
  wire and_dcpl_187;
  wire and_dcpl_188;
  wire and_dcpl_190;
  wire and_dcpl_191;
  wire and_dcpl_193;
  wire and_dcpl_194;
  wire and_dcpl_196;
  wire and_dcpl_197;
  wire and_dcpl_199;
  wire and_dcpl_200;
  wire and_dcpl_203;
  wire and_dcpl_204;
  wire and_dcpl_207;
  wire and_dcpl_209;
  wire or_dcpl_87;
  wire and_dcpl_210;
  wire or_dcpl_91;
  wire and_dcpl_211;
  wire and_dcpl_215;
  wire and_dcpl_216;
  wire and_dcpl_217;
  wire and_dcpl_219;
  wire and_dcpl_221;
  wire or_tmp_33;
  wire and_dcpl_228;
  wire and_dcpl_241;
  wire and_dcpl_242;
  wire and_dcpl_246;
  wire and_dcpl_248;
  wire and_dcpl_266;
  wire mux_tmp_25;
  wire or_tmp_43;
  wire and_dcpl_281;
  wire and_dcpl_282;
  wire and_dcpl_293;
  wire and_dcpl_294;
  wire or_tmp_206;
  wire not_tmp_203;
  wire or_tmp_215;
  wire mux_tmp_108;
  wire and_dcpl_312;
  wire not_tmp_217;
  wire and_dcpl_329;
  wire and_dcpl_355;
  wire and_dcpl_376;
  wire or_tmp_334;
  wire and_dcpl_389;
  wire and_dcpl_398;
  wire and_dcpl_401;
  wire and_dcpl_419;
  wire and_dcpl_420;
  wire mux_tmp_182;
  wire and_dcpl_431;
  wire and_dcpl_459;
  wire and_dcpl_467;
  wire or_tmp_341;
  wire or_tmp_342;
  wire and_dcpl_469;
  wire or_tmp_347;
  wire not_tmp_312;
  wire or_tmp_352;
  wire not_tmp_314;
  wire or_tmp_358;
  wire not_tmp_316;
  wire or_tmp_364;
  wire or_tmp_365;
  wire not_tmp_319;
  wire not_tmp_322;
  wire not_tmp_325;
  wire or_tmp_382;
  wire or_dcpl_603;
  wire and_dcpl_504;
  wire and_dcpl_505;
  wire or_dcpl_606;
  wire and_dcpl_525;
  wire or_dcpl_615;
  wire and_dcpl_529;
  wire and_dcpl_532;
  wire and_dcpl_533;
  wire and_dcpl_543;
  wire and_dcpl_547;
  wire and_dcpl_550;
  wire and_dcpl_554;
  wire and_dcpl_557;
  wire and_dcpl_561;
  wire and_dcpl_564;
  wire and_dcpl_568;
  wire or_dcpl_616;
  wire or_dcpl_627;
  wire or_dcpl_628;
  wire or_dcpl_632;
  wire or_dcpl_635;
  wire or_dcpl_658;
  wire and_dcpl_580;
  wire and_dcpl_582;
  wire and_dcpl_584;
  wire and_dcpl_588;
  wire and_dcpl_592;
  wire or_dcpl_665;
  wire and_dcpl_611;
  wire and_dcpl_612;
  wire and_dcpl_616;
  wire nor_tmp_39;
  wire or_tmp_415;
  wire nor_tmp_41;
  wire mux_tmp_277;
  wire mux_tmp_280;
  wire mux_tmp_283;
  wire not_tmp_469;
  wire or_tmp_427;
  wire or_tmp_430;
  wire or_tmp_432;
  wire mux_tmp_293;
  wire mux_tmp_294;
  wire mux_tmp_295;
  wire or_tmp_443;
  wire or_tmp_451;
  wire mux_tmp_305;
  wire or_tmp_458;
  wire and_dcpl_625;
  wire or_tmp_465;
  wire mux_tmp_313;
  wire mux_tmp_314;
  wire mux_tmp_319;
  wire nor_tmp_89;
  wire or_tmp_472;
  wire or_tmp_473;
  wire or_tmp_474;
  wire or_tmp_476;
  wire mux_tmp_320;
  wire nor_tmp_95;
  wire or_tmp_478;
  wire or_tmp_479;
  wire or_tmp_480;
  wire mux_tmp_321;
  wire or_tmp_486;
  wire or_tmp_487;
  wire mux_tmp_327;
  wire or_tmp_489;
  wire mux_tmp_328;
  wire mux_tmp_330;
  wire mux_tmp_332;
  wire mux_tmp_333;
  wire mux_tmp_342;
  wire and_dcpl_626;
  wire or_dcpl_677;
  wire or_tmp_511;
  wire mux_tmp_353;
  wire or_tmp_517;
  wire and_dcpl_629;
  wire and_dcpl_631;
  wire or_tmp_521;
  wire mux_tmp_359;
  wire or_tmp_526;
  wire mux_tmp_360;
  wire mux_tmp_361;
  wire mux_tmp_362;
  wire and_dcpl_632;
  wire and_dcpl_639;
  wire or_tmp_528;
  wire or_tmp_530;
  wire mux_tmp_366;
  wire nor_tmp_123;
  wire or_tmp_532;
  wire or_tmp_533;
  wire or_tmp_534;
  wire or_tmp_536;
  wire nor_tmp_129;
  wire or_tmp_538;
  wire or_tmp_539;
  wire or_tmp_540;
  wire or_tmp_542;
  wire or_tmp_544;
  wire or_tmp_545;
  wire or_tmp_547;
  wire or_tmp_548;
  wire mux_tmp_370;
  wire mux_tmp_371;
  wire and_dcpl_641;
  wire or_tmp_564;
  wire or_tmp_566;
  wire mux_tmp_387;
  wire nor_tmp_143;
  wire or_tmp_568;
  wire or_tmp_569;
  wire or_tmp_570;
  wire or_tmp_572;
  wire nor_tmp_149;
  wire or_tmp_574;
  wire or_tmp_575;
  wire or_tmp_576;
  wire or_tmp_578;
  wire or_tmp_580;
  wire or_tmp_581;
  wire or_tmp_583;
  wire or_tmp_584;
  wire mux_tmp_391;
  wire mux_tmp_392;
  wire and_dcpl_642;
  wire or_tmp_600;
  wire or_tmp_602;
  wire mux_tmp_408;
  wire nor_tmp_163;
  wire or_tmp_604;
  wire or_tmp_605;
  wire or_tmp_606;
  wire or_tmp_608;
  wire nor_tmp_169;
  wire or_tmp_610;
  wire or_tmp_611;
  wire or_tmp_612;
  wire or_tmp_614;
  wire or_tmp_616;
  wire or_tmp_617;
  wire or_tmp_619;
  wire or_tmp_620;
  wire mux_tmp_412;
  wire mux_tmp_413;
  wire and_dcpl_643;
  wire or_tmp_636;
  wire or_tmp_638;
  wire mux_tmp_429;
  wire or_tmp_642;
  wire or_tmp_644;
  wire or_tmp_648;
  wire or_tmp_650;
  wire or_tmp_652;
  wire or_tmp_653;
  wire or_tmp_655;
  wire or_tmp_656;
  wire mux_tmp_435;
  wire mux_tmp_436;
  wire or_tmp_665;
  wire or_tmp_668;
  wire and_dcpl_644;
  wire or_tmp_678;
  wire or_tmp_680;
  wire mux_tmp_454;
  wire or_tmp_685;
  wire or_tmp_690;
  wire and_dcpl_645;
  wire or_tmp_692;
  wire or_tmp_693;
  wire or_tmp_694;
  wire or_tmp_696;
  wire or_tmp_697;
  wire or_tmp_698;
  wire mux_tmp_458;
  wire mux_tmp_459;
  wire and_dcpl_646;
  wire and_dcpl_651;
  wire or_dcpl_678;
  wire while_and_24_cse;
  wire [3:0] pe_config_manager_counter_sva_mx1;
  wire [4:0] operator_4_false_acc_sdt_sva_1;
  wire [5:0] nl_operator_4_false_acc_sdt_sva_1;
  reg [3:0] pe_config_num_manager_sva;
  wire state_0_sva_mx1;
  wire while_if_and_tmp_1;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  wire PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_nor_1_cse_1;
  reg PECore_DecodeAxiWrite_switch_lp_equal_tmp_1;
  reg PECore_DecodeAxiWrite_switch_lp_equal_tmp_2;
  reg PECore_DecodeAxiWrite_switch_lp_nor_tmp_1;
  reg pe_config_is_valid_sva;
  reg pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_nor_mdf_sva_st_1;
  wire pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_if_nor_mdf_sva_1;
  reg pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1;
  reg PECore_UpdateFSM_switch_lp_and_7_itm_1;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_1;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_3_1;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_5_1;
  reg PECore_UpdateFSM_switch_lp_nor_7_itm_1;
  reg [8:0] operator_8_false_acc_sdt_sva_1;
  wire [9:0] nl_operator_8_false_acc_sdt_sva_1;
  wire PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva_mx1;
  wire PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_cse_1;
  wire PECore_RunFSM_switch_lp_equal_tmp_1_mx0w1;
  reg PECore_RunFSM_switch_lp_nor_tmp_1;
  reg [1:0] state_2_1_sva;
  reg state_0_sva;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_11_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_10_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_14_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_13_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_12_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_9_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_7_1_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_7_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_7_4_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_7_2_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_7_5_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_7_6_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_7_7_sva_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_7_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_7_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_11_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_10_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_14_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_13_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_12_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_9_7_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_6_1_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_6_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_6_4_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_6_2_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_6_5_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_6_6_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_6_7_sva_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_6_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_6_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_11_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_13_6_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_5_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_5_4_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_5_6_sva_mx1;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_5_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_5_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_11_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_10_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_14_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_13_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_12_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_9_5_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_4_1_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_4_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_4_4_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_4_2_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_4_5_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_4_6_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_4_7_sva_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_4_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_4_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_11_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_10_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_14_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_13_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_12_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_9_4_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_3_1_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_3_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_3_4_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_3_2_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_3_5_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_3_6_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_3_7_sva_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_3_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_3_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_11_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_10_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_14_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_13_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_12_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_9_3_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_2_1_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_2_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_2_4_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_2_2_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_2_5_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_2_6_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_2_7_sva_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_2_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_2_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_11_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_10_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_14_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_13_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_12_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_9_2_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_1_1_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_1_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_1_4_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_1_2_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_1_5_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_1_6_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_1_7_sva_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_1_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_1_lpi_1_dfm_mx0;
  wire Arbiter_8U_Roundrobin_pick_1_priority_14_1_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_priority_13_1_sva_1;
  wire weight_mem_read_arbxbar_arbiters_next_0_2_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_0_5_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_0_6_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_0_7_sva_mx0;
  reg PECore_RunFSM_switch_lp_equal_tmp_1_2;
  reg weight_mem_run_3_for_land_lpi_1_dfm_2;
  reg weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  reg weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  reg weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  reg weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  reg weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  wire weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_3_m1c_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  reg weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  reg weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  reg weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  reg input_read_req_valid_lpi_1_dfm_1_9;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7;
  reg rva_in_reg_rw_sva_9;
  wire PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_m1c_1;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_9;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_9;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_9;
  wire PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_and_5;
  wire PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0;
  wire PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0;
  wire PECore_UpdateFSM_switch_lp_equal_tmp_6;
  wire PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_1_cse_1;
  wire PECore_RunScale_PECore_RunScale_if_and_1_svs_1;
  wire PECore_UpdateFSM_switch_lp_nor_tmp_1;
  wire PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_1_cse_1;
  wire [7:0] pe_config_input_counter_sva_mx1;
  wire [8:0] operator_16_false_acc_sdt_sva_1;
  wire [9:0] nl_operator_16_false_acc_sdt_sva_1;
  reg [7:0] pe_manager_num_input_sva;
  reg [7:0] pe_config_num_output_sva;
  wire PECore_PushOutput_PECore_PushOutput_if_and_svs_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_5_1;
  wire Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_3_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_2_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_6_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_15;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_15;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_15;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_15;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_5_1;
  wire Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_2_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_3_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_6_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_14;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_14;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_14;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_14;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_3_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_6_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_5_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_13;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_13;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_13;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_13;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1;
  wire Arbiter_8U_Roundrobin_pick_1_unequal_tmp_15;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_8;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_8;
  reg weight_mem_run_3_for_land_lpi_1_dfm_1;
  reg weight_mem_run_3_for_land_6_lpi_1_dfm_1;
  reg weight_mem_run_3_for_land_4_lpi_1_dfm_1;
  reg weight_mem_run_3_for_land_2_lpi_1_dfm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3;
  wire PECore_DecodeAxiWrite_switch_lp_nor_tmp_1_1;
  wire PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_mx0w0;
  reg PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_1_1;
  wire weight_mem_run_3_for_land_lpi_1_dfm_1_1;
  wire weight_mem_run_3_for_land_6_lpi_1_dfm_1_1;
  reg pe_manager_base_weight_slc_pe_manager_base_weight_2_0_178_itm_1;
  reg weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  wire weight_mem_run_3_for_land_4_lpi_1_dfm_1_1;
  wire weight_mem_run_3_for_land_2_lpi_1_dfm_1_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_6_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_6_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_4_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_4_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4_1;
  wire Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4_1;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_6;
  reg Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_4;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_0_2_lpi_1_dfm_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_2;
  wire Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_2;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_0_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_0_1;
  wire Arbiter_8U_Roundrobin_pick_1_unequal_tmp_10;
  wire Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11;
  wire Arbiter_8U_Roundrobin_pick_1_unequal_tmp_12;
  wire Arbiter_8U_Roundrobin_pick_1_unequal_tmp_13;
  wire Arbiter_8U_Roundrobin_pick_1_unequal_tmp_14;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_8;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_8;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1;
  reg pe_manager_base_weight_slc_pe_manager_base_weight_2_0_95_itm_1;
  reg pe_manager_base_weight_slc_pe_manager_base_weight_2_0_93_itm_1;
  reg pe_manager_base_weight_slc_pe_manager_base_weight_2_0_122_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_1_itm_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1_1;
  wire weight_mem_run_3_for_land_1_lpi_1_dfm_1_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_11_itm_1;
  reg rva_in_reg_rw_sva_5;
  wire PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_127_sva_1;
  reg input_write_req_valid_lpi_1_dfm_1_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_127_sva_1;
  wire input_write_req_valid_lpi_1_dfm_5;
  wire input_mem_banks_write_if_for_if_and_stg_6_126_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_126_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_125_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_125_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_124_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_124_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_123_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_123_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_122_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_122_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_121_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_121_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_120_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_120_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_119_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_119_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_118_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_118_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_117_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_117_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_116_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_116_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_115_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_115_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_114_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_114_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_113_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_113_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_112_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_112_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_111_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_111_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_110_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_110_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_109_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_109_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_108_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_108_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_107_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_107_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_106_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_106_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_105_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_105_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_104_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_104_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_103_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_103_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_102_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_102_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_101_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_101_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_100_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_100_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_99_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_99_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_98_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_98_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_97_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_97_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_96_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_96_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_95_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_95_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_94_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_94_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_93_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_93_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_92_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_92_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_91_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_91_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_90_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_90_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_89_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_89_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_88_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_88_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_87_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_87_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_86_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_86_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_85_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_85_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_84_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_84_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_83_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_83_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_82_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_82_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_81_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_81_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_80_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_80_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_79_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_79_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_78_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_78_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_77_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_77_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_76_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_76_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_75_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_75_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_74_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_74_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_73_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_73_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_72_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_72_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_71_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_71_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_70_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_70_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_69_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_69_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_68_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_68_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_67_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_67_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_66_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_66_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_65_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_65_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_64_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_64_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_63_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_63_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_62_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_62_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_61_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_61_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_60_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_60_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_59_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_59_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_58_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_58_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_57_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_57_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_56_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_56_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_55_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_55_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_54_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_54_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_53_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_53_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_52_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_52_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_51_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_51_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_50_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_50_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_49_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_49_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_48_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_48_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_47_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_47_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_46_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_46_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_45_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_45_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_44_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_44_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_43_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_43_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_42_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_42_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_41_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_41_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_40_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_40_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_39_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_39_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_38_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_38_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_37_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_37_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_36_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_36_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_35_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_35_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_34_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_34_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_33_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_33_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_32_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_32_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_31_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_31_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_30_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_30_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_29_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_29_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_28_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_28_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_27_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_27_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_26_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_26_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_25_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_25_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_24_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_24_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_23_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_23_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_22_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_22_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_21_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_21_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_20_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_20_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_19_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_19_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_18_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_18_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_17_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_17_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_16_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_16_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_15_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_15_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_14_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_14_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_13_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_13_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_12_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_12_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_11_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_11_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_10_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_10_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_9_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_9_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_8_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_8_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_7_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_7_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_6_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_6_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_5_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_5_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_4_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_4_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_3_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_3_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_2_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_2_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_1_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_1_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_6_0_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_6_0_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_0_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_1_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_2_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_3_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_4_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_5_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_6_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_7_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_8_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_9_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_10_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_11_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_12_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_13_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_14_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_15_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_16_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_17_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_18_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_19_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_20_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_21_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_22_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_23_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_24_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_25_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_26_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_27_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_28_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_29_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_30_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_31_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_32_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_33_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_34_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_35_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_36_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_37_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_38_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_39_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_40_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_41_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_42_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_43_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_44_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_45_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_46_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_47_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_48_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_49_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_50_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_51_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_52_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_53_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_54_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_55_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_56_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_57_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_58_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_59_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_60_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_61_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_62_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_5_63_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_0_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_1_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_2_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_3_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_4_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_5_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_6_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_7_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_8_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_9_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_10_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_11_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_12_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_13_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_14_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_15_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_16_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_17_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_18_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_19_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_20_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_21_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_22_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_23_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_24_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_25_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_26_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_27_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_28_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_29_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_30_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_4_31_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_0_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_1_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_2_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_3_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_4_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_5_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_6_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_7_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_8_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_9_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_10_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_11_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_12_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_13_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_14_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_3_15_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_0_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_1_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_2_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_3_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_4_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_5_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_6_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_2_7_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_1_0_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_1_1_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_1_2_sva_1;
  wire input_mem_banks_write_if_for_if_and_stg_1_3_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_0_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_1_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_2_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_3_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_4_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_5_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_6_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_7_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_8_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_9_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_10_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_11_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_12_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_13_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_14_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_15_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_16_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_17_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_18_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_19_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_20_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_21_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_22_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_23_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_24_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_25_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_26_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_27_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_28_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_29_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_30_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_31_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_32_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_33_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_34_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_35_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_36_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_37_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_38_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_39_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_40_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_41_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_42_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_43_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_44_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_45_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_46_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_47_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_48_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_49_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_50_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_51_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_52_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_53_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_54_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_55_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_56_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_57_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_58_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_59_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_60_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_61_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_62_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_5_63_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_0_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_1_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_2_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_3_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_4_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_5_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_6_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_7_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_8_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_9_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_10_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_11_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_12_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_13_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_14_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_15_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_16_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_17_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_18_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_19_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_20_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_21_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_22_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_23_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_24_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_25_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_26_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_27_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_28_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_29_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_30_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_4_31_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_0_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_1_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_2_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_3_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_4_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_5_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_6_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_7_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_8_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_9_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_10_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_11_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_12_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_13_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_14_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_3_15_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_0_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_1_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_2_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_3_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_4_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_5_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_6_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_2_7_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_1_0_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_1_1_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_1_2_sva_1;
  wire input_mem_banks_write_1_if_for_if_and_stg_1_3_sva_1;
  reg [14:0] pe_manager_base_input_sva;
  reg PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_2;
  wire PECore_DecodeAxiRead_switch_lp_equal_tmp_4;
  wire PECore_DecodeAxiRead_switch_lp_nor_tmp_mx0w0;
  wire PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_mx0w0;
  reg accum_vector_data_7_sva_1_load;
  reg accum_vector_data_6_sva_1_load;
  reg accum_vector_data_5_sva_1_load;
  reg accum_vector_data_4_sva_1_load;
  reg accum_vector_data_3_sva_1_load;
  reg accum_vector_data_2_sva_1_load;
  reg accum_vector_data_1_sva_1_load;
  reg accum_vector_data_0_sva_1_load;
  reg rva_in_reg_rw_sva_st_1_9;
  reg input_read_req_valid_lpi_1_dfm_1_8;
  reg rva_in_reg_rw_sva_8;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6;
  reg rva_in_reg_rw_sva_st_1_8;
  reg rva_in_reg_rw_sva_st_8;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_8;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_8;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_8;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_7;
  reg while_stage_0_10;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_8;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_8;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7;
  reg rva_in_reg_rw_sva_st_1_6;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_st_5;
  reg weight_mem_run_3_for_land_3_lpi_1_dfm_2;
  reg while_stage_0_7;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4;
  reg rva_in_reg_rw_sva_st_1_5;
  reg rva_in_reg_rw_sva_st_5;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_5;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_5;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_5;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_44_itm_1;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4;
  reg while_stage_0_6;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_54_itm_1;
  reg weight_mem_run_3_for_land_3_lpi_1_dfm_1;
  reg weight_mem_run_3_for_land_5_lpi_1_dfm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_78_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_1;
  reg weight_mem_run_3_for_land_7_lpi_1_dfm_1;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3;
  reg rva_in_reg_rw_sva_st_1_4;
  reg weight_mem_run_3_for_land_1_lpi_1_dfm_2;
  reg weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  reg while_stage_0_5;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_44_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_76_itm_1;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_3;
  reg ProductSum_for_asn_16_itm_3;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_st_3;
  reg ProductSum_for_asn_25_itm_3;
  reg ProductSum_for_asn_42_itm_3;
  reg ProductSum_for_asn_51_itm_3;
  reg ProductSum_for_asn_64_itm_3;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_1;
  reg ProductSum_for_asn_73_itm_3;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_1;
  reg while_stage_0_4;
  reg while_stage_0_3;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2;
  reg PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5;
  reg while_stage_0_9;
  reg rva_in_reg_rw_sva_st_1_7;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_7;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_st_7;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_st_7;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_st_6;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_6;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_st_6;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_st_5;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_5;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_st_3;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_3;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_st_2;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_1_1;
  reg while_stage_0_8;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_46_itm_1;
  reg rva_in_reg_rw_sva_st_7;
  reg input_read_req_valid_lpi_1_dfm_1_7;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_6;
  reg rva_in_reg_rw_sva_7;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_3;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_3;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_7;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_7;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_7;
  reg accum_vector_operator_1_for_asn_70_itm_6;
  reg accum_vector_operator_1_for_asn_61_itm_6;
  reg accum_vector_operator_1_for_asn_52_itm_6;
  reg accum_vector_operator_1_for_asn_43_itm_6;
  reg accum_vector_operator_1_for_asn_34_itm_6;
  reg accum_vector_operator_1_for_asn_25_itm_6;
  reg accum_vector_operator_1_for_asn_16_itm_6;
  reg accum_vector_operator_1_for_asn_7_itm_6;
  reg input_read_req_valid_lpi_1_dfm_1_6;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_4;
  reg rva_in_reg_rw_sva_4;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_17_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_95_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_86_itm_1;
  reg [2:0] crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_1;
  reg rva_in_reg_rw_sva_st_4;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_4;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_4;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_4;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2;
  reg rva_in_reg_rw_sva_st_6;
  reg PECore_RunMac_PECore_RunMac_if_and_svs_st_2;
  reg rva_in_reg_rw_sva_6;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_5;
  reg accum_vector_operator_1_for_asn_7_itm_1;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_6;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_6;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_6;
  reg ProductSum_for_asn_64_itm_1;
  reg rva_in_reg_rw_sva_st_3;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_2;
  reg rva_in_reg_rw_sva_3;
  reg input_read_req_valid_lpi_1_dfm_1_3;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_5;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_3;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2_3;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_3;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_1;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3_2;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_2;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_2;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_3;
  reg PECore_DecodeAxiRead_switch_lp_nor_tmp_1;
  reg [3:0] while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_1;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_3;
  reg weight_mem_run_3_for_5_and_108_itm_1;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_3;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_7_itm_1;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_1;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_20_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_19_itm_1;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_3;
  reg [1:0] state_2_1_sva_dfm_1;
  reg while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_9;
  reg while_stage_0_11;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_9;
  reg weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  reg weight_mem_run_3_for_land_3_lpi_1_dfm_3;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_2;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_2;
  reg PECore_RunScale_PECore_RunScale_if_and_1_svs_8;
  reg weight_mem_run_3_for_land_7_lpi_1_dfm_2;
  reg weight_mem_run_3_for_land_5_lpi_1_dfm_2;
  reg while_and_1126_itm_1;
  reg [7:0] weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1;
  reg weight_mem_read_arbxbar_arbiters_next_7_5_sva;
  reg Arbiter_8U_Roundrobin_pick_1_mux_538_itm_1;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_7_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_7_4_sva;
  reg Arbiter_8U_Roundrobin_pick_1_mux_542_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_537_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_541_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_540_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_539_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_6_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_5_sva;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_464_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_465_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_496_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_6_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_6_4_sva;
  reg Arbiter_8U_Roundrobin_pick_1_mux_468_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_469_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_466_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_6_3_sva;
  reg Arbiter_8U_Roundrobin_pick_1_mux_467_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_5_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_4_sva;
  reg Arbiter_8U_Roundrobin_pick_1_mux_394_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_393_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_5_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_5_sva;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_4_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_4_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_5_sva;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_3_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_3_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_5_sva;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_2_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_2_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_5_sva;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_1_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_1_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_4_sva;
  reg weight_mem_read_arbxbar_arbiters_next_1_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_5_sva;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1;
  reg weight_mem_read_arbxbar_arbiters_next_0_6_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_1_sva;
  reg weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs;
  wire operator_7_false_1_operator_7_false_1_or_mdf_sva_1;
  wire operator_7_false_1_operator_7_false_1_or_mdf_7_sva_1;
  wire operator_7_false_1_operator_7_false_1_or_mdf_5_sva_1;
  wire operator_7_false_1_operator_7_false_1_or_mdf_4_sva_1;
  wire operator_7_false_1_operator_7_false_1_or_mdf_3_sva_1;
  wire operator_7_false_1_operator_7_false_1_or_mdf_2_sva_1;
  reg [2:0] weight_read_addrs_7_lpi_1_dfm_3_2_0;
  reg [2:0] weight_read_addrs_5_lpi_1_dfm_3_2_0;
  reg [2:0] weight_read_addrs_3_lpi_1_dfm_3_2_0;
  reg [2:0] weight_read_addrs_7_lpi_1_dfm_2_2_0;
  reg [2:0] weight_read_addrs_5_lpi_1_dfm_2_2_0;
  reg [2:0] weight_read_addrs_3_lpi_1_dfm_2_2_0;
  reg [14:0] weight_read_addrs_7_lpi_1_dfm_1;
  reg [14:0] weight_read_addrs_5_lpi_1_dfm_1;
  reg [14:0] pe_manager_base_weight_sva;
  reg [14:0] weight_read_addrs_3_lpi_1_dfm_1;
  reg [14:0] weight_read_addrs_1_lpi_1_dfm_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112_mx0w0;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97_mx0w0;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82_mx0w0;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67_mx0w0;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52_mx0w0;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37_mx0w0;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22_mx0w0;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7_mx0w0;
  reg Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7;
  wire [10:0] PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1;
  wire [11:0] nl_PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1;
  reg [2:0] crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1;
  wire [2:0] crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1_1;
  reg [3:0] weight_read_addrs_0_3_0_lpi_1_dfm_1_2;
  wire [14:0] pe_manager_base_weight_sva_mx2;
  wire [3:0] pe_manager_base_weight_sva_mx1_3_0;
  reg [7:0] while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4;
  wire [7:0] input_write_addrs_lpi_1_dfm_2;
  wire PECore_UpdateFSM_next_state_0_lpi_1_dfm_4;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_41_mx1w0;
  reg Arbiter_8U_Roundrobin_pick_1_mux_396_itm_1;
  wire while_and_1123_rgt;
  wire weight_mem_banks_read_1_for_mux_cse;
  wire weight_mem_banks_read_1_for_mux_1_cse;
  wire weight_mem_banks_read_1_for_mux_4_cse;
  wire weight_mem_banks_read_1_for_mux_5_cse;
  wire weight_mem_banks_read_1_for_mux_8_cse;
  wire weight_mem_banks_read_1_for_mux_9_cse;
  wire weight_mem_banks_read_1_for_mux_12_cse;
  wire weight_mem_banks_read_1_for_mux_13_cse;
  wire weight_mem_banks_read_1_for_mux_16_cse;
  wire weight_mem_banks_read_1_for_mux_17_cse;
  wire weight_mem_banks_read_1_for_mux_20_cse;
  wire weight_mem_banks_read_1_for_mux_21_cse;
  wire weight_mem_banks_read_1_for_mux_24_cse;
  wire weight_mem_banks_read_1_for_mux_25_cse;
  wire weight_mem_banks_read_1_for_mux_28_cse;
  wire weight_mem_banks_read_1_for_mux_29_cse;
  wire weight_mem_banks_write_if_for_if_mux_8_cse;
  wire weight_mem_banks_write_if_for_if_mux_9_cse;
  wire weight_mem_banks_read_for_mux_cse;
  wire weight_mem_banks_read_for_mux_1_cse;
  wire weight_mem_banks_write_if_for_if_mux_12_cse;
  wire weight_mem_banks_write_if_for_if_mux_13_cse;
  wire weight_mem_banks_read_for_mux_4_cse;
  wire weight_mem_banks_read_for_mux_5_cse;
  wire weight_mem_banks_write_if_for_if_mux_16_cse;
  wire weight_mem_banks_write_if_for_if_mux_17_cse;
  wire weight_mem_banks_read_for_mux_8_cse;
  wire weight_mem_banks_read_for_mux_9_cse;
  wire weight_mem_banks_write_if_for_if_mux_20_cse;
  wire weight_mem_banks_write_if_for_if_mux_21_cse;
  wire weight_mem_banks_read_for_mux_12_cse;
  wire weight_mem_banks_read_for_mux_13_cse;
  wire weight_mem_banks_write_if_for_if_mux_24_cse;
  wire weight_mem_banks_write_if_for_if_mux_25_cse;
  wire weight_mem_banks_read_for_mux_16_cse;
  wire weight_mem_banks_read_for_mux_17_cse;
  wire weight_mem_banks_write_if_for_if_mux_28_cse;
  wire weight_mem_banks_write_if_for_if_mux_29_cse;
  wire weight_mem_banks_read_for_mux_20_cse;
  wire weight_mem_banks_read_for_mux_21_cse;
  wire weight_mem_banks_write_if_for_if_mux_32_cse;
  wire weight_mem_banks_write_if_for_if_mux_33_cse;
  wire weight_mem_banks_read_for_mux_24_cse;
  wire weight_mem_banks_read_for_mux_25_cse;
  wire weight_mem_banks_write_if_for_if_mux_36_cse;
  wire weight_mem_banks_write_if_for_if_mux_37_cse;
  wire weight_mem_banks_read_for_mux_28_cse;
  wire weight_mem_banks_read_for_mux_29_cse;
  wire input_mem_banks_write_1_if_for_if_mux_cse;
  wire input_mem_banks_write_1_if_for_if_mux_1_cse;
  wire input_mem_banks_read_1_for_mux_cse;
  wire input_mem_banks_read_1_for_mux_1_cse;
  wire input_mem_banks_write_if_for_if_mux_cse;
  wire input_mem_banks_write_if_for_if_mux_1_cse;
  wire input_mem_banks_read_for_mux_cse;
  wire input_mem_banks_read_for_mux_1_cse;
  reg reg_PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_cgo_ir_cse;
  reg reg_PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_cse;
  reg reg_weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_cse;
  reg reg_rva_out_Push_mioi_iswt0_cse;
  reg reg_start_PopNB_mioi_iswt0_cse;
  reg reg_act_port_Push_mioi_iswt0_cse;
  reg reg_rva_in_PopNB_mioi_iswt0_cse;
  wire rva_out_reg_data_and_cse;
  wire weight_port_read_out_data_and_1_cse;
  wire weight_port_read_out_data_and_3_cse;
  wire weight_port_read_out_data_and_5_cse;
  wire weight_port_read_out_data_and_8_cse;
  wire weight_port_read_out_data_and_14_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_cse;
  reg reg_rva_in_reg_rw_sva_st_1_1_cse;
  reg [2:0] reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse;
  wire weight_port_read_out_data_and_7_cse;
  wire weight_port_read_out_data_and_60_cse;
  wire operator_15_false_1_and_cse;
  wire pe_config_num_manager_and_cse;
  wire PECore_DecodeAxiWrite_switch_lp_and_cse;
  reg reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse;
  wire or_196_cse;
  wire or_162_cse;
  wire or_186_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_cse;
  wire nor_340_cse;
  reg reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_3_1_itm_2_cse;
  reg reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_2_itm_2_cse;
  wire and_680_cse;
  reg reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_0_1_itm_2_cse;
  reg reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_2_1_itm_2_cse;
  wire pe_manager_num_input_and_cse;
  wire or_999_cse;
  wire Arbiter_8U_Roundrobin_pick_nand_54_cse;
  wire Arbiter_8U_Roundrobin_pick_and_37_cse;
  wire Arbiter_8U_Roundrobin_pick_nand_42_cse;
  wire Arbiter_8U_Roundrobin_pick_and_31_cse;
  wire Arbiter_8U_Roundrobin_pick_nand_30_cse;
  wire Arbiter_8U_Roundrobin_pick_and_25_cse;
  wire Arbiter_8U_Roundrobin_pick_nand_18_cse;
  wire Arbiter_8U_Roundrobin_pick_and_19_cse;
  wire Arbiter_8U_Roundrobin_pick_nand_6_cse;
  wire Arbiter_8U_Roundrobin_pick_and_13_cse;
  wire [1:0] state_mux_1_cse;
  wire and_321_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_or_cse;
  wire and_703_cse;
  wire and_702_cse;
  wire and_700_cse;
  wire and_516_cse;
  wire and_692_cse;
  wire weight_mem_read_arbxbar_xbar_1_for_3_8_for_2_or_cse;
  wire or_362_cse;
  wire nor_464_cse;
  wire while_and_23_cse;
  wire nor_17_cse;
  wire nor_18_cse;
  wire nor_469_cse;
  wire and_704_cse;
  wire and_149_cse;
  wire nor_227_cse;
  wire nor_230_cse;
  wire nor_231_cse;
  wire nor_228_cse;
  wire nor_229_cse;
  wire and_114_cse;
  wire nor_238_cse;
  wire nor_239_cse;
  wire nor_236_cse;
  wire nor_237_cse;
  wire nor_242_cse;
  wire nor_243_cse;
  wire nor_240_cse;
  wire nor_241_cse;
  wire nor_246_cse;
  wire nor_247_cse;
  wire nor_244_cse;
  wire nor_245_cse;
  wire nor_250_cse;
  wire nor_251_cse;
  wire nor_248_cse;
  wire nor_249_cse;
  wire nand_36_cse;
  wire while_while_nor_259_cse;
  wire nand_27_cse;
  wire and_714_cse;
  wire and_716_cse;
  wire and_720_cse;
  wire and_721_cse;
  wire and_722_cse;
  wire and_728_cse;
  wire and_729_cse;
  wire and_730_cse;
  wire and_732_cse;
  wire and_737_cse;
  wire and_755_cse;
  wire and_757_cse;
  wire and_756_cse;
  wire and_758_cse;
  wire and_775_cse;
  wire and_776_cse;
  wire and_777_cse;
  wire and_778_cse;
  wire and_779_cse;
  wire and_780_cse;
  wire and_781_cse;
  wire and_789_cse;
  wire and_791_cse;
  wire and_790_cse;
  wire and_792_cse;
  wire and_809_cse;
  wire and_811_cse;
  wire and_810_cse;
  wire and_812_cse;
  wire and_829_cse;
  wire and_831_cse;
  wire and_830_cse;
  wire and_832_cse;
  wire and_855_cse;
  wire and_849_cse;
  wire and_861_cse;
  wire and_851_cse;
  wire and_850_cse;
  wire and_852_cse;
  wire and_853_cse;
  wire and_859_cse;
  wire and_873_cse;
  wire and_874_cse;
  wire and_875_cse;
  wire and_876_cse;
  wire and_879_cse;
  wire and_880_cse;
  wire and_883_cse;
  wire and_884_cse;
  reg Arbiter_8U_Roundrobin_pick_1_mux_31_itm_1;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_6_mx1w0;
  reg Arbiter_8U_Roundrobin_pick_1_mux_30_itm_1;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_5_mx1w0;
  reg accum_vector_operator_1_for_asn_70_itm_5;
  reg accum_vector_operator_1_for_asn_70_itm_4;
  reg accum_vector_operator_1_for_asn_70_itm_3;
  reg accum_vector_operator_1_for_asn_70_itm_2;
  reg accum_vector_operator_1_for_asn_70_itm_1;
  reg accum_vector_operator_1_for_asn_61_itm_5;
  reg accum_vector_operator_1_for_asn_61_itm_4;
  reg accum_vector_operator_1_for_asn_61_itm_3;
  reg accum_vector_operator_1_for_asn_61_itm_2;
  reg PECore_DecodeAxiWrite_switch_lp_equal_tmp_1_2;
  reg accum_vector_operator_1_for_asn_52_itm_5;
  reg accum_vector_operator_1_for_asn_52_itm_4;
  reg accum_vector_operator_1_for_asn_52_itm_3;
  reg accum_vector_operator_1_for_asn_43_itm_5;
  reg accum_vector_operator_1_for_asn_43_itm_4;
  reg accum_vector_operator_1_for_asn_43_itm_3;
  reg accum_vector_operator_1_for_asn_34_itm_5;
  reg accum_vector_operator_1_for_asn_34_itm_4;
  reg accum_vector_operator_1_for_asn_34_itm_3;
  reg accum_vector_operator_1_for_asn_34_itm_2;
  reg accum_vector_operator_1_for_asn_25_itm_5;
  reg accum_vector_operator_1_for_asn_25_itm_4;
  reg accum_vector_operator_1_for_asn_25_itm_3;
  reg accum_vector_operator_1_for_asn_25_itm_2;
  reg accum_vector_operator_1_for_asn_16_itm_5;
  reg accum_vector_operator_1_for_asn_16_itm_4;
  reg accum_vector_operator_1_for_asn_16_itm_3;
  reg accum_vector_operator_1_for_asn_16_itm_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_2;
  reg accum_vector_operator_1_for_asn_7_itm_5;
  reg accum_vector_operator_1_for_asn_7_itm_4;
  reg accum_vector_operator_1_for_asn_7_itm_3;
  wire while_if_and_2_m1c;
  wire PECore_DecodeAxiRead_switch_lp_nor_2_cse;
  wire pe_config_is_valid_and_cse;
  wire weight_mem_run_3_for_5_and_175_cse;
  wire weight_mem_run_3_for_5_and_176_cse;
  wire weight_mem_run_3_for_5_and_177_cse;
  wire weight_mem_run_3_for_5_and_178_cse;
  wire weight_mem_run_3_for_5_and_180_cse;
  wire weight_mem_run_3_for_5_and_181_cse;
  wire Arbiter_8U_Roundrobin_pick_nand_cse;
  wire Arbiter_8U_Roundrobin_pick_and_40_cse;
  wire Arbiter_8U_Roundrobin_pick_nand_69_cse;
  wire Arbiter_8U_Roundrobin_pick_and_52_cse;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_nand_cse;
  wire Arbiter_8U_Roundrobin_pick_and_1_cse;
  wire pe_config_input_counter_and_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_1_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_2_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_cse;
  wire while_and_4_cse;
  wire and_100_cse;
  wire or_1099_cse;
  wire PECore_DecodeAxiWrite_case_4_switch_lp_or_cse_1;
  wire PECore_DecodeAxiWrite_switch_lp_or_5_cse_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_65_cse;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0;
  wire and_514_rmff;
  wire and_510_rmff;
  wire and_506_rmff;
  wire and_502_rmff;
  wire and_498_rmff;
  wire and_494_rmff;
  wire and_490_rmff;
  wire and_487_rmff;
  wire and_483_rmff;
  wire and_480_rmff;
  wire and_518_rmff;
  wire and_520_rmff;
  reg [7:0] pe_config_output_counter_sva;
  reg [7:0] pe_config_input_counter_sva;
  reg rva_out_reg_data_63_sva_dfm_4_4;
  reg [6:0] rva_out_reg_data_62_56_sva_dfm_4_4;
  reg rva_out_reg_data_47_sva_dfm_4_4;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_4_4;
  reg weight_port_read_out_data_slc_weight_port_read_out_data_0_2_0_itm_1;
  reg weight_port_read_out_data_slc_weight_port_read_out_data_0_1_0_itm_1;
  reg weight_port_read_out_data_slc_weight_port_read_out_data_0_0_0_itm_1;
  reg [19:0] act_port_reg_data_243_224_sva_dfm_1_1;
  reg [19:0] act_port_reg_data_211_192_sva_dfm_1_1;
  reg [19:0] act_port_reg_data_179_160_sva_dfm_1_1;
  reg [19:0] act_port_reg_data_147_128_sva_dfm_1_1;
  reg [19:0] act_port_reg_data_115_96_sva_dfm_1_1;
  reg [19:0] act_port_reg_data_83_64_sva_dfm_1_1;
  reg [19:0] act_port_reg_data_51_32_sva_dfm_1_1;
  reg [19:0] act_port_reg_data_19_0_sva_dfm_1_1;
  reg [10:0] weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_11_1;
  reg [10:0] weight_read_addrs_0_14_4_lpi_1_dfm_1_4;
  reg weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_0;
  reg weight_read_addrs_slc_weight_read_addrs_0_3_0_3_23_itm_1;
  reg [10:0] weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_11_1;
  reg weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_0;
  reg weight_read_addrs_4_14_2_lpi_1_dfm_2_0;
  reg [10:0] weight_read_addrs_0_14_4_lpi_1_dfm_1_3;
  reg [13:0] weight_read_addrs_2_14_1_lpi_1_dfm_1;
  reg [12:0] weight_read_addrs_4_14_2_lpi_1_dfm_1;
  reg [13:0] weight_read_addrs_6_14_1_lpi_1_dfm_1;
  reg weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3;
  wire [7:0] weight_port_read_out_data_7_1_sva_dfm_2;
  reg [63:0] input_mem_banks_read_1_read_data_lpi_1_dfm_1_4;
  reg ProductSum_for_asn_16_itm_5;
  wire [7:0] weight_port_read_out_data_7_0_sva_dfm_2;
  reg [7:0] weight_port_read_out_data_7_5_sva_dfm_1;
  reg [47:0] input_mem_banks_read_1_read_data_lpi_1_dfm_1_5_63_16;
  reg [7:0] weight_port_read_out_data_7_2_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_7_3_sva_dfm_1;
  reg ProductSum_for_asn_12_itm_6;
  reg [7:0] weight_port_read_out_data_7_6_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_7_7_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_7_4_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_6_1_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_2_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
  reg ProductSum_for_asn_25_itm_5;
  reg [7:0] weight_port_read_out_data_6_0_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_1_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
  reg [7:0] weight_mem_run_3_for_5_mux_53_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_50_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_51_itm_1;
  reg ProductSum_for_asn_23_itm_6;
  reg [7:0] weight_mem_run_3_for_5_mux_54_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_55_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_52_itm_1;
  wire [7:0] weight_port_read_out_data_5_1_sva_dfm_2;
  reg ProductSum_for_asn_42_itm_5;
  wire [7:0] weight_port_read_out_data_5_0_sva_dfm_2;
  reg [7:0] weight_port_read_out_data_5_5_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_5_2_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_5_3_sva_dfm_1;
  reg ProductSum_for_asn_38_itm_6;
  reg [7:0] weight_port_read_out_data_5_6_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_5_7_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_5_4_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_4_1_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_2_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
  reg ProductSum_for_asn_51_itm_5;
  reg [7:0] weight_port_read_out_data_4_0_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_1_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
  reg [7:0] weight_mem_run_3_for_5_mux_37_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_34_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_35_itm_1;
  reg ProductSum_for_asn_49_itm_6;
  reg [7:0] weight_mem_run_3_for_5_mux_38_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_39_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_36_itm_1;
  reg [7:0] weight_port_read_out_data_3_1_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000000;
  reg ProductSum_for_asn_64_itm_5;
  reg [7:0] weight_port_read_out_data_3_0_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000001;
  reg [7:0] weight_port_read_out_data_3_5_sva_dfm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_26_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_27_itm_1;
  reg ProductSum_for_asn_62_itm_6;
  reg [7:0] weight_port_read_out_data_3_6_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_3_7_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_3_4_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_2_1_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000000;
  reg ProductSum_for_asn_73_itm_5;
  reg [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000001;
  reg [7:0] weight_port_read_out_data_2_0_sva_dfm_1;
  reg [7:0] input_mem_banks_read_1_read_data_lpi_1_dfm_1_5_7_0;
  reg ProductSum_for_asn_72_itm_6;
  reg [7:0] weight_mem_run_3_for_5_mux_21_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_18_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_19_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_22_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_23_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_20_itm_1;
  reg [7:0] weight_port_read_out_data_1_1_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000000;
  reg ProductSum_for_asn_82_itm_5;
  reg [7:0] weight_port_read_out_data_1_0_sva_dfm_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000001;
  reg [7:0] weight_mem_run_3_for_5_mux_13_itm_1;
  reg ProductSum_for_asn_80_itm_6;
  reg [7:0] weight_mem_run_3_for_5_mux_14_itm_1;
  reg [7:0] weight_mem_run_3_for_5_mux_15_itm_1;
  reg ProductSum_for_asn_98_itm_5;
  reg ProductSum_for_asn_94_itm_6;
  reg [7:0] weight_write_data_data_0_7_lpi_1_dfm_1_2_6;
  reg [7:0] weight_write_data_data_0_6_lpi_1_dfm_1_2_6;
  reg [7:0] weight_write_data_data_0_5_lpi_1_dfm_1_2_6;
  reg [7:0] weight_write_data_data_0_4_lpi_1_dfm_1_2_6;
  reg [7:0] weight_write_data_data_0_3_lpi_1_dfm_1_2_6;
  reg [7:0] weight_write_data_data_0_2_lpi_1_dfm_1_2_6;
  reg [7:0] weight_write_data_data_0_1_lpi_1_dfm_1_2_6;
  reg [7:0] weight_write_data_data_0_0_lpi_1_dfm_1_2_6;
  reg [14:0] weight_write_addrs_lpi_1_dfm_1_2;
  reg [7:0] weight_write_data_data_0_7_lpi_1_dfm_1_3_2;
  reg [7:0] weight_write_data_data_0_6_lpi_1_dfm_1_3_2;
  reg [7:0] weight_write_data_data_0_5_lpi_1_dfm_1_3_2;
  reg [7:0] weight_write_data_data_0_4_lpi_1_dfm_1_3_2;
  reg [7:0] weight_write_data_data_0_3_lpi_1_dfm_1_3_2;
  reg [7:0] weight_write_data_data_0_2_lpi_1_dfm_1_3_2;
  reg [7:0] weight_write_data_data_0_1_lpi_1_dfm_1_3_2;
  reg [7:0] weight_write_data_data_0_0_lpi_1_dfm_1_3_2;
  reg [11:0] weight_write_addrs_lpi_1_dfm_1_3_14_3;
  wire or_dcpl_679;
  wire nor_tmp;
  wire and_dcpl_664;
  wire or_dcpl_683;
  wire and_dcpl_665;
  wire or_dcpl_684;
  reg [63:0] input_mem_banks_read_read_data_lpi_1_dfm_1_4;
  reg [63:0] weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1;
  reg [63:0] weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1;
  reg [63:0] weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1;
  reg [63:0] weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1;
  reg [63:0] weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1;
  wire [63:0] weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0;
  wire [55:0] weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0;
  reg [7:0] weight_mem_write_arbxbar_xbar_for_empty_sva_2;
  reg [1:0] pe_manager_base_weight_slc_pe_manager_base_weight_1_0_1_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_79_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_44_itm_2;
  wire or_1401_tmp;
  wire or_1407_tmp;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_1_4;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_1_4;
  reg [5:0] rva_out_reg_data_30_25_sva_dfm_2;
  reg [6:0] rva_out_reg_data_23_17_sva_dfm_2;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_4;
  wire and_923_cse;
  wire and_924_cse;
  wire and_925_cse;
  wire and_926_cse;
  wire and_927_cse;
  wire and_928_cse;
  wire nor_523_cse;
  wire and_931_cse;
  wire and_932_cse;
  wire and_933_cse;
  wire and_934_cse;
  wire and_935_cse;
  wire and_936_cse;
  wire and_937_cse;
  wire nor_524_cse;
  reg pe_config_is_zero_first_sva;
  reg pe_manager_zero_active_sva;
  wire [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm;
  wire [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm;
  wire mux_188_itm;
  wire mux_230_itm;
  wire mux_306_itm;
  wire mux_330_itm;
  wire mux_343_itm;
  wire mux_373_itm;
  wire mux_380_itm;
  wire mux_394_itm;
  wire mux_401_itm;
  wire mux_415_itm;
  wire mux_422_itm;
  wire mux_438_itm;
  wire mux_445_itm;
  wire mux_461_itm;
  reg weight_mem_read_arbxbar_arbiters_next_5_2_sva;
  reg weight_mem_read_arbxbar_arbiters_next_5_5_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_3_sva;
  reg weight_mem_read_arbxbar_arbiters_next_0_4_sva;
  reg [14:0] pe_manager_base_bias_sva;
  reg pe_config_is_cluster_sva;
  reg pe_config_is_bias_sva;
  reg [3:0] pe_config_manager_counter_sva;
  reg [22:0] accum_vector_data_3_sva;
  wire [23:0] nl_accum_vector_data_3_sva;
  reg [22:0] accum_vector_data_4_sva;
  wire [23:0] nl_accum_vector_data_4_sva;
  reg [22:0] accum_vector_data_2_sva;
  wire [23:0] nl_accum_vector_data_2_sva;
  reg [22:0] accum_vector_data_5_sva;
  wire [23:0] nl_accum_vector_data_5_sva;
  reg [22:0] accum_vector_data_1_sva;
  wire [23:0] nl_accum_vector_data_1_sva;
  reg [22:0] accum_vector_data_6_sva;
  wire [23:0] nl_accum_vector_data_6_sva;
  reg [22:0] accum_vector_data_0_sva;
  wire [23:0] nl_accum_vector_data_0_sva;
  reg [22:0] accum_vector_data_7_sva;
  wire [23:0] nl_accum_vector_data_7_sva;
  reg [19:0] act_port_reg_data_115_96_sva;
  reg [19:0] act_port_reg_data_147_128_sva;
  reg [19:0] act_port_reg_data_83_64_sva;
  reg [19:0] act_port_reg_data_179_160_sva;
  reg [19:0] act_port_reg_data_51_32_sva;
  reg [19:0] act_port_reg_data_211_192_sva;
  reg [19:0] act_port_reg_data_19_0_sva;
  reg [19:0] act_port_reg_data_243_224_sva;
  reg [7:0] BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_8;
  reg [63:0] input_mem_banks_bank_a_0_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_1_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_2_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_3_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_4_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_5_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_6_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_7_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_8_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_9_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_10_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_11_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_12_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_13_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_14_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_15_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_16_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_17_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_18_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_19_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_20_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_21_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_22_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_23_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_24_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_25_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_26_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_27_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_28_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_29_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_30_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_31_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_32_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_33_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_34_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_35_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_36_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_37_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_38_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_39_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_40_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_41_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_42_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_43_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_44_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_45_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_46_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_47_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_48_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_49_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_50_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_51_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_52_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_53_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_54_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_55_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_56_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_57_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_58_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_59_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_60_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_61_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_62_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_63_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_64_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_65_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_66_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_67_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_68_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_69_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_70_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_71_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_72_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_73_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_74_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_75_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_76_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_77_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_78_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_79_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_80_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_81_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_82_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_83_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_84_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_85_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_86_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_87_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_88_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_89_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_90_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_91_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_92_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_93_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_94_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_95_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_96_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_97_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_98_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_99_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_100_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_101_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_102_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_103_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_104_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_105_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_106_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_107_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_108_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_109_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_110_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_111_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_112_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_113_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_114_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_115_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_116_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_117_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_118_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_119_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_120_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_121_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_122_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_123_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_124_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_125_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_126_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_127_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_128_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_129_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_130_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_131_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_132_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_133_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_134_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_135_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_136_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_137_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_138_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_139_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_140_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_141_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_142_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_143_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_144_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_145_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_146_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_147_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_148_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_149_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_150_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_151_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_152_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_153_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_154_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_155_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_156_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_157_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_158_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_159_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_160_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_161_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_162_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_163_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_164_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_165_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_166_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_167_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_168_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_169_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_170_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_171_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_172_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_173_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_174_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_175_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_176_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_177_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_178_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_179_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_180_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_181_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_182_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_183_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_184_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_185_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_186_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_187_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_188_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_189_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_190_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_191_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_192_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_193_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_194_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_195_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_196_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_197_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_198_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_199_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_200_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_201_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_202_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_203_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_204_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_205_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_206_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_207_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_208_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_209_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_210_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_211_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_212_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_213_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_214_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_215_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_216_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_217_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_218_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_219_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_220_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_221_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_222_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_223_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_224_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_225_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_226_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_227_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_228_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_229_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_230_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_231_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_232_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_233_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_234_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_235_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_236_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_237_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_238_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_239_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_240_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_241_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_242_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_243_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_244_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_245_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_246_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_247_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_248_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_249_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_250_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_251_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_252_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_253_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_254_sva_dfm_2;
  reg [63:0] input_mem_banks_bank_a_255_sva_dfm_2;
  reg [7:0] weight_port_read_out_data_1_2_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_1_3_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_1_4_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_1_5_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_1_6_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_1_7_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_2_2_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_2_3_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_2_4_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_2_5_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_2_6_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_2_7_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_3_2_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_3_3_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_3_4_sva_dfm_1_1;
  reg [7:0] weight_port_read_out_data_3_5_sva_dfm_1_1;
  reg [7:0] weight_port_read_out_data_3_6_sva_dfm_1_1;
  reg [7:0] weight_port_read_out_data_3_7_sva_dfm_1_1;
  reg [7:0] weight_port_read_out_data_4_2_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_4_3_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_4_4_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_4_5_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_4_6_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_4_7_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_5_0_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_5_1_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_5_2_sva_dfm_1_1;
  reg [7:0] weight_port_read_out_data_5_3_sva_dfm_1_1;
  reg [7:0] weight_port_read_out_data_5_4_sva_dfm_1_1;
  reg [7:0] weight_port_read_out_data_5_5_sva_dfm_1_1;
  reg [7:0] weight_port_read_out_data_5_6_sva_dfm_1_1;
  reg [7:0] weight_port_read_out_data_5_7_sva_dfm_1_1;
  reg [7:0] weight_port_read_out_data_6_2_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_6_3_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_6_4_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_6_5_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_6_6_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_6_7_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_7_0_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_7_1_sva_dfm_1;
  reg [7:0] weight_port_read_out_data_7_2_sva_dfm_1_1;
  reg [7:0] weight_port_read_out_data_7_3_sva_dfm_1_1;
  reg [7:0] weight_port_read_out_data_7_4_sva_dfm_1_1;
  reg [7:0] weight_port_read_out_data_7_5_sva_dfm_1_1;
  reg [7:0] weight_port_read_out_data_7_6_sva_dfm_1_1;
  reg [7:0] weight_port_read_out_data_7_7_sva_dfm_1_1;
  reg rva_out_reg_data_24_sva_dfm_6;
  reg rva_out_reg_data_31_sva_dfm_6;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_6;
  reg rva_out_reg_data_16_sva_dfm_6;
  reg rva_out_reg_data_8_sva_dfm_6;
  reg rva_out_reg_data_0_sva_dfm_6;
  reg [63:0] weight_mem_banks_read_1_read_data_1_lpi_1_dfm_1;
  reg [63:0] weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1_1;
  reg [63:0] weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1_1;
  reg [63:0] weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1_1;
  reg [63:0] weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1_1;
  reg [63:0] weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1_1;
  reg [63:0] weight_mem_banks_read_1_read_data_7_lpi_1_dfm_1;
  reg [6:0] rva_out_reg_data_62_56_sva_dfm_6;
  reg [22:0] accum_vector_data_7_sva_4;
  reg [22:0] accum_vector_data_7_sva_5;
  reg [22:0] accum_vector_data_7_sva_6;
  reg [22:0] accum_vector_data_7_sva_7;
  reg [22:0] accum_vector_data_6_sva_4;
  reg [22:0] accum_vector_data_6_sva_5;
  reg [22:0] accum_vector_data_6_sva_6;
  reg [22:0] accum_vector_data_6_sva_7;
  reg [22:0] accum_vector_data_5_sva_4;
  reg [22:0] accum_vector_data_5_sva_5;
  reg [22:0] accum_vector_data_5_sva_6;
  reg [22:0] accum_vector_data_5_sva_7;
  reg [22:0] accum_vector_data_4_sva_4;
  reg [22:0] accum_vector_data_4_sva_5;
  reg [22:0] accum_vector_data_4_sva_6;
  reg [22:0] accum_vector_data_4_sva_7;
  reg [22:0] accum_vector_data_3_sva_4;
  reg [22:0] accum_vector_data_3_sva_5;
  reg [22:0] accum_vector_data_3_sva_6;
  reg [22:0] accum_vector_data_3_sva_7;
  reg [22:0] accum_vector_data_2_sva_4;
  reg [22:0] accum_vector_data_2_sva_5;
  reg [22:0] accum_vector_data_2_sva_6;
  reg [22:0] accum_vector_data_2_sva_7;
  reg [22:0] accum_vector_data_1_sva_4;
  reg [22:0] accum_vector_data_1_sva_5;
  reg [22:0] accum_vector_data_1_sva_6;
  reg [22:0] accum_vector_data_1_sva_7;
  reg [22:0] accum_vector_data_0_sva_4;
  reg [22:0] accum_vector_data_0_sva_5;
  reg [22:0] accum_vector_data_0_sva_6;
  reg [22:0] accum_vector_data_0_sva_7;
  reg weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  reg weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2;
  reg PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8;
  reg PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1;
  reg [3:0] pe_config_manager_counter_sva_dfm_3_1;
  reg [7:0] input_read_addrs_sva_1_1;
  wire [8:0] nl_input_read_addrs_sva_1_1;
  reg [6:0] rva_out_reg_data_62_56_sva_dfm_4_1;
  reg [6:0] rva_out_reg_data_62_56_sva_dfm_4_2;
  reg [6:0] rva_out_reg_data_62_56_sva_dfm_4_3;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_4_1;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_4_2;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_4_3;
  reg [63:0] input_mem_banks_read_read_data_sva_1;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_1_2;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_1_3;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_1_4;
  reg [7:0] rva_out_reg_data_55_48_sva_dfm_1_5;
  reg [6:0] rva_out_reg_data_62_56_sva_dfm_1_1;
  reg [6:0] rva_out_reg_data_62_56_sva_dfm_1_2;
  reg [6:0] rva_out_reg_data_62_56_sva_dfm_1_3;
  reg [6:0] rva_out_reg_data_62_56_sva_dfm_1_4;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_1_1;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_1_2;
  reg [6:0] rva_out_reg_data_46_40_sva_dfm_1_3;
  reg [3:0] rva_out_reg_data_39_36_sva_dfm_1_1;
  reg [3:0] rva_out_reg_data_39_36_sva_dfm_1_2;
  reg [3:0] rva_out_reg_data_39_36_sva_dfm_1_3;
  reg [3:0] rva_out_reg_data_39_36_sva_dfm_1_4;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_1_1;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_1_2;
  reg [3:0] rva_out_reg_data_35_32_sva_dfm_1_3;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_1;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_2;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_3;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_7;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_8;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_9;
  reg [6:0] rva_out_reg_data_23_17_sva_dfm_1;
  reg [6:0] rva_out_reg_data_23_17_sva_dfm_5;
  reg [6:0] rva_out_reg_data_23_17_sva_dfm_6;
  reg [6:0] rva_out_reg_data_23_17_sva_dfm_7;
  reg [5:0] rva_out_reg_data_30_25_sva_dfm_1;
  reg [5:0] rva_out_reg_data_30_25_sva_dfm_5;
  reg [5:0] rva_out_reg_data_30_25_sva_dfm_6;
  reg [5:0] rva_out_reg_data_30_25_sva_dfm_7;
  reg [7:0] pe_config_output_counter_sva_dfm_1;
  reg [7:0] pe_config_input_counter_sva_dfm_1;
  reg [63:0] rva_in_reg_data_sva_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1;
  reg [7:0] weight_write_data_data_0_0_lpi_1_dfm_1_1;
  reg [7:0] weight_write_data_data_0_1_lpi_1_dfm_1_1;
  reg [7:0] weight_write_data_data_0_2_lpi_1_dfm_1_1;
  reg [7:0] weight_write_data_data_0_3_lpi_1_dfm_1_1;
  reg [7:0] weight_write_data_data_0_4_lpi_1_dfm_1_1;
  reg [7:0] weight_write_data_data_0_5_lpi_1_dfm_1_1;
  reg [7:0] weight_write_data_data_0_6_lpi_1_dfm_1_1;
  reg [7:0] weight_write_data_data_0_7_lpi_1_dfm_1_1;
  reg [10:0] weight_read_addrs_0_14_4_lpi_1_dfm_1_1;
  reg [10:0] weight_read_addrs_0_14_4_lpi_1_dfm_1_2;
  reg [3:0] weight_read_addrs_0_3_0_lpi_1_dfm_1_1;
  reg [7:0] weight_mem_write_arbxbar_xbar_for_empty_sva_1;
  reg [10:0] PEManager_15U_GetWeightAddr_else_acc_3_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_2_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_1_1;
  reg [63:0] input_mem_banks_read_1_read_data_lpi_1_dfm_1_1;
  reg [63:0] input_mem_banks_read_1_read_data_lpi_1_dfm_1_2;
  reg [63:0] input_mem_banks_read_1_read_data_lpi_1_dfm_1_3;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_4;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_5;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_6;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_7;
  reg PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  reg [14:0] pe_manager_base_weight_sva_dfm_3_1;
  reg [14:0] pe_manager_base_input_sva_dfm_3_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_asn_1_itm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_asn_1_itm_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_4;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_5;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_6;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_7;
  reg PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_3;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_4;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_5;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_6;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_7;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_3;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_4;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_5;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_6;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_7;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_8;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_9;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_3;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_4;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_1;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_2;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_3;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_4;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_5;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_6;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_7;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_8;
  reg PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_9;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_6_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_22_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_30_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_38_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_46_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_and_8_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_25_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_41_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_and_15_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_26_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_42_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_3_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_27_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_43_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_4_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_28_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_44_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_5_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_21_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_29_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_45_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_for_and_45_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_7_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_23_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_31_itm_1;
  reg [7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_47_itm_1;
  reg [5:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_1;
  reg [5:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_1;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_2;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_1;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_2;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_1;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_1;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_2;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_1;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_1;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_2;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_1;
  reg [6:0] input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_1;
  reg input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_2;
  reg [7:0] weight_mem_banks_load_store_1_for_3_result_val_Marshall_64U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1;
  reg [7:0] weight_mem_banks_load_store_1_for_5_result_val_Marshall_64U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_3;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_14_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_15_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_17_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_3;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_19_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_20_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_2_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_2_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_34_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_34_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_35_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_35_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_44_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_54_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_56_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_56_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_46_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_47_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_48_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_6_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_6_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_60_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_62_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_2;
  reg pe_manager_base_weight_slc_pe_manager_base_weight_0_12_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_71_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_72_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_76_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_78_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_80_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_10_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_84_itm_1;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_86_itm_2;
  reg crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_95_itm_2;
  reg [1:0] pe_manager_base_weight_slc_pe_manager_base_weight_1_0_1_itm_1;
  reg weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_20_itm_1;
  reg weight_mem_run_3_for_5_and_162_itm_1;
  reg weight_mem_run_3_for_5_and_162_itm_2;
  reg weight_mem_run_3_for_5_and_163_itm_1;
  reg weight_mem_run_3_for_5_and_164_itm_1;
  reg weight_mem_run_3_for_5_and_164_itm_2;
  reg weight_mem_run_3_for_5_and_165_itm_1;
  reg weight_mem_run_3_for_5_and_166_itm_1;
  reg weight_mem_run_3_for_5_and_167_itm_1;
  reg weight_mem_run_3_for_5_and_168_itm_1;
  reg weight_mem_run_3_for_5_and_8_itm_1;
  reg weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_1;
  reg weight_mem_run_3_for_5_and_20_itm_1;
  reg weight_mem_run_3_for_5_and_20_itm_2;
  reg weight_mem_run_3_for_5_and_22_itm_1;
  reg weight_mem_run_3_for_5_and_23_itm_1;
  reg weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_3_itm_1;
  reg weight_mem_run_3_for_5_and_28_itm_1;
  reg weight_mem_run_3_for_5_and_30_itm_1;
  reg weight_mem_run_3_for_5_and_30_itm_2;
  reg weight_mem_run_3_for_5_and_31_itm_1;
  reg weight_mem_run_3_for_5_and_31_itm_2;
  reg weight_mem_run_3_for_5_and_38_itm_1;
  reg weight_mem_run_3_for_5_and_39_itm_1;
  reg weight_mem_run_3_for_5_and_39_itm_2;
  reg weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_5_itm_1;
  reg weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_5_itm_2;
  reg weight_mem_run_3_for_5_and_44_itm_1;
  reg weight_mem_run_3_for_5_and_44_itm_2;
  reg weight_mem_run_3_for_5_and_46_itm_1;
  reg weight_mem_run_3_for_5_and_46_itm_2;
  reg weight_mem_run_3_for_5_and_47_itm_1;
  reg weight_mem_run_3_for_5_and_48_itm_1;
  reg weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_10_itm_1;
  reg weight_mem_run_3_for_5_and_84_itm_1;
  reg weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_12_itm_1;
  reg weight_mem_run_3_for_5_and_102_itm_1;
  reg weight_mem_run_3_for_5_and_102_itm_2;
  reg weight_mem_run_3_for_5_and_103_itm_1;
  reg weight_mem_run_3_for_5_and_103_itm_2;
  reg weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_13_itm_1;
  reg weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_13_itm_2;
  reg weight_mem_run_3_for_5_and_110_itm_1;
  reg weight_mem_run_3_for_5_and_111_itm_1;
  reg weight_mem_run_3_for_5_and_112_itm_1;
  reg weight_mem_run_3_for_5_and_156_itm_1;
  reg weight_mem_run_3_for_5_and_156_itm_2;
  reg ProductSum_for_asn_98_itm_1;
  reg ProductSum_for_asn_98_itm_2;
  reg ProductSum_for_asn_98_itm_3;
  reg ProductSum_for_asn_98_itm_4;
  reg ProductSum_for_asn_82_itm_1;
  reg ProductSum_for_asn_82_itm_2;
  reg ProductSum_for_asn_82_itm_3;
  reg ProductSum_for_asn_82_itm_4;
  reg ProductSum_for_asn_73_itm_1;
  reg ProductSum_for_asn_73_itm_2;
  reg ProductSum_for_asn_73_itm_4;
  reg ProductSum_for_asn_64_itm_2;
  reg ProductSum_for_asn_64_itm_4;
  reg ProductSum_for_asn_51_itm_2;
  reg ProductSum_for_asn_51_itm_4;
  reg ProductSum_for_asn_42_itm_2;
  reg ProductSum_for_asn_42_itm_4;
  reg ProductSum_for_asn_25_itm_2;
  reg ProductSum_for_asn_25_itm_4;
  reg ProductSum_for_asn_16_itm_2;
  reg ProductSum_for_asn_16_itm_4;
  reg accum_vector_operator_1_for_asn_1_itm_7;
  reg accum_vector_operator_1_for_asn_10_itm_7;
  reg accum_vector_operator_1_for_asn_22_itm_7;
  reg accum_vector_operator_1_for_asn_28_itm_7;
  reg accum_vector_operator_1_for_asn_37_itm_7;
  reg accum_vector_operator_1_for_asn_46_itm_7;
  reg accum_vector_operator_1_for_asn_55_itm_7;
  reg accum_vector_operator_1_for_asn_64_itm_7;
  reg [14:0] PEManager_15U_PEManagerWrite_slc_rva_in_reg_data_30_16_itm_1;
  reg while_if_mux_19_itm_1;
  reg PECore_PushAxiRsp_mux_10_itm_1;
  reg PECore_PushAxiRsp_mux_13_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_57_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_26_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_27_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_28_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_29_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_131_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_99_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_100_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_101_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_102_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_103_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_104_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_204_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_172_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_173_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_174_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_175_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_176_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_177_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_277_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_245_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_246_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_247_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_248_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_249_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_250_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_350_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_318_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_319_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_320_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_321_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_322_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_323_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_423_itm_1;
  reg Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_391_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_392_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_395_itm_1;
  reg Arbiter_8U_Roundrobin_pick_1_mux_576_itm_1;
  reg [22:0] accum_vector_data_acc_10_itm_1;
  wire [23:0] nl_accum_vector_data_acc_10_itm_1;
  reg [22:0] accum_vector_data_acc_13_itm_1;
  wire [23:0] nl_accum_vector_data_acc_13_itm_1;
  reg [22:0] accum_vector_data_acc_19_itm_1;
  wire [23:0] nl_accum_vector_data_acc_19_itm_1;
  reg [22:0] accum_vector_data_acc_22_itm_1;
  wire [23:0] nl_accum_vector_data_acc_22_itm_1;
  reg [22:0] accum_vector_data_acc_25_itm_1;
  wire [23:0] nl_accum_vector_data_acc_25_itm_1;
  reg [22:0] accum_vector_data_acc_28_itm_1;
  wire [23:0] nl_accum_vector_data_acc_28_itm_1;
  reg [22:0] accum_vector_data_acc_30_itm_1;
  wire [23:0] nl_accum_vector_data_acc_30_itm_1;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_2;
  reg weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_2;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_2;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_5;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_6;
  reg PECore_PushOutput_PECore_PushOutput_if_and_svs_st_7;
  reg [55:0] weight_mem_banks_read_1_read_data_lpi_1_dfm_1_63_8;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_2;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_0;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_3;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1_1;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_0;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_3;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_2;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_0;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_0;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_0;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_3;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_2;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_0;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_3;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_3;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_2;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_0;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_3;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_1;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_3;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_2;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_0;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_3;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_3;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_2;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_1;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_0;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_3;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_0;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_2;
  reg Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_0;
  reg [31:0] input_mem_banks_read_read_data_lpi_1_dfm_1_5_31_0;
  reg [31:0] input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0;
  reg [1:0] weight_read_addrs_2_14_1_lpi_1_dfm_2_1_0;
  reg [1:0] weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0;
  reg weight_read_addrs_4_14_2_lpi_1_dfm_3_0;
  reg [1:0] weight_read_addrs_6_14_1_lpi_1_dfm_2_1_0;
  reg [1:0] weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_6;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_5;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_4;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_3;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_2;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_1;
  reg nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_0;
  wire [7:0] weight_port_read_out_data_7_3_sva_dfm_2;
  wire [7:0] weight_port_read_out_data_7_2_sva_dfm_2;
  wire [7:0] weight_port_read_out_data_7_5_sva_dfm_2;
  wire [7:0] weight_port_read_out_data_7_4_sva_dfm_2;
  wire [7:0] weight_port_read_out_data_7_7_sva_dfm_2;
  wire [7:0] weight_port_read_out_data_7_6_sva_dfm_2;
  wire [7:0] weight_port_read_out_data_5_3_sva_dfm_2;
  wire [7:0] weight_port_read_out_data_5_2_sva_dfm_2;
  wire [7:0] weight_port_read_out_data_5_5_sva_dfm_2;
  wire [7:0] weight_port_read_out_data_5_4_sva_dfm_2;
  wire [7:0] weight_port_read_out_data_5_7_sva_dfm_2;
  wire [7:0] weight_port_read_out_data_5_6_sva_dfm_2;
  wire [7:0] weight_port_read_out_data_3_5_sva_dfm_2;
  wire [7:0] weight_port_read_out_data_3_4_sva_dfm_2;
  wire [7:0] weight_port_read_out_data_3_7_sva_dfm_2;
  wire [7:0] weight_port_read_out_data_3_6_sva_dfm_2;
  wire PECore_PushAxiRsp_if_else_mux_13_mx0w2;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_10_itm_mx0w0;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_84_itm_mx0w0;
  wire weight_mem_read_arbxbar_arbiters_next_5_2_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_5_5_sva_mx1;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_36_mx1w0;
  wire weight_mem_read_arbxbar_arbiters_next_5_7_sva_mx0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_34_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_33_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_32_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_31_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_30_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_29_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_27_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_26_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_25_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_24_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_23_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_22_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_20_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_19_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_18_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_17_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_16_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_15_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_13_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_12_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_11_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_10_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_9_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_8_mx1w0;
  wire weight_mem_read_arbxbar_arbiters_next_0_3_sva_mx1;
  wire weight_mem_read_arbxbar_arbiters_next_0_4_sva_mx1;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_2_mx1w0;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_1_mx1w0;
  wire [14:0] weight_read_addrs_1_lpi_1_dfm_1_1;
  wire [13:0] weight_read_addrs_2_14_1_lpi_1_dfm_1_1;
  wire [14:0] weight_read_addrs_3_lpi_1_dfm_1_1;
  wire [12:0] weight_read_addrs_4_14_2_lpi_1_dfm_1_1;
  wire [14:0] weight_read_addrs_5_lpi_1_dfm_1_1;
  wire [13:0] weight_read_addrs_6_14_1_lpi_1_dfm_1_1;
  wire [14:0] weight_read_addrs_7_lpi_1_dfm_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_0_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_2_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_6_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_0_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_5_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_2_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_3_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_6_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_0_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_5_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_2_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_3_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_6_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_0_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_5_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_2_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_3_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_6_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_0_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_5_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_4_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_2_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_3_1;
  wire accum_vector_data_6_sva_1_load_mx0w1;
  wire [7:0] pe_config_output_counter_sva_mx1;
  wire pe_config_is_zero_first_sva_mx1;
  wire pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1_1;
  wire [19:0] act_port_reg_data_19_0_sva_mx1;
  wire [19:0] act_port_reg_data_51_32_sva_mx1;
  wire [19:0] act_port_reg_data_83_64_sva_mx1;
  wire [19:0] act_port_reg_data_115_96_sva_mx1;
  wire [19:0] act_port_reg_data_147_128_sva_mx1;
  wire [19:0] act_port_reg_data_179_160_sva_mx1;
  wire [19:0] act_port_reg_data_211_192_sva_mx1;
  wire [19:0] act_port_reg_data_243_224_sva_mx1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_94_itm_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_71_itm_1_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_72_itm_1_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6_mx1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0_mx1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5_mx1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1_mx1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4_mx1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2_mx1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3_mx1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_9_itm_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_7_itm_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_6_itm_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_95_itm_mx0w0;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_mx0w0;
  wire [22:0] accum_vector_data_7_sva_5_mx1w0;
  wire [22:0] accum_vector_data_7_sva_4_mx0w0;
  wire [22:0] accum_vector_data_6_sva_5_mx1w0;
  wire [22:0] accum_vector_data_6_sva_4_mx0w0;
  wire [22:0] accum_vector_data_5_sva_5_mx0w0;
  wire [22:0] accum_vector_data_5_sva_4_mx1w0;
  wire [22:0] accum_vector_data_4_sva_5_mx1w0;
  wire [22:0] accum_vector_data_4_sva_4_mx1w0;
  wire [22:0] accum_vector_data_3_sva_5_mx1w0;
  wire [22:0] accum_vector_data_3_sva_4_mx1w0;
  wire [22:0] accum_vector_data_2_sva_6_mx1w0;
  wire [22:0] accum_vector_data_2_sva_5_mx1w0;
  wire [22:0] accum_vector_data_2_sva_4_mx1w0;
  wire [22:0] accum_vector_data_1_sva_5_mx1w0;
  wire [22:0] accum_vector_data_1_sva_4_mx1w0;
  wire [22:0] accum_vector_data_0_sva_5_mx1w0;
  wire [22:0] accum_vector_data_0_sva_4_mx1w0;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_1_1;
  wire [22:0] accum_vector_data_7_sva_7_mx1w0;
  wire [22:0] accum_vector_data_7_sva_6_mx1w0;
  wire [22:0] accum_vector_data_6_sva_7_mx1w0;
  wire [22:0] accum_vector_data_6_sva_6_mx1w0;
  wire [22:0] accum_vector_data_5_sva_7_mx1w0;
  wire [22:0] accum_vector_data_5_sva_6_mx1w0;
  wire [22:0] accum_vector_data_4_sva_7_mx1w0;
  wire [22:0] accum_vector_data_4_sva_6_mx1w0;
  wire [22:0] accum_vector_data_3_sva_7_mx1w0;
  wire [22:0] accum_vector_data_3_sva_6_mx1w0;
  wire [22:0] accum_vector_data_1_sva_7_mx1w0;
  wire [22:0] accum_vector_data_1_sva_6_mx1w0;
  wire [22:0] accum_vector_data_0_sva_7_mx1w0;
  wire [22:0] accum_vector_data_0_sva_6_mx1w0;
  wire PECore_PushAxiRsp_if_else_mux_10_mx0w2;
  wire [6:0] rva_out_reg_data_62_56_sva_dfm_6_mx1;
  wire [3:0] rva_out_reg_data_35_32_sva_dfm_6_mx1;
  wire PECore_PushAxiRsp_mux_13_itm_1_mx0c1;
  wire [63:0] input_mem_banks_bank_a_0_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_1_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_2_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_3_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_4_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_5_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_6_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_7_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_8_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_9_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_10_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_11_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_12_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_13_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_14_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_15_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_16_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_17_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_18_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_19_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_20_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_21_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_22_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_23_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_24_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_25_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_26_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_27_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_28_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_29_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_30_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_31_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_32_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_33_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_34_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_35_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_36_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_37_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_38_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_39_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_40_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_41_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_42_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_43_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_44_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_45_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_46_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_47_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_48_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_49_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_50_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_51_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_52_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_53_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_54_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_55_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_56_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_57_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_58_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_59_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_60_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_61_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_62_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_63_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_64_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_65_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_66_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_67_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_68_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_69_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_70_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_71_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_72_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_73_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_74_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_75_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_76_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_77_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_78_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_79_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_80_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_81_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_82_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_83_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_84_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_85_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_86_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_87_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_88_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_89_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_90_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_91_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_92_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_93_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_94_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_95_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_96_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_97_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_98_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_99_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_100_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_101_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_102_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_103_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_104_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_105_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_106_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_107_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_108_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_109_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_110_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_111_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_112_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_113_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_114_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_115_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_116_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_117_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_118_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_119_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_120_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_121_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_122_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_123_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_124_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_125_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_126_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_127_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_128_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_129_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_130_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_131_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_132_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_133_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_134_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_135_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_136_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_137_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_138_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_139_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_140_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_141_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_142_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_143_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_144_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_145_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_146_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_147_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_148_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_149_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_150_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_151_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_152_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_153_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_154_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_155_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_156_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_157_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_158_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_159_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_160_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_161_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_162_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_163_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_164_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_165_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_166_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_167_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_168_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_169_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_170_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_171_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_172_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_173_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_174_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_175_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_176_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_177_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_178_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_179_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_180_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_181_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_182_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_183_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_184_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_185_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_186_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_187_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_188_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_189_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_190_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_191_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_192_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_193_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_194_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_195_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_196_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_197_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_198_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_199_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_200_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_201_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_202_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_203_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_204_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_205_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_206_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_207_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_208_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_209_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_210_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_211_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_212_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_213_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_214_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_215_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_216_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_217_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_218_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_219_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_220_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_221_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_222_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_223_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_224_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_225_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_226_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_227_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_228_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_229_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_230_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_231_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_232_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_233_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_234_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_235_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_236_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_237_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_238_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_239_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_240_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_241_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_242_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_243_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_244_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_245_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_246_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_247_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_248_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_249_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_250_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_251_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_252_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_253_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_254_sva_dfm_2_mx1;
  wire [63:0] input_mem_banks_bank_a_255_sva_dfm_2_mx1;
  wire accum_vector_data_3_sva_1_load_mx0w0;
  wire accum_vector_data_2_sva_1_load_mx0w0;
  wire accum_vector_data_1_sva_1_load_mx0w0;
  wire accum_vector_data_0_sva_1_load_mx0w0;
  wire [14:0] pe_manager_base_input_sva_mx2;
  wire accum_vector_data_7_sva_1_load_mx0w1;
  wire accum_vector_data_5_sva_1_load_mx0w1;
  wire accum_vector_data_4_sva_1_load_mx0w1;
  wire PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  wire [7:0] BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1;
  wire weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_1_m1c_1;
  wire weight_mem_banks_load_store_1_for_else_else_and_10_m1c_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_sva_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_7_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_7_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_7_sva_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_6_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_6_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_6_sva_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_5_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_5_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_5_sva_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_4_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_4_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_4_sva_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_3_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_3_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_3_sva_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_2_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_2_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_2_sva_1;
  wire operator_2_false_3_operator_2_false_3_or_mdf_1_sva_1;
  wire operator_2_false_4_operator_2_false_4_or_mdf_1_sva_1;
  wire operator_2_false_5_operator_2_false_5_or_mdf_1_sva_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_3_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_4_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_5_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_6_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_0_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_2_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_1_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_3_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_4_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_5_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_6_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_0_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_2_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_1_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_3_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_4_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_5_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_6_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_0_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_2_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_1_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_3_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_4_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_5_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_6_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_0_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_2_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_1_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_3_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_4_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_5_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_6_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_0_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_2_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_1_mx0;
  wire weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1;
  wire [3:0] weight_read_addrs_0_3_0_lpi_1_dfm_4;
  wire while_and_1129_cse_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_pmx_sva_1;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000002;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000003;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000004;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000005;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000006;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_6_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_5_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_3_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_6_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_5_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_3_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000002;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000003;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000002;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000003;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000004;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000005;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_pmx_000000;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000006;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000000;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000001;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000002;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000003;
  wire [7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000004;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_3_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_4_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_5_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_6_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_0_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_2_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_1_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_3_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_4_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_5_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_6_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_0_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_2_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_1_mx0;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_0_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_9;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_9;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_9;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_9;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_10;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_10;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_10;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_10;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_11;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_11;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_11;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_11;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_12;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_12;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_12;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_12;
  wire rva_out_reg_data_63_sva_dfm_7;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_257_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_255_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_256_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_254_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_255_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_253_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_254_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_252_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_253_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_251_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_252_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_250_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_251_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_249_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_250_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_248_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_249_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_247_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_248_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_246_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_247_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_245_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_246_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_244_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_245_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_243_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_244_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_242_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_243_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_241_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_242_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_240_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_241_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_239_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_240_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_238_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_239_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_237_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_238_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_236_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_237_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_235_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_236_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_234_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_235_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_233_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_234_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_232_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_233_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_231_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_232_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_230_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_231_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_229_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_230_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_228_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_229_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_227_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_228_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_226_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_227_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_225_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_226_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_224_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_225_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_223_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_224_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_222_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_223_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_221_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_222_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_220_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_221_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_219_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_220_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_218_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_219_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_217_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_218_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_216_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_217_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_215_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_216_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_214_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_215_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_213_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_214_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_212_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_213_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_211_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_212_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_210_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_211_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_209_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_210_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_208_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_209_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_207_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_208_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_206_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_207_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_205_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_206_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_204_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_205_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_203_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_204_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_202_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_203_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_201_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_202_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_200_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_201_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_199_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_200_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_198_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_199_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_197_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_198_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_196_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_197_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_195_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_196_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_194_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_195_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_193_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_194_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_192_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_193_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_191_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_192_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_190_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_191_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_189_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_190_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_188_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_189_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_187_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_188_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_186_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_187_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_185_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_186_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_184_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_185_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_183_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_184_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_182_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_183_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_181_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_182_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_180_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_181_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_179_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_180_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_178_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_179_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_177_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_178_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_176_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_177_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_175_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_176_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_174_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_175_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_173_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_174_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_172_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_173_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_171_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_172_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_170_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_171_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_169_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_170_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_168_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_169_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_167_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_168_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_166_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_167_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_165_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_166_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_164_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_165_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_163_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_164_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_162_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_163_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_161_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_162_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_160_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_161_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_159_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_160_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_158_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_159_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_157_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_158_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_156_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_157_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_155_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_156_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_154_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_155_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_153_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_154_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_152_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_153_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_151_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_152_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_150_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_151_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_149_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_150_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_148_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_149_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_147_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_148_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_146_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_147_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_145_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_146_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_144_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_145_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_143_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_144_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_142_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_143_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_141_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_142_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_140_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_141_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_139_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_140_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_138_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_139_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_137_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_138_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_136_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_137_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_135_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_136_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_134_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_135_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_133_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_134_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_132_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_133_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_131_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_132_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_130_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_131_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_129_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_130_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_128_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_129_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_127_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_128_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_126_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_127_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_125_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_126_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_124_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_125_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_123_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_124_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_122_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_123_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_121_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_122_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_120_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_121_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_119_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_120_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_118_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_119_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_117_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_118_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_116_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_117_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_115_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_116_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_114_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_115_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_113_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_114_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_112_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_113_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_111_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_112_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_110_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_111_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_109_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_110_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_108_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_109_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_107_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_108_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_106_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_107_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_105_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_106_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_104_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_105_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_103_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_104_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_102_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_103_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_101_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_102_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_100_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_101_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_99_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_100_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_98_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_99_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_97_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_98_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_96_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_97_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_95_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_96_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_94_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_95_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_93_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_94_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_92_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_93_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_91_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_92_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_90_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_91_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_89_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_90_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_88_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_89_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_87_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_88_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_86_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_87_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_85_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_86_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_84_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_85_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_83_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_84_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_82_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_83_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_81_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_82_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_80_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_81_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_79_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_80_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_78_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_79_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_77_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_78_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_76_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_77_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_75_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_76_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_74_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_75_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_73_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_74_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_72_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_73_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_71_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_72_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_70_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_71_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_69_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_70_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_68_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_69_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_67_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_68_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_66_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_67_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_65_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_66_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_64_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_65_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_63_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_64_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_62_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_63_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_61_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_62_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_60_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_61_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_59_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_60_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_58_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_59_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_57_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_58_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_56_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_57_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_55_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_56_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_54_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_55_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_53_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_54_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_52_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_53_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_51_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_52_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_50_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_51_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_49_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_50_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_48_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_49_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_47_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_48_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_46_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_47_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_45_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_46_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_44_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_45_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_43_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_44_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_42_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_43_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_41_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_42_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_40_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_41_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_39_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_40_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_38_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_39_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_37_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_38_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_36_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_37_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_35_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_36_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_34_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_35_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_33_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_34_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_32_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_33_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_31_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_32_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_30_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_31_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_29_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_30_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_28_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_29_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_27_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_28_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_26_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_27_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_25_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_26_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_24_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_25_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_23_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_24_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_22_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_23_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_21_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_22_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_20_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_21_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_19_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_20_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_18_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_19_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_17_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_18_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_16_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_17_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_15_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_16_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_14_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_15_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_13_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_14_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_12_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_13_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_11_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_12_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_10_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_11_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_9_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_10_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_8_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_9_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_7_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_8_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_6_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_7_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_5_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_6_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_4_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_5_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_3_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_4_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_2_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_3_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_1_tmp_1;
  wire input_mem_write_arbxbar_xbar_1_for_3_if_1_and_2_tmp_1;
  wire input_mem_write_arbxbar_xbar_for_3_if_1_and_tmp_1;
  wire PECore_DecodeAxiRead_case_4_switch_lp_nor_5_cse_1;
  wire PECore_DecodeAxiRead_switch_lp_nor_13_cse_1;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_not_185;
  wire PECore_PushAxiRsp_if_asn_55;
  wire PECore_PushAxiRsp_if_asn_57;
  wire PECore_PushAxiRsp_if_asn_59;
  wire weight_mem_run_3_for_5_asn_309;
  wire weight_mem_run_3_for_5_asn_311;
  wire weight_mem_run_3_for_5_asn_313;
  wire weight_mem_run_3_for_5_asn_315;
  wire weight_mem_run_3_for_5_asn_317;
  wire weight_mem_run_3_for_5_asn_319;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_118;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_120;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_122;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_124;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_asn_56;
  wire weight_mem_run_3_for_5_asn_321;
  wire weight_mem_run_3_for_5_asn_323;
  wire PECore_PushAxiRsp_if_asn_61;
  wire PECore_PushAxiRsp_if_asn_63;
  wire PECore_PushAxiRsp_if_asn_65;
  wire weight_mem_run_3_for_5_and_166;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_98;
  wire weight_mem_run_3_for_5_and_168;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_100;
  wire weight_mem_run_3_for_5_and_172;
  wire weight_mem_run_3_for_5_and_174;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_and_52;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_and_54;
  wire [7:0] pe_manager_base_input_sva_mx1_7_0;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_0;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_2;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_1;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_0;
  wire mux_246_cse;
  wire PECore_PushAxiRsp_if_mux1h_15;
  wire PECore_PushAxiRsp_if_mux1h_17;
  reg reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_20_itm_2_cse;
  reg reg_weight_mem_run_3_for_5_and_163_itm_2_cse;
  reg reg_weight_mem_run_3_for_5_and_165_itm_2_cse;
  reg reg_weight_mem_run_3_for_5_and_166_itm_2_cse;
  reg reg_weight_mem_run_3_for_5_and_167_itm_2_cse;
  reg reg_weight_mem_run_3_for_5_and_168_itm_2_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_5_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_1_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_2_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_3_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_5_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_5_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_6_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_5_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_4_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_5_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_cse;
  reg reg_rva_in_reg_rw_sva_2_cse;
  reg reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_2_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_5_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_5_cse;
  reg reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4_cse;
  reg reg_PECore_RunMac_PECore_RunMac_if_and_svs_st_8_cse;
  wire weight_mem_run_3_for_5_and_161_cse;
  wire nor_320_cse;
  reg weight_mem_run_3_for_5_mux_10_itm_1_7;
  reg [6:0] weight_mem_run_3_for_5_mux_10_itm_1_6_0;
  wire weight_mem_run_3_for_5_and_209_ssc;
  reg weight_mem_run_3_for_5_mux_11_itm_1_7;
  reg [6:0] weight_mem_run_3_for_5_mux_11_itm_1_6_0;
  reg [1:0] weight_mem_run_3_for_5_mux_12_itm_1_7_6;
  reg [5:0] weight_mem_run_3_for_5_mux_12_itm_1_5_0;
  wire weight_mem_banks_load_store_for_else_and_4_ssc;
  reg [3:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1_7_4;
  reg [3:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1_3_0;
  wire weight_mem_banks_load_store_for_else_and_27_ssc;
  reg weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1_7;
  reg [6:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1_6_0;
  reg weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_itm_1_7;
  reg [6:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_itm_1_6_0;
  reg weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1_7;
  reg [6:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1_6_0;
  wire weight_mem_banks_load_store_for_else_and_20_ssc;
  reg [1:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_itm_1_7_6;
  reg [5:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_itm_1_5_0;
  reg [3:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1_7_4;
  reg [3:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1_3_0;
  wire weight_mem_banks_load_store_for_else_and_10_ssc;
  reg weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1_7;
  reg [6:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1_6_0;
  wire and_922_ssc;
  wire weight_port_read_out_data_0_0_sva_dfm_mx0w0_7;
  wire [6:0] weight_port_read_out_data_0_0_sva_dfm_mx0w0_6_0;
  wire weight_port_read_out_data_0_1_sva_dfm_mx0w0_7;
  wire [6:0] weight_port_read_out_data_0_1_sva_dfm_mx0w0_6_0;
  wire and_940_ssc;
  wire weight_port_read_out_data_0_2_sva_dfm_mx0w0_7;
  wire weight_port_read_out_data_0_2_sva_dfm_mx0w0_6;
  wire [5:0] weight_port_read_out_data_0_2_sva_dfm_mx0w0_5_0;
  wire weight_port_read_out_data_0_3_sva_dfm_mx0w0_7;
  wire [2:0] weight_port_read_out_data_0_3_sva_dfm_mx0w0_6_4;
  wire [3:0] weight_port_read_out_data_0_3_sva_dfm_mx0w0_3_0;
  wire [3:0] crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_8_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_64_63_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_2_0_8_7_0_sdt_47_40_sva_1_7_4;
  wire [3:0] crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_8_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_64_63_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_2_0_8_7_0_sdt_47_40_sva_1_3_0;
  wire weight_port_read_out_data_0_7_sva_dfm_3_7;
  wire [6:0] weight_port_read_out_data_0_7_sva_dfm_3_6_0;
  wire and_967_ssc;
  wire and_968_ssc;
  wire and_969_ssc;
  wire and_970_ssc;
  wire and_971_ssc;
  wire and_972_ssc;
  wire and_973_ssc;
  wire nor_528_ssc;
  wire [3:0] weight_port_read_out_data_0_5_sva_dfm_3_7_4;
  wire [3:0] weight_port_read_out_data_0_5_sva_dfm_3_3_0;
  wire and_976_ssc;
  wire and_979_ssc;
  wire and_980_ssc;
  wire weight_port_read_out_data_0_4_sva_dfm_3_7;
  wire weight_port_read_out_data_0_4_sva_dfm_3_6;
  wire [5:0] weight_port_read_out_data_0_4_sva_dfm_3_5_0;
  reg weight_port_read_out_data_0_1_sva_dfm_2_7;
  reg [6:0] weight_port_read_out_data_0_1_sva_dfm_2_6_0;
  reg weight_port_read_out_data_0_3_sva_dfm_1_7;
  reg [2:0] weight_port_read_out_data_0_3_sva_dfm_1_6_4;
  reg [3:0] weight_port_read_out_data_0_3_sva_dfm_1_3_0;
  wire weight_port_read_out_data_and_100_ssc;
  reg weight_port_read_out_data_0_0_sva_dfm_1_7;
  reg weight_port_read_out_data_0_1_sva_dfm_1_7;
  reg weight_port_read_out_data_0_2_sva_dfm_1_7;
  reg weight_port_read_out_data_0_2_sva_dfm_1_6;
  reg [5:0] weight_port_read_out_data_0_2_sva_dfm_1_5_0;
  reg weight_port_read_out_data_0_0_sva_dfm_2_7;
  reg [6:0] weight_port_read_out_data_0_0_sva_dfm_2_6_0;
  reg weight_port_read_out_data_0_2_sva_dfm_2_7;
  reg weight_port_read_out_data_0_2_sva_dfm_2_6;
  reg [5:0] weight_port_read_out_data_0_2_sva_dfm_2_5_0;
  reg weight_port_read_out_data_0_3_sva_dfm_2_7;
  reg [2:0] weight_port_read_out_data_0_3_sva_dfm_2_6_4;
  reg [3:0] weight_port_read_out_data_0_3_sva_dfm_2_3_0;
  reg weight_port_read_out_data_0_4_sva_dfm_2_7;
  reg weight_port_read_out_data_0_4_sva_dfm_2_6;
  reg [5:0] weight_port_read_out_data_0_4_sva_dfm_2_5_0;
  reg [3:0] weight_port_read_out_data_0_5_sva_dfm_2_7_4;
  reg [3:0] weight_port_read_out_data_0_5_sva_dfm_2_3_0;
  wire weight_port_read_out_data_and_42_ssc;
  reg [3:0] weight_port_read_out_data_0_6_sva_dfm_2_7_4;
  reg [3:0] weight_port_read_out_data_0_6_sva_dfm_2_3_0;
  reg weight_port_read_out_data_0_7_sva_dfm_2_7;
  reg [6:0] weight_port_read_out_data_0_7_sva_dfm_2_6_0;
  reg [3:0] rva_out_reg_data_55_48_sva_dfm_4_1_7_4;
  reg [3:0] rva_out_reg_data_55_48_sva_dfm_4_1_3_0;
  reg [2:0] rva_out_reg_data_46_40_sva_dfm_4_1_6_4;
  reg [3:0] rva_out_reg_data_46_40_sva_dfm_4_1_3_0;
  reg rva_out_reg_data_39_36_sva_dfm_4_1_3;
  reg rva_out_reg_data_39_36_sva_dfm_4_1_2;
  reg [1:0] rva_out_reg_data_39_36_sva_dfm_4_1_1_0;
  wire weight_mem_run_3_for_5_and_179_ssc;
  wire PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_a_mx1_7;
  wire [6:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_a_mx1_6_0;
  wire weight_port_read_out_data_0_0_sva_dfm_3_7;
  wire [6:0] weight_port_read_out_data_0_0_sva_dfm_3_6_0;
  reg [3:0] weight_mem_run_3_for_5_mux_6_itm_1_7_4;
  reg [3:0] weight_mem_run_3_for_5_mux_6_itm_1_3_0;
  reg [3:0] rva_out_reg_data_55_48_sva_dfm_4_2_7_4;
  reg [3:0] rva_out_reg_data_55_48_sva_dfm_4_2_3_0;
  reg [2:0] rva_out_reg_data_46_40_sva_dfm_4_2_6_4;
  reg [3:0] rva_out_reg_data_46_40_sva_dfm_4_2_3_0;
  reg rva_out_reg_data_39_36_sva_dfm_4_2_3;
  reg rva_out_reg_data_39_36_sva_dfm_4_2_2;
  reg [1:0] rva_out_reg_data_39_36_sva_dfm_4_2_1_0;
  reg weight_port_read_out_data_0_3_sva_dfm_2_7_1;
  reg [2:0] weight_port_read_out_data_0_3_sva_dfm_2_6_4_1;
  reg [3:0] weight_port_read_out_data_0_3_sva_dfm_2_3_0_1;
  reg weight_port_read_out_data_0_2_sva_dfm_2_7_1;
  reg weight_port_read_out_data_0_2_sva_dfm_2_6_1;
  reg [5:0] weight_port_read_out_data_0_2_sva_dfm_2_5_0_1;
  reg weight_port_read_out_data_0_1_sva_dfm_2_7_1;
  wire weight_port_read_out_data_and_96_ssc;
  reg weight_port_read_out_data_0_0_sva_dfm_2_7_1;
  wire weight_mem_run_3_for_5_and_182_ssc;
  wire weight_mem_run_3_for_5_and_187_ssc;
  wire weight_port_read_out_data_0_7_sva_dfm_1_1_mx0_7;
  wire [6:0] weight_port_read_out_data_0_7_sva_dfm_1_1_mx0_6_0;
  wire [3:0] rva_out_reg_data_55_48_sva_dfm_6_mx1_7_4;
  wire [3:0] rva_out_reg_data_55_48_sva_dfm_6_mx1_3_0;
  wire [2:0] rva_out_reg_data_46_40_sva_dfm_6_mx1_6_4;
  wire [3:0] rva_out_reg_data_46_40_sva_dfm_6_mx1_3_0;
  wire rva_out_reg_data_39_36_sva_dfm_6_mx1_3;
  wire rva_out_reg_data_39_36_sva_dfm_6_mx1_2;
  wire [1:0] rva_out_reg_data_39_36_sva_dfm_6_mx1_1_0;
  reg weight_port_read_out_data_0_0_sva_dfm_1_6;
  reg [5:0] weight_port_read_out_data_0_0_sva_dfm_1_5_0;
  reg [2:0] weight_port_read_out_data_0_1_sva_dfm_1_6_4;
  reg [3:0] weight_port_read_out_data_0_1_sva_dfm_1_3_0;
  wire rva_out_reg_data_and_14_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_2_cse;
  wire rva_out_reg_data_and_17_cse;
  wire input_mem_banks_read_read_data_and_cse;
  wire weight_port_read_out_data_and_68_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_cse;
  wire rva_in_reg_rw_and_cse;
  wire ProductSum_for_and_cse;
  wire weight_mem_run_3_for_aelse_and_cse;
  wire weight_mem_banks_read_1_read_data_and_8_cse;
  wire ProductSum_for_and_8_cse;
  wire weight_mem_run_3_for_aelse_and_1_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_101_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_105_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_108_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_cse;
  wire weight_mem_read_arbxbar_xbar_1_for_3_and_8_cse;
  wire weight_mem_read_arbxbar_xbar_1_for_3_and_10_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_50_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_56_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_62_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_67_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_73_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_79_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_85_cse;
  wire weight_mem_read_arbxbar_arbiters_next_and_91_cse;
  wire weight_read_addrs_and_9_cse;
  wire weight_write_data_data_and_cse;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_cse;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_14_cse;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_18_cse;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_22_cse;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_26_cse;
  wire PECore_RunFSM_switch_lp_and_cse;
  wire Arbiter_8U_Roundrobin_pick_1_and_15_cse;
  wire Arbiter_8U_Roundrobin_pick_1_and_22_cse;
  wire Arbiter_8U_Roundrobin_pick_and_cse;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_13_cse;
  wire Arbiter_8U_Roundrobin_pick_1_and_64_cse;
  wire weight_write_data_data_and_8_cse;
  wire PECore_DecodeAxiWrite_switch_lp_and_2_cse;
  wire rva_in_reg_rw_and_6_cse;
  wire PECore_UpdateFSM_switch_lp_and_9_cse;
  wire state_and_cse;
  wire PECore_PushOutput_if_and_cse;
  wire weight_port_read_out_data_and_92_cse;
  wire accum_vector_data_and_40_cse;
  wire weight_read_addrs_and_19_cse;
  wire while_if_and_10_cse;
  wire nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_30_cse;
  wire PECore_RunMac_if_and_cse;
  wire rva_in_reg_rw_and_2_cse;
  wire ProductSum_for_and_16_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_122_cse;
  wire input_mem_banks_read_read_data_and_9_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_4_cse;
  wire while_if_and_14_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_7_cse;
  wire while_if_and_6_cse;
  wire rva_out_reg_data_and_24_cse;
  wire input_read_req_valid_and_1_cse;
  wire PECore_RunScale_if_and_cse;
  wire weight_mem_banks_load_store_for_else_and_3_cse;
  wire weight_mem_banks_load_store_for_else_and_cse;
  wire weight_mem_banks_load_store_for_else_and_1_cse;
  wire weight_mem_banks_load_store_for_else_and_9_cse;
  wire weight_mem_banks_load_store_for_else_and_2_cse;
  wire weight_mem_banks_load_store_for_else_and_17_cse;
  wire weight_mem_banks_load_store_for_else_and_22_cse;
  wire rva_in_reg_rw_and_7_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_cse;
  wire PECore_RunMac_if_and_1_cse;
  wire rva_in_reg_rw_and_3_cse;
  wire ProductSum_for_and_24_cse;
  wire ProductSum_for_and_30_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_73_cse;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_72_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_8_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_11_cse;
  wire while_if_and_7_cse;
  wire rva_out_reg_data_and_32_cse;
  wire input_read_req_valid_and_2_cse;
  wire PECore_RunScale_if_and_3_cse;
  wire weight_mem_read_arbxbar_xbar_requests_transpose_and_14_cse;
  wire PECore_RunMac_if_and_2_cse;
  wire rva_in_reg_rw_and_8_cse;
  wire ProductSum_for_and_32_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_12_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_15_cse;
  wire rva_out_reg_data_and_40_cse;
  wire input_read_req_valid_and_3_cse;
  wire rva_out_reg_data_and_45_cse;
  wire rva_in_reg_rw_and_4_cse;
  wire PECore_RunScale_if_and_5_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_16_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_19_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_19_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_23_cse;
  wire rva_out_reg_data_and_51_cse;
  wire rva_out_reg_data_and_54_cse;
  wire PECore_RunMac_if_and_5_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_24_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_25_cse;
  wire rva_out_reg_data_and_59_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_27_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_29_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_30_cse;
  wire PECore_DecodeAxiRead_switch_lp_and_31_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_33_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_34_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_37_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_39_cse;
  wire PECore_DecodeAxiRead_case_4_switch_lp_and_41_cse;
  reg weight_port_read_out_data_0_7_sva_dfm_1_1_rsp_0;
  reg [6:0] weight_port_read_out_data_0_7_sva_dfm_1_1_rsp_1;
  reg weight_port_read_out_data_0_0_sva_dfm_3_rsp_0;
  reg weight_port_read_out_data_0_1_sva_dfm_3_rsp_0;
  reg weight_port_read_out_data_0_2_sva_dfm_3_rsp_0;
  reg weight_port_read_out_data_0_2_sva_dfm_3_rsp_1;
  reg [5:0] weight_port_read_out_data_0_2_sva_dfm_3_rsp_2;
  reg weight_port_read_out_data_0_3_sva_dfm_3_rsp_0;
  reg [2:0] weight_port_read_out_data_0_3_sva_dfm_3_rsp_1;
  reg [3:0] weight_port_read_out_data_0_3_sva_dfm_3_rsp_2;
  reg rva_out_reg_data_39_36_sva_dfm_4_3_rsp_0;
  reg rva_out_reg_data_39_36_sva_dfm_4_3_rsp_1;
  reg [1:0] rva_out_reg_data_39_36_sva_dfm_4_3_rsp_2;
  reg [2:0] rva_out_reg_data_46_40_sva_dfm_4_3_rsp_0;
  reg [3:0] rva_out_reg_data_46_40_sva_dfm_4_3_rsp_1;
  reg [3:0] rva_out_reg_data_55_48_sva_dfm_4_3_rsp_0;
  reg [3:0] rva_out_reg_data_55_48_sva_dfm_4_3_rsp_1;
  reg [3:0] rva_out_reg_data_55_48_sva_dfm_6_rsp_0;
  reg [3:0] rva_out_reg_data_55_48_sva_dfm_6_rsp_1;
  reg [2:0] rva_out_reg_data_46_40_sva_dfm_6_rsp_0;
  reg [3:0] rva_out_reg_data_46_40_sva_dfm_6_rsp_1;
  reg rva_out_reg_data_39_36_sva_dfm_6_rsp_0;
  reg rva_out_reg_data_39_36_sva_dfm_6_rsp_1;
  reg [1:0] rva_out_reg_data_39_36_sva_dfm_6_rsp_2;
  reg [3:0] reg_rva_out_reg_data_55_48_sva_dfm_4_4_ftd;
  reg [3:0] reg_rva_out_reg_data_55_48_sva_dfm_4_4_ftd_1;
  reg [2:0] reg_rva_out_reg_data_46_40_sva_dfm_4_4_ftd;
  reg [3:0] reg_rva_out_reg_data_46_40_sva_dfm_4_4_ftd_1;
  reg reg_rva_out_reg_data_39_36_sva_dfm_4_4_ftd;
  reg reg_rva_out_reg_data_39_36_sva_dfm_4_4_ftd_1;
  reg [1:0] reg_rva_out_reg_data_39_36_sva_dfm_4_4_ftd_2;
  reg reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_1_ftd;
  reg reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_1_ftd;
  reg reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_ftd;
  reg reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_ftd_1;
  reg [4:0] reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_ftd_2;
  reg reg_weight_port_read_out_data_0_3_sva_dfm_4_ftd;
  reg [2:0] reg_weight_port_read_out_data_0_3_sva_dfm_4_ftd_1;
  reg [3:0] reg_weight_port_read_out_data_0_3_sva_dfm_4_ftd_2;
  reg reg_weight_port_read_out_data_0_0_sva_dfm_2_1_ftd;
  reg [5:0] reg_weight_port_read_out_data_0_0_sva_dfm_2_1_ftd_1;
  reg [2:0] reg_weight_port_read_out_data_0_1_sva_dfm_2_1_ftd;
  reg [3:0] reg_weight_port_read_out_data_0_1_sva_dfm_2_1_ftd_1;
  wire PECore_PushAxiRsp_if_mux1h_10_6;
  wire PECore_PushAxiRsp_if_mux1h_12_6;
  wire PECore_PushAxiRsp_if_mux1h_14_6;
  wire PECore_PushAxiRsp_if_mux1h_14_5;
  wire [4:0] PECore_PushAxiRsp_if_mux1h_14_4_0;
  wire [2:0] PECore_PushAxiRsp_if_mux1h_16_5_3;
  wire [2:0] PECore_PushAxiRsp_if_mux1h_16_2_0;
  reg weight_port_read_out_data_0_0_sva_dfm_3_rsp_1_6;
  reg [5:0] weight_port_read_out_data_0_0_sva_dfm_3_rsp_1_5_0;
  reg [2:0] weight_port_read_out_data_0_1_sva_dfm_3_rsp_1_6_4;
  reg [3:0] weight_port_read_out_data_0_1_sva_dfm_3_rsp_1_3_0;
  reg rva_out_reg_data_7_1_sva_dfm_6_rsp_0;
  reg reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_1_ftd_1_rsp_0;
  reg [4:0] reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_1_ftd_1_rsp_1;
  reg rva_out_reg_data_15_9_sva_dfm_6_rsp_0;
  reg [2:0] reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_1_ftd_1_rsp_0;
  reg [2:0] reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_1_ftd_1_rsp_1;
  reg rva_out_reg_data_23_17_sva_dfm_6_rsp_0;
  reg rva_out_reg_data_23_17_sva_dfm_6_rsp_1;
  reg [4:0] rva_out_reg_data_23_17_sva_dfm_6_rsp_2;
  reg [2:0] rva_out_reg_data_30_25_sva_dfm_6_rsp_0;
  reg [2:0] rva_out_reg_data_30_25_sva_dfm_6_rsp_1;
  wire PECore_PushAxiRsp_if_mux1h_10_5;
  wire [4:0] PECore_PushAxiRsp_if_mux1h_10_4_0;
  wire [2:0] PECore_PushAxiRsp_if_mux1h_12_5_3;
  wire [2:0] PECore_PushAxiRsp_if_mux1h_12_2_0;
  reg rva_out_reg_data_7_1_sva_dfm_6_rsp_1_rsp_0;
  reg [4:0] rva_out_reg_data_7_1_sva_dfm_6_rsp_1_rsp_1;
  reg [2:0] rva_out_reg_data_15_9_sva_dfm_6_rsp_1_rsp_0;
  reg [2:0] rva_out_reg_data_15_9_sva_dfm_6_rsp_1_rsp_1;
  wire or_dcpl_717;
  wire or_dcpl_718;
  wire or_dcpl_727;
  wire or_tmp_720;
  wire mux_tmp_481;
  wire mux_tmp_482;
  wire mux_tmp_483;
  wire and_dcpl_759;
  wire or_dcpl_751;
  wire or_dcpl_779;
  wire or_dcpl_801;
  wire or_dcpl_824;
  wire and_dcpl_885;
  wire or_tmp_745;
  wire or_dcpl_826;
  wire or_tmp_762;
  wire or_dcpl_828;
  wire or_tmp_779;
  wire or_tmp_796;
  wire or_tmp_830;
  wire or_tmp_864;
  wire or_tmp_915;
  wire or_tmp_949;
  wire and_dcpl_964;
  wire [7:0] PEManager_15U_GetInputAddr_acc_tmp;
  wire [8:0] nl_PEManager_15U_GetInputAddr_acc_tmp;
  wire mux_tmp_1225;
  wire or_tmp_2755;
  wire or_tmp_2762;
  wire or_tmp_2778;
  wire not_tmp_1925;
  wire and_1002_cse;
  wire mux_501_cse;
  wire and_1048_cse;
  wire or_1491_cse;
  wire nor_912_cse;
  wire and_1098_cse;
  wire and_1129_cse;
  wire xor_7_cse;
  wire and_1177_cse;
  wire xor_13_cse;
  wire nor_910_cse;
  wire nor_929_cse;
  wire and_1402_cse;
  wire and_1411_cse;
  wire or_2088_cse;
  wire nand_407_cse;
  wire nand_408_cse;
  wire nand_410_cse;
  wire nand_414_cse;
  wire nand_422_cse;
  wire nor_922_cse;
  wire nor_907_cse;
  wire nor_909_cse;
  wire nand_372_cse;
  wire and_1065_cse;
  wire and_2257_cse;
  wire nor_894_cse;
  wire nor_896_cse;
  wire nor_536_cse;
  wire or_3652_cse;
  wire or_3651_cse;
  wire or_3659_cse;
  wire or_3658_cse;
  wire and_1040_cse;
  wire and_1044_cse;
  wire and_1162_cse;
  wire and_1166_cse;
  wire and_1250_cse;
  wire and_1262_cse;
  wire and_1274_cse;
  wire and_1292_cse;
  wire and_1304_cse;
  wire mux_537_cse;
  wire mux_545_cse;
  wire mux_553_cse;
  wire mux_561_cse;
  wire mux_577_cse;
  wire mux_617_cse;
  wire mux_633_cse;
  wire mux_743_cse;
  wire mux_773_cse;
  wire mux_799_cse;
  wire or_3653_cse;
  wire or_3650_cse;
  wire or_3657_cse;
  wire and_1138_cse;
  wire and_1320_cse;
  wire and_1332_cse;
  wire and_1344_cse;
  wire and_1356_cse;
  wire and_1368_cse;
  wire and_1380_cse;
  wire and_1392_cse;
  wire and_2218_cse;
  wire mux_1268_cse;
  reg reg_rva_out_reg_data_15_9_sva_dfm_8_enexo;
  reg reg_rva_out_reg_data_23_17_sva_dfm_6_enexo;
  reg reg_rva_out_reg_data_30_25_sva_dfm_6_enexo;
  reg reg_rva_out_reg_data_62_56_sva_dfm_4_3_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_4_3_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_4_3_1_enexo;
  reg reg_rva_out_reg_data_46_40_sva_dfm_4_3_1_enexo;
  reg reg_rva_out_reg_data_35_32_sva_dfm_4_3_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_1_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_1_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_1_enexo;
  reg reg_weight_port_read_out_data_0_2_sva_dfm_3_2_enexo;
  reg reg_weight_port_read_out_data_0_3_sva_dfm_3_2_enexo;
  reg reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_1_enexo;
  reg reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_4_enexo;
  reg reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_4_enexo_1;
  reg reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_000000;
  reg reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_3_enexo;
  reg reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo;
  reg reg_Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1_enexo;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0_enexo;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_3_enexo;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1_enexo;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0_enexo;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_3_enexo;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_3_enexo;
  reg reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_1;
  reg reg_Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1_enexo_1;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_0_enexo;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0_enexo_1;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_3_enexo_1;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1_enexo_1;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0_enexo_1;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_3_enexo_1;
  reg reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_3_enexo_1;
  reg reg_weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs_enexo;
  reg reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_2;
  reg reg_weight_write_data_data_0_7_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_6_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_5_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_4_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_3_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_2_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_1_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_data_data_0_0_lpi_1_dfm_1_2_6_enexo;
  reg reg_weight_write_addrs_lpi_1_dfm_1_2_enexo;
  reg reg_weight_write_data_data_0_7_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_6_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_5_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_4_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_3_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_2_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_1_lpi_1_dfm_1_1_enexo;
  reg reg_weight_write_data_data_0_0_lpi_1_dfm_1_1_enexo;
  reg reg_pe_manager_base_input_enexo;
  reg reg_weight_read_addrs_0_3_0_lpi_1_dfm_1_1_enexo;
  reg reg_pe_config_num_output_enexo;
  reg reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_1_enexo;
  reg reg_rva_in_reg_data_sva_1_enexo;
  reg reg_input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0_enexo;
  reg reg_input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0_enexo_1;
  reg reg_input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0_enexo_2;
  reg reg_input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0_enexo_3;
  reg reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_30_25_sva_dfm_5_enexo;
  reg reg_rva_out_reg_data_23_17_sva_dfm_5_enexo;
  reg reg_rva_out_reg_data_15_9_sva_dfm_7_enexo;
  reg reg_rva_out_reg_data_35_32_sva_dfm_4_2_enexo;
  reg reg_rva_out_reg_data_62_56_sva_dfm_4_2_enexo;
  reg reg_input_mem_banks_read_read_data_lpi_1_dfm_1_5_31_0_enexo;
  reg reg_weight_mem_write_arbxbar_xbar_for_empty_sva_1_enexo;
  reg reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_1_enexo;
  reg reg_weight_mem_run_3_for_5_mux_12_itm_1_1_enexo;
  reg reg_weight_mem_run_3_for_5_mux_11_itm_1_1_enexo;
  reg reg_weight_mem_run_3_for_5_mux_10_itm_1_1_enexo;
  reg reg_rva_out_reg_data_35_32_sva_dfm_4_1_enexo;
  reg reg_rva_out_reg_data_62_56_sva_dfm_4_1_enexo;
  reg reg_input_mem_banks_bank_a_167_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_86_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_242_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_165_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_186_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_110_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_187_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_246_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_129_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_175_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_239_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_227_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_138_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_174_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_11_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_79_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_71_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_82_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_97_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_188_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_162_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_205_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_93_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_54_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_38_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_192_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_209_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_220_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_139_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_196_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_207_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_224_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_204_sva_dfm_2_enexo;
  reg reg_input_write_req_valid_lpi_1_dfm_1_1_enexo;
  reg reg_input_mem_banks_bank_a_51_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_72_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_111_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_2_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_99_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_65_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_101_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_52_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_182_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_109_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_60_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_83_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_214_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_33_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_23_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_173_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_141_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_114_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_236_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_238_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_151_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_243_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_245_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_131_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_94_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_226_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_168_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_26_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_124_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_45_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_89_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_75_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_163_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_61_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_13_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_62_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_32_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_6_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_210_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_31_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_118_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_230_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_250_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_217_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_253_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_212_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_132_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_43_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_160_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_42_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_85_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_4_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_16_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_25_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_46_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_50_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_40_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_117_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_134_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_155_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_254_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_17_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_208_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_185_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_219_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_125_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_68_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_24_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_12_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_59_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_199_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_156_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_77_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_216_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_34_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_251_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_228_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_78_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_67_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_19_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_27_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_81_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_164_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_183_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_179_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_189_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_213_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_234_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_248_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_249_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_112_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_232_sva_dfm_2_enexo;
  reg reg_input_read_addrs_sva_1_1_enexo;
  reg reg_input_mem_banks_bank_a_181_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_18_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_218_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_80_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_121_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_15_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_92_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_152_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_203_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_0_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_44_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_237_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_105_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_84_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_193_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_225_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_21_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_143_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_57_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_154_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_63_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_106_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_87_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_177_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_201_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_122_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_113_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_88_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_74_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_90_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_41_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_7_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_235_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_126_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_146_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_229_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_223_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_161_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_206_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_130_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_195_sva_dfm_2_enexo;
  reg reg_input_mem_banks_read_read_data_sva_1_enexo;
  reg reg_input_mem_banks_bank_a_103_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_100_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_157_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_127_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_49_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_47_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_240_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_222_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_120_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_66_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_35_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_133_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_172_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_69_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_108_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_14_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_159_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_76_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_241_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_171_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_200_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_98_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_233_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_148_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_104_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_55_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_123_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_119_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_135_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_116_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_128_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_194_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_30_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_136_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_255_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_221_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_244_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_28_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_231_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_180_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_145_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_150_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_96_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_140_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_8_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_91_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_202_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_20_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_169_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_176_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_158_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_149_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_147_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_53_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_29_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_153_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_252_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_3_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_102_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_107_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_9_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_137_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_115_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_170_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_211_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_10_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_197_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_64_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_166_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_191_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_198_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_190_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_5_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_184_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_215_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_37_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_247_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_36_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_142_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_178_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_73_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_144_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_22_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_48_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_56_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_39_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_58_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_1_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_95_sva_dfm_2_enexo;
  reg reg_input_mem_banks_bank_a_70_sva_dfm_2_enexo;
  reg reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo;
  reg reg_rva_out_reg_data_30_25_sva_dfm_1_enexo;
  reg reg_rva_out_reg_data_23_17_sva_dfm_1_enexo;
  reg reg_rva_out_reg_data_15_9_sva_dfm_3_enexo;
  reg reg_rva_out_reg_data_35_32_sva_dfm_1_3_enexo;
  reg reg_rva_out_reg_data_39_36_sva_dfm_1_3_enexo;
  reg reg_rva_out_reg_data_46_40_sva_dfm_1_3_enexo;
  reg reg_rva_out_reg_data_62_56_sva_dfm_1_3_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_1_3_enexo;
  reg reg_rva_out_reg_data_15_9_sva_dfm_2_enexo;
  reg reg_rva_out_reg_data_35_32_sva_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_39_36_sva_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_46_40_sva_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_62_56_sva_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_15_9_sva_dfm_1_enexo;
  reg reg_rva_out_reg_data_35_32_sva_dfm_1_1_enexo;
  reg reg_rva_out_reg_data_39_36_sva_dfm_1_1_enexo;
  reg reg_rva_out_reg_data_46_40_sva_dfm_1_1_enexo;
  reg reg_rva_out_reg_data_62_56_sva_dfm_1_1_enexo;
  reg reg_pe_config_input_counter_sva_dfm_1_enexo;
  reg reg_weight_port_read_out_data_0_2_sva_dfm_2_2_enexo;
  reg reg_weight_port_read_out_data_0_3_sva_dfm_2_2_enexo;
  reg reg_rva_out_reg_data_46_40_sva_dfm_4_2_1_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_4_2_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_4_2_1_enexo;
  reg reg_weight_port_read_out_data_0_0_sva_dfm_1_2_enexo;
  reg reg_weight_port_read_out_data_0_1_sva_dfm_1_2_enexo;
  reg reg_weight_port_read_out_data_0_2_sva_dfm_1_2_enexo;
  reg reg_weight_port_read_out_data_0_3_sva_dfm_1_2_enexo;
  reg reg_rva_out_reg_data_46_40_sva_dfm_4_1_1_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_4_1_enexo;
  reg reg_rva_out_reg_data_55_48_sva_dfm_4_1_1_enexo;
  reg reg_weight_port_read_out_data_0_0_sva_dfm_3_2_enexo;
  reg reg_weight_port_read_out_data_0_0_sva_dfm_2_2_enexo;
  reg reg_weight_port_read_out_data_0_1_sva_dfm_2_2_enexo;
  wire rva_out_reg_data_and_78_enex5;
  wire rva_out_reg_data_and_79_enex5;
  wire rva_out_reg_data_and_80_enex5;
  wire rva_out_reg_data_and_81_enex5;
  wire rva_out_reg_data_and_82_enex5;
  wire rva_out_reg_data_and_83_enex5;
  wire rva_out_reg_data_and_84_enex5;
  wire rva_out_reg_data_and_85_enex5;
  wire input_mem_banks_read_read_data_and_22_enex5;
  wire input_mem_banks_read_read_data_and_23_enex5;
  wire input_mem_banks_read_read_data_and_24_enex5;
  wire weight_port_read_out_data_and_104_enex5;
  wire weight_port_read_out_data_and_105_enex5;
  wire input_mem_banks_read_read_data_and_25_enex5;
  wire input_mem_banks_read_1_read_data_and_enex5;
  wire input_mem_banks_read_1_read_data_and_6_enex5;
  wire weight_port_read_out_data_and_enex5;
  wire input_mem_banks_read_1_read_data_and_7_enex5;
  wire weight_read_addrs_and_7_enex5;
  wire weight_mem_read_arbxbar_xbar_1_for_3_and_enex5;
  wire weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5;
  wire weight_write_data_data_and_24_enex5;
  wire weight_write_data_data_and_25_enex5;
  wire weight_write_data_data_and_26_enex5;
  wire weight_write_data_data_and_27_enex5;
  wire weight_write_data_data_and_28_enex5;
  wire weight_write_data_data_and_29_enex5;
  wire weight_write_data_data_and_30_enex5;
  wire weight_write_data_data_and_31_enex5;
  wire weight_write_addrs_and_enex5;
  wire weight_write_data_data_and_32_enex5;
  wire weight_write_data_data_and_33_enex5;
  wire weight_write_data_data_and_34_enex5;
  wire weight_write_data_data_and_35_enex5;
  wire weight_write_data_data_and_36_enex5;
  wire weight_write_data_data_and_37_enex5;
  wire weight_write_data_data_and_38_enex5;
  wire weight_write_data_data_and_39_enex5;
  wire weight_write_addrs_and_2_enex5;
  wire weight_read_addrs_and_28_enex5;
  wire pe_config_UpdateManagerCounter_if_if_and_enex5;
  wire weight_read_addrs_and_29_enex5;
  wire PEManager_15U_PEManagerWrite_and_enex5;
  wire input_mem_banks_read_read_data_and_26_enex5;
  wire input_mem_banks_read_read_data_and_27_enex5;
  wire input_mem_banks_read_read_data_and_28_enex5;
  wire input_mem_banks_read_read_data_and_29_enex5;
  wire input_mem_banks_read_1_read_data_and_3_enex5;
  wire rva_out_reg_data_and_86_enex5;
  wire rva_out_reg_data_and_87_enex5;
  wire rva_out_reg_data_and_88_enex5;
  wire rva_out_reg_data_and_89_enex5;
  wire rva_out_reg_data_and_90_enex5;
  wire input_mem_banks_read_read_data_and_18_enex5;
  wire weight_mem_write_arbxbar_xbar_for_empty_and_enex5;
  wire input_mem_banks_read_1_read_data_and_4_enex5;
  wire rva_out_reg_data_and_91_enex5;
  wire rva_out_reg_data_and_92_enex5;
  wire rva_out_reg_data_and_93_enex5;
  wire rva_out_reg_data_and_94_enex5;
  wire rva_out_reg_data_and_95_enex5;
  wire input_mem_banks_read_1_read_data_and_5_enex5;
  wire input_mem_banks_read_read_data_and_19_enex5;
  wire rva_out_reg_data_and_96_enex5;
  wire rva_out_reg_data_and_97_enex5;
  wire rva_out_reg_data_and_98_enex5;
  wire rva_out_reg_data_and_99_enex5;
  wire rva_out_reg_data_and_100_enex5;
  wire rva_out_reg_data_and_101_enex5;
  wire rva_out_reg_data_and_102_enex5;
  wire rva_out_reg_data_and_103_enex5;
  wire rva_out_reg_data_and_104_enex5;
  wire rva_out_reg_data_and_105_enex5;
  wire rva_out_reg_data_and_106_enex5;
  wire rva_out_reg_data_and_107_enex5;
  wire rva_out_reg_data_and_108_enex5;
  wire rva_out_reg_data_and_109_enex5;
  wire rva_out_reg_data_and_67_enex5;
  wire rva_out_reg_data_and_110_enex5;
  wire rva_out_reg_data_and_111_enex5;
  wire rva_out_reg_data_and_112_enex5;
  wire rva_out_reg_data_and_113_enex5;
  wire rva_out_reg_data_and_114_enex5;
  wire weight_port_read_out_data_and_106_enex5;
  wire weight_port_read_out_data_and_107_enex5;
  wire rva_out_reg_data_and_115_enex5;
  wire rva_out_reg_data_and_116_enex5;
  wire rva_out_reg_data_and_117_enex5;
  wire weight_port_read_out_data_and_108_enex5;
  wire weight_port_read_out_data_and_109_enex5;
  wire weight_port_read_out_data_and_110_enex5;
  wire weight_port_read_out_data_and_111_enex5;
  wire rva_out_reg_data_and_118_enex5;
  wire rva_out_reg_data_and_119_enex5;
  wire rva_out_reg_data_and_120_enex5;
  wire weight_port_read_out_data_and_112_enex5;
  wire weight_port_read_out_data_and_113_enex5;
  wire weight_port_read_out_data_and_114_enex5;
  wire data_in_tmp_operator_2_for_and_tmp;
  wire pe_manager_base_input_and_tmp;
  wire rva_in_reg_data_and_tmp;
  wire and_1920_tmp;
  wire and_1677_tmp;
  wire and_2145_tmp;
  wire and_1914_tmp;
  wire and_1977_tmp;
  wire and_1749_tmp;
  wire and_1980_tmp;
  wire and_2157_tmp;
  wire and_1806_tmp;
  wire and_1944_tmp;
  wire and_2136_tmp;
  wire and_2100_tmp;
  wire and_1833_tmp;
  wire and_1941_tmp;
  wire and_1452_tmp;
  wire and_1656_tmp;
  wire and_1632_tmp;
  wire and_1665_tmp;
  wire and_1710_tmp;
  wire and_1983_tmp;
  wire and_1905_tmp;
  wire and_2034_tmp;
  wire and_1698_tmp;
  wire and_1581_tmp;
  wire and_1533_tmp;
  wire and_1995_tmp;
  wire and_2046_tmp;
  wire and_2079_tmp;
  wire and_1836_tmp;
  wire and_2007_tmp;
  wire and_2040_tmp;
  wire and_2091_tmp;
  wire and_2031_tmp;
  wire and_1572_tmp;
  wire and_1635_tmp;
  wire and_1752_tmp;
  wire and_1425_tmp;
  wire and_1716_tmp;
  wire and_1614_tmp;
  wire and_1722_tmp;
  wire and_1575_tmp;
  wire and_1965_tmp;
  wire and_1746_tmp;
  wire and_1599_tmp;
  wire and_1668_tmp;
  wire and_2061_tmp;
  wire and_1518_tmp;
  wire and_1488_tmp;
  wire and_1938_tmp;
  wire and_1842_tmp;
  wire and_1761_tmp;
  wire and_2127_tmp;
  wire and_2133_tmp;
  wire and_1872_tmp;
  wire and_2148_tmp;
  wire and_2154_tmp;
  wire and_1812_tmp;
  wire and_1701_tmp;
  wire and_2097_tmp;
  wire and_1923_tmp;
  wire and_1497_tmp;
  wire and_1791_tmp;
  wire and_1554_tmp;
  wire and_1686_tmp;
  wire and_1644_tmp;
  wire and_1908_tmp;
  wire and_1602_tmp;
  wire and_1458_tmp;
  wire and_1605_tmp;
  wire and_1515_tmp;
  wire and_1437_tmp;
  wire and_2049_tmp;
  wire and_1512_tmp;
  wire and_1773_tmp;
  wire and_2109_tmp;
  wire and_2169_tmp;
  wire and_2070_tmp;
  wire and_2178_tmp;
  wire and_2055_tmp;
  wire and_1815_tmp;
  wire and_1548_tmp;
  wire and_1899_tmp;
  wire and_1545_tmp;
  wire and_1674_tmp;
  wire and_1431_tmp;
  wire and_1467_tmp;
  wire and_1494_tmp;
  wire and_1557_tmp;
  wire and_1569_tmp;
  wire and_1539_tmp;
  wire and_1770_tmp;
  wire and_1821_tmp;
  wire and_1884_tmp;
  wire and_2181_tmp;
  wire and_1470_tmp;
  wire and_2043_tmp;
  wire and_1974_tmp;
  wire and_2076_tmp;
  wire and_1794_tmp;
  wire and_1623_tmp;
  wire and_1491_tmp;
  wire and_1455_tmp;
  wire and_1596_tmp;
  wire and_2016_tmp;
  wire and_1887_tmp;
  wire and_1650_tmp;
  wire and_2067_tmp;
  wire and_1521_tmp;
  wire and_2172_tmp;
  wire and_2103_tmp;
  wire and_1653_tmp;
  wire and_1620_tmp;
  wire and_1476_tmp;
  wire and_1500_tmp;
  wire and_1662_tmp;
  wire and_1911_tmp;
  wire and_1968_tmp;
  wire and_1956_tmp;
  wire and_1986_tmp;
  wire and_2058_tmp;
  wire and_2121_tmp;
  wire and_2163_tmp;
  wire and_2166_tmp;
  wire and_1755_tmp;
  wire and_2115_tmp;
  wire and_1962_tmp;
  wire and_1473_tmp;
  wire and_2073_tmp;
  wire and_1659_tmp;
  wire and_1782_tmp;
  wire and_1464_tmp;
  wire and_1695_tmp;
  wire and_1875_tmp;
  wire and_2028_tmp;
  wire and_1419_tmp;
  wire and_1551_tmp;
  wire and_2130_tmp;
  wire and_1734_tmp;
  wire and_1671_tmp;
  wire and_1998_tmp;
  wire and_2094_tmp;
  wire and_1482_tmp;
  wire and_1848_tmp;
  wire and_1590_tmp;
  wire and_1881_tmp;
  wire and_1608_tmp;
  wire and_1737_tmp;
  wire and_1680_tmp;
  wire and_1950_tmp;
  wire and_2022_tmp;
  wire and_1785_tmp;
  wire and_1758_tmp;
  wire and_1683_tmp;
  wire and_1641_tmp;
  wire and_1689_tmp;
  wire and_1542_tmp;
  wire and_1440_tmp;
  wire and_2124_tmp;
  wire and_1797_tmp;
  wire and_1857_tmp;
  wire and_2106_tmp;
  wire and_2088_tmp;
  wire and_1902_tmp;
  wire and_2037_tmp;
  wire and_1809_tmp;
  wire and_2004_tmp;
  wire input_mem_banks_read_read_data_and_21_tmp;
  wire and_1728_tmp;
  wire and_1719_tmp;
  wire and_1890_tmp;
  wire and_1800_tmp;
  wire and_1566_tmp;
  wire and_1560_tmp;
  wire and_2139_tmp;
  wire and_2085_tmp;
  wire and_1779_tmp;
  wire and_1617_tmp;
  wire and_1524_tmp;
  wire and_1818_tmp;
  wire and_1935_tmp;
  wire and_1626_tmp;
  wire and_1743_tmp;
  wire and_1461_tmp;
  wire and_1896_tmp;
  wire and_1647_tmp;
  wire and_2142_tmp;
  wire and_1932_tmp;
  wire and_2019_tmp;
  wire and_1713_tmp;
  wire and_2118_tmp;
  wire and_1863_tmp;
  wire and_1731_tmp;
  wire and_1584_tmp;
  wire and_1788_tmp;
  wire and_1776_tmp;
  wire and_1824_tmp;
  wire and_1767_tmp;
  wire and_1803_tmp;
  wire and_2001_tmp;
  wire and_1509_tmp;
  wire and_1827_tmp;
  wire and_2184_tmp;
  wire and_2082_tmp;
  wire and_2151_tmp;
  wire and_1503_tmp;
  wire and_2112_tmp;
  wire and_1959_tmp;
  wire and_1854_tmp;
  wire and_1869_tmp;
  wire and_1707_tmp;
  wire and_1839_tmp;
  wire and_1443_tmp;
  wire and_1692_tmp;
  wire and_2025_tmp;
  wire and_1479_tmp;
  wire and_1926_tmp;
  wire and_1947_tmp;
  wire and_1893_tmp;
  wire and_1866_tmp;
  wire and_1860_tmp;
  wire and_1578_tmp;
  wire and_1506_tmp;
  wire and_1878_tmp;
  wire and_2175_tmp;
  wire and_1428_tmp;
  wire and_1725_tmp;
  wire and_1740_tmp;
  wire and_1446_tmp;
  wire and_1830_tmp;
  wire and_1764_tmp;
  wire and_1929_tmp;
  wire and_2052_tmp;
  wire and_1449_tmp;
  wire and_2010_tmp;
  wire and_1611_tmp;
  wire and_1917_tmp;
  wire and_1992_tmp;
  wire and_2013_tmp;
  wire and_1989_tmp;
  wire and_1434_tmp;
  wire and_1971_tmp;
  wire and_2064_tmp;
  wire and_1530_tmp;
  wire and_2160_tmp;
  wire and_1527_tmp;
  wire and_1845_tmp;
  wire and_1953_tmp;
  wire and_1638_tmp;
  wire and_1851_tmp;
  wire and_1485_tmp;
  wire and_1563_tmp;
  wire and_1587_tmp;
  wire and_1536_tmp;
  wire and_1593_tmp;
  wire and_1422_tmp;
  wire and_1704_tmp;
  wire and_1629_tmp;
  wire input_mem_banks_read_read_data_and_20_tmp;
  wire and_1217_tmp;
  wire mux_498_itm;
  wire PECore_PushAxiRsp_if_else_mux_14_itm;
  wire PECore_PushAxiRsp_if_else_mux_15_itm;
  wire PECore_PushAxiRsp_if_else_mux_16_itm;

  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_1;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_1;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_1;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_1;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_2;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_2;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_2;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_2;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_3;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_3;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_3;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_3;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_4;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_4;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_4;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_4;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_5;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_5;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_5;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_5;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_6;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_6;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_6;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_6;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_7;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_7;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_7;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_7;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_8;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_8;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_8;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_8;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_9;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_9;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_9;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_9;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_10;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_10;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_10;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_10;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_1;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_1;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_11;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_11;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_11;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_11;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_12;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_12;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_12;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_12;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_2;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_2;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_13;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_13;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_13;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_13;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_14;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_14;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_14;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_14;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_3;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_3;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_15;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_15;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_15;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_15;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_16;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_16;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_16;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_16;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_4;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_4;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_17;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_17;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_17;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_17;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_18;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_18;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_18;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_18;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_5;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_5;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_19;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_19;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_19;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_19;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_20;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_20;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_20;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_20;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_6;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_6;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_21;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_21;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_21;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_21;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_22;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_22;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_22;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_22;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_7;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_7;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_23;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_23;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_23;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_23;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_24;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_24;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_24;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_24;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_8;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_8;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_25;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_25;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_25;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_25;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_26;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_26;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_26;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_26;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_9;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_9;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_27;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_27;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_27;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_27;
  wire mux_192_nl;
  wire and_486_nl;
  wire mux_191_nl;
  wire mux_190_nl;
  wire mux_189_nl;
  wire or_945_nl;
  wire or_944_nl;
  wire mux_197_nl;
  wire and_489_nl;
  wire mux_196_nl;
  wire mux_195_nl;
  wire mux_194_nl;
  wire or_951_nl;
  wire or_950_nl;
  wire mux_203_nl;
  wire and_493_nl;
  wire mux_202_nl;
  wire or_959_nl;
  wire mux_201_nl;
  wire mux_200_nl;
  wire or_958_nl;
  wire mux_198_nl;
  wire or_956_nl;
  wire or_955_nl;
  wire mux_209_nl;
  wire and_497_nl;
  wire mux_208_nl;
  wire or_966_nl;
  wire mux_207_nl;
  wire mux_206_nl;
  wire or_965_nl;
  wire mux_204_nl;
  wire or_963_nl;
  wire or_962_nl;
  wire mux_215_nl;
  wire and_501_nl;
  wire mux_214_nl;
  wire mux_213_nl;
  wire mux_212_nl;
  wire or_972_nl;
  wire mux_210_nl;
  wire or_971_nl;
  wire or_970_nl;
  wire mux_221_nl;
  wire and_505_nl;
  wire mux_220_nl;
  wire or_979_nl;
  wire mux_219_nl;
  wire mux_218_nl;
  wire or_978_nl;
  wire mux_216_nl;
  wire or_976_nl;
  wire or_975_nl;
  wire mux_227_nl;
  wire and_509_nl;
  wire mux_226_nl;
  wire or_985_nl;
  wire mux_225_nl;
  wire mux_224_nl;
  wire or_984_nl;
  wire mux_222_nl;
  wire or_982_nl;
  wire or_981_nl;
  wire mux_234_nl;
  wire and_513_nl;
  wire mux_233_nl;
  wire or_992_nl;
  wire mux_232_nl;
  wire mux_231_nl;
  wire or_991_nl;
  wire mux_228_nl;
  wire or_988_nl;
  wire or_987_nl;
  wire nor_19_nl;
  wire and_985_nl;
  wire and_705_nl;
  wire mux_245_nl;
  wire mux_244_nl;
  wire mux_243_nl;
  wire and_709_nl;
  wire mux_239_nl;
  wire mux_242_nl;
  wire mux_241_nl;
  wire mux_240_nl;
  wire mux_493_nl;
  wire or_997_nl;
  wire or_996_nl;
  wire mux_248_nl;
  wire mux_247_nl;
  wire or_995_nl;
  wire or_994_nl;
  wire[30:0] PECore_RunScale_if_for_8_mul_1_nl;
  wire signed [31:0] nl_PECore_RunScale_if_for_8_mul_1_nl;
  wire[30:0] PECore_RunScale_if_for_1_mul_1_nl;
  wire signed [31:0] nl_PECore_RunScale_if_for_1_mul_1_nl;
  wire[30:0] PECore_RunScale_if_for_7_mul_1_nl;
  wire signed [31:0] nl_PECore_RunScale_if_for_7_mul_1_nl;
  wire[30:0] PECore_RunScale_if_for_2_mul_1_nl;
  wire signed [31:0] nl_PECore_RunScale_if_for_2_mul_1_nl;
  wire[30:0] PECore_RunScale_if_for_6_mul_1_nl;
  wire signed [31:0] nl_PECore_RunScale_if_for_6_mul_1_nl;
  wire[30:0] PECore_RunScale_if_for_3_mul_1_nl;
  wire signed [31:0] nl_PECore_RunScale_if_for_3_mul_1_nl;
  wire[30:0] PECore_RunScale_if_for_5_mul_1_nl;
  wire signed [31:0] nl_PECore_RunScale_if_for_5_mul_1_nl;
  wire[30:0] PECore_RunScale_if_for_4_mul_1_nl;
  wire signed [31:0] nl_PECore_RunScale_if_for_4_mul_1_nl;
  wire mux_5_nl;
  wire mux_4_nl;
  wire or_14_nl;
  wire mux_6_nl;
  wire mux_7_nl;
  wire or_21_nl;
  wire mux_9_nl;
  wire or_22_nl;
  wire mux_8_nl;
  wire weight_mem_run_3_for_5_and_100_nl;
  wire mux_500_nl;
  wire mux_505_nl;
  wire mux_504_nl;
  wire mux_10_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_20_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_6_nl;
  wire mux_512_nl;
  wire or_1485_nl;
  wire mux_511_nl;
  wire or_1483_nl;
  wire or_1466_nl;
  wire[7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_24_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_123_nl;
  wire mux_12_nl;
  wire nor_331_nl;
  wire[7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_40_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_109_nl;
  wire mux_13_nl;
  wire nor_332_nl;
  wire mux_14_nl;
  wire or_32_nl;
  wire or_31_nl;
  wire mux_15_nl;
  wire or_34_nl;
  wire or_33_nl;
  wire mux_16_nl;
  wire mux_514_nl;
  wire mux_513_nl;
  wire nor_900_nl;
  wire nor_901_nl;
  wire[10:0] PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_6_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_nl;
  wire[3:0] PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_and_nl;
  wire and_601_nl;
  wire[3:0] operator_4_false_acc_nl;
  wire[4:0] nl_operator_4_false_acc_nl;
  wire pe_config_UpdateManagerCounter_if_not_7_nl;
  wire mux_515_nl;
  wire mux_516_nl;
  wire[1:0] PECore_UpdateFSM_switch_lp_and_1_nl;
  wire[1:0] PECore_UpdateFSM_switch_lp_mux1h_18_nl;
  wire PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_or_nl;
  wire PECore_UpdateFSM_switch_lp_or_nl;
  wire PECore_UpdateFSM_switch_lp_nor_8_nl;
  wire mux_26_nl;
  wire mux_25_nl;
  wire mux_24_nl;
  wire mux_23_nl;
  wire mux_22_nl;
  wire mux_21_nl;
  wire mux_20_nl;
  wire nor_259_nl;
  wire nor_260_nl;
  wire nor_261_nl;
  wire nor_262_nl;
  wire nor_263_nl;
  wire nor_264_nl;
  wire nor_265_nl;
  wire nor_266_nl;
  wire[22:0] accum_vector_data_acc_29_nl;
  wire[23:0] nl_accum_vector_data_acc_29_nl;
  wire[22:0] accum_vector_data_mux_12_nl;
  wire[22:0] accum_vector_data_mux_9_nl;
  wire[22:0] accum_vector_data_acc_9_nl;
  wire[23:0] nl_accum_vector_data_acc_9_nl;
  wire[22:0] accum_vector_data_mux_54_nl;
  wire[22:0] accum_vector_data_mux_51_nl;
  wire[22:0] accum_vector_data_acc_27_nl;
  wire[23:0] nl_accum_vector_data_acc_27_nl;
  wire[22:0] accum_vector_data_mux_17_nl;
  wire[22:0] accum_vector_data_mux_14_nl;
  wire[22:0] accum_vector_data_acc_12_nl;
  wire[23:0] nl_accum_vector_data_acc_12_nl;
  wire[22:0] accum_vector_data_mux_48_nl;
  wire[22:0] accum_vector_data_mux_45_nl;
  wire[22:0] accum_vector_data_acc_24_nl;
  wire[23:0] nl_accum_vector_data_acc_24_nl;
  wire[22:0] accum_vector_data_mux_21_nl;
  wire[22:0] accum_vector_data_mux_19_nl;
  wire[22:0] accum_vector_data_acc_15_nl;
  wire[23:0] nl_accum_vector_data_acc_15_nl;
  wire[22:0] accum_vector_data_mux_42_nl;
  wire[22:0] accum_vector_data_mux_39_nl;
  wire[22:0] accum_vector_data_acc_16_nl;
  wire[23:0] nl_accum_vector_data_acc_16_nl;
  wire[22:0] accum_vector_data_mux_36_nl;
  wire[22:0] accum_vector_data_acc_21_nl;
  wire[23:0] nl_accum_vector_data_acc_21_nl;
  wire[22:0] accum_vector_data_mux_27_nl;
  wire[22:0] accum_vector_data_mux_24_nl;
  wire[22:0] accum_vector_data_acc_18_nl;
  wire[23:0] nl_accum_vector_data_acc_18_nl;
  wire[22:0] accum_vector_data_mux_33_nl;
  wire[22:0] accum_vector_data_mux_30_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_122_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_108_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_130_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_15_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_16_nl;
  wire[7:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_20_nl;
  wire[7:0] PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_and_1_nl;
  wire PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_mux_19_nl;
  wire PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_mux_6_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_1_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_7_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_and_16_nl;
  wire mux_31_nl;
  wire mux_30_nl;
  wire nor_338_nl;
  wire mux_531_nl;
  wire mux_536_nl;
  wire mux_535_nl;
  wire mux_534_nl;
  wire mux_533_nl;
  wire mux_532_nl;
  wire or_1608_nl;
  wire or_1605_nl;
  wire or_1603_nl;
  wire or_1601_nl;
  wire or_1599_nl;
  wire or_1597_nl;
  wire or_1595_nl;
  wire mux_538_nl;
  wire or_1593_nl;
  wire mux_544_nl;
  wire mux_543_nl;
  wire mux_542_nl;
  wire mux_541_nl;
  wire mux_540_nl;
  wire or_1627_nl;
  wire or_1624_nl;
  wire or_1622_nl;
  wire or_1620_nl;
  wire or_1618_nl;
  wire or_1616_nl;
  wire or_1614_nl;
  wire mux_546_nl;
  wire or_1612_nl;
  wire mux_552_nl;
  wire mux_551_nl;
  wire mux_550_nl;
  wire mux_549_nl;
  wire mux_548_nl;
  wire or_1647_nl;
  wire or_1644_nl;
  wire or_1642_nl;
  wire or_1640_nl;
  wire or_1638_nl;
  wire or_1636_nl;
  wire or_1634_nl;
  wire mux_554_nl;
  wire or_1632_nl;
  wire mux_560_nl;
  wire mux_559_nl;
  wire mux_558_nl;
  wire mux_557_nl;
  wire mux_556_nl;
  wire or_1665_nl;
  wire or_1662_nl;
  wire or_1660_nl;
  wire or_1658_nl;
  wire or_1656_nl;
  wire or_1654_nl;
  wire or_1652_nl;
  wire mux_562_nl;
  wire or_1650_nl;
  wire mux_576_nl;
  wire mux_575_nl;
  wire mux_574_nl;
  wire mux_573_nl;
  wire mux_572_nl;
  wire or_1701_nl;
  wire or_1698_nl;
  wire or_1696_nl;
  wire or_1694_nl;
  wire or_1692_nl;
  wire or_1690_nl;
  wire or_1688_nl;
  wire mux_578_nl;
  wire or_1686_nl;
  wire mux_594_nl;
  wire mux_593_nl;
  wire mux_592_nl;
  wire mux_591_nl;
  wire mux_590_nl;
  wire mux_589_nl;
  wire mux_588_nl;
  wire or_1737_nl;
  wire or_1734_nl;
  wire or_1732_nl;
  wire or_1730_nl;
  wire or_1728_nl;
  wire or_1726_nl;
  wire or_1724_nl;
  wire or_1722_nl;
  wire mux_616_nl;
  wire mux_615_nl;
  wire mux_614_nl;
  wire mux_613_nl;
  wire mux_612_nl;
  wire or_1791_nl;
  wire or_1788_nl;
  wire or_1786_nl;
  wire or_1784_nl;
  wire or_1782_nl;
  wire or_1780_nl;
  wire or_1778_nl;
  wire mux_618_nl;
  wire or_1776_nl;
  wire mux_632_nl;
  wire mux_631_nl;
  wire mux_630_nl;
  wire mux_629_nl;
  wire mux_628_nl;
  wire or_1827_nl;
  wire or_1824_nl;
  wire or_1822_nl;
  wire or_1820_nl;
  wire or_1818_nl;
  wire or_1816_nl;
  wire or_1814_nl;
  wire mux_634_nl;
  wire or_1812_nl;
  wire[22:0] accum_vector_data_mux_62_nl;
  wire[22:0] accum_vector_data_mux_59_nl;
  wire[22:0] accum_vector_data_mux_68_nl;
  wire[22:0] accum_vector_data_mux_65_nl;
  wire[22:0] accum_vector_data_mux_74_nl;
  wire[22:0] accum_vector_data_mux_71_nl;
  wire[22:0] accum_vector_data_mux_80_nl;
  wire[22:0] accum_vector_data_mux_77_nl;
  wire[22:0] accum_vector_data_mux_86_nl;
  wire[22:0] accum_vector_data_mux_83_nl;
  wire accum_vector_operator_1_for_not_13_nl;
  wire[22:0] accum_vector_data_mux_92_nl;
  wire[22:0] accum_vector_data_mux_89_nl;
  wire[22:0] accum_vector_data_mux_98_nl;
  wire[22:0] accum_vector_data_mux_95_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_131_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_103_nl;
  wire mux_103_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_117_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_124_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_96_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_110_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_132_nl;
  wire mux_108_nl;
  wire mux_107_nl;
  wire mux_106_nl;
  wire mux_105_nl;
  wire mux_104_nl;
  wire weight_mem_banks_load_store_for_else_mux1h_11_nl;
  wire[6:0] weight_mem_banks_load_store_for_else_mux1h_38_nl;
  wire not_2441_nl;
  wire mux_474_nl;
  wire[7:0] mux1h_2_nl;
  wire and_918_nl;
  wire and_919_nl;
  wire and_612_nl;
  wire not_2450_nl;
  wire mux_110_nl;
  wire mux_109_nl;
  wire nor_350_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_125_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_111_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_133_nl;
  wire[3:0] weight_mem_banks_load_store_for_else_mux1h_18_nl;
  wire not_2442_nl;
  wire[3:0] weight_mem_banks_load_store_for_else_mux1h_39_nl;
  wire not_2443_nl;
  wire[7:0] mux_489_nl;
  wire[7:0] weight_mem_banks_load_store_for_else_or_nl;
  wire[7:0] weight_mem_banks_load_store_for_else_mux1h_20_nl;
  wire and_613_nl;
  wire and_615_nl;
  wire and_619_nl;
  wire and_623_nl;
  wire and_624_nl;
  wire and_616_nl;
  wire or_1404_nl;
  wire nor_522_nl;
  wire mux_475_nl;
  wire or_1402_nl;
  wire mux_117_nl;
  wire mux_116_nl;
  wire mux_115_nl;
  wire mux_114_nl;
  wire mux_113_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_126_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_112_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_134_nl;
  wire mux_120_nl;
  wire nor_291_nl;
  wire mux_119_nl;
  wire mux_118_nl;
  wire[1:0] weight_mem_banks_load_store_for_else_mux1h_25_nl;
  wire not_2444_nl;
  wire[5:0] weight_mem_banks_load_store_for_else_mux1h_40_nl;
  wire not_2445_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_127_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_113_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_135_nl;
  wire weight_mem_banks_load_store_for_else_mux1h_30_nl;
  wire[6:0] weight_mem_banks_load_store_for_else_mux1h_41_nl;
  wire not_2447_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_128_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_114_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_78_nl;
  wire mux_121_nl;
  wire weight_mem_banks_load_store_for_else_mux1h_35_nl;
  wire[6:0] weight_mem_banks_load_store_for_else_mux1h_42_nl;
  wire not_2449_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_76_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_72_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_and_7_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_and_9_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_14_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_4_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_for_and_5_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_28_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_35_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_34_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_nl;
  wire mux_122_nl;
  wire mux_123_nl;
  wire and_698_nl;
  wire mux_173_nl;
  wire nor_353_nl;
  wire[63:0] input_mem_banks_read_1_for_mux_4_nl;
  wire and_629_nl;
  wire weight_port_read_out_data_mux_20_nl;
  wire[7:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_1_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_129_nl;
  wire nor_963_nl;
  wire nor_1000_nl;
  wire nor_1001_nl;
  wire or_2278_nl;
  wire or_2276_nl;
  wire while_if_while_if_and_12_nl;
  wire mux_176_nl;
  wire[14:0] while_if_while_if_and_2_nl;
  wire mux_278_nl;
  wire or_1095_nl;
  wire mux_277_nl;
  wire and_649_nl;
  wire or_1096_nl;
  wire mux_177_nl;
  wire mux_180_nl;
  wire mux_179_nl;
  wire mux_178_nl;
  wire and_699_nl;
  wire or_921_nl;
  wire mux_184_nl;
  wire mux_183_nl;
  wire mux_182_nl;
  wire mux_181_nl;
  wire and_701_nl;
  wire or_923_nl;
  wire nor_354_nl;
  wire mux_185_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_nl;
  wire PECore_DecodeAxiRead_case_4_switch_lp_mux_2_nl;
  wire PECore_DecodeAxiRead_case_4_switch_lp_mux_3_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_1_nl;
  wire PECore_DecodeAxiRead_case_4_switch_lp_mux_7_nl;
  wire PECore_DecodeAxiRead_case_4_switch_lp_mux_8_nl;
  wire[3:0] PECore_DecodeAxiRead_case_4_switch_lp_mux_9_nl;
  wire[6:0] PECore_DecodeAxiRead_case_4_switch_lp_mux_10_nl;
  wire weight_mem_run_3_for_5_and_81_nl;
  wire weight_mem_run_3_for_5_and_7_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_56_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_57_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_58_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_59_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_60_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_61_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_62_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_63_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_64_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_65_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_66_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_67_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_69_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_70_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_71_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_72_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_100_nl;
  wire Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_101_nl;
  wire[14:0] PECore_RunFSM_case_2_for_2_operator_15_false_acc_nl;
  wire[15:0] nl_PECore_RunFSM_case_2_for_2_operator_15_false_acc_nl;
  wire[13:0] operator_15_false_acc_nl;
  wire[14:0] nl_operator_15_false_acc_nl;
  wire[14:0] PECore_RunFSM_case_2_for_4_operator_15_false_acc_nl;
  wire[15:0] nl_PECore_RunFSM_case_2_for_4_operator_15_false_acc_nl;
  wire[12:0] operator_15_false_acc_1_nl;
  wire[13:0] nl_operator_15_false_acc_1_nl;
  wire[14:0] PECore_RunFSM_case_2_for_6_operator_15_false_acc_nl;
  wire[15:0] nl_PECore_RunFSM_case_2_for_6_operator_15_false_acc_nl;
  wire[13:0] operator_15_false_acc_2_nl;
  wire[14:0] nl_operator_15_false_acc_2_nl;
  wire[14:0] PECore_RunFSM_case_2_for_8_operator_15_false_acc_nl;
  wire[15:0] nl_PECore_RunFSM_case_2_for_8_operator_15_false_acc_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_22_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_20_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_18_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_16_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_14_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_12_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_10_nl;
  wire Arbiter_8U_Roundrobin_pick_1_if_1_mux_8_nl;
  wire[7:0] pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_and_nl;
  wire[7:0] operator_8_false_acc_nl;
  wire[8:0] nl_operator_8_false_acc_nl;
  wire pe_config_UpdateInputCounter_not_nl;
  wire pe_config_input_counter_nand_nl;
  wire[7:0] pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_and_1_nl;
  wire[7:0] operator_8_false_1_acc_nl;
  wire[8:0] nl_operator_8_false_1_acc_nl;
  wire pe_config_UpdateManagerCounter_if_not_9_nl;
  wire pe_config_output_counter_nand_nl;
  wire while_and_63_nl;
  wire pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_and_nl;
  wire while_if_or_nl;
  wire while_if_and_4_nl;
  wire[19:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_15_nl;
  wire PECore_UpdateFSM_switch_lp_not_23_nl;
  wire[19:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_14_nl;
  wire PECore_UpdateFSM_switch_lp_not_24_nl;
  wire[19:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_13_nl;
  wire PECore_UpdateFSM_switch_lp_not_25_nl;
  wire[19:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_12_nl;
  wire PECore_UpdateFSM_switch_lp_not_26_nl;
  wire[19:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_11_nl;
  wire PECore_UpdateFSM_switch_lp_not_27_nl;
  wire[19:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_10_nl;
  wire PECore_UpdateFSM_switch_lp_not_28_nl;
  wire[19:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_9_nl;
  wire PECore_UpdateFSM_switch_lp_not_29_nl;
  wire[19:0] PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_8_nl;
  wire PECore_UpdateFSM_switch_lp_not_19_nl;
  wire[22:0] ProductSum_for_mux_nl;
  wire accum_vector_operator_1_for_not_61_nl;
  wire[22:0] ProductSum_for_mux_1_nl;
  wire accum_vector_operator_1_for_not_38_nl;
  wire[22:0] ProductSum_for_mux_2_nl;
  wire accum_vector_operator_1_for_not_62_nl;
  wire[22:0] ProductSum_for_mux_3_nl;
  wire accum_vector_operator_1_for_not_40_nl;
  wire[22:0] ProductSum_for_mux_4_nl;
  wire accum_vector_operator_1_for_not_63_nl;
  wire[22:0] ProductSum_for_mux_5_nl;
  wire accum_vector_operator_1_for_not_42_nl;
  wire[22:0] ProductSum_for_mux_6_nl;
  wire accum_vector_operator_1_for_not_64_nl;
  wire[22:0] ProductSum_for_mux_7_nl;
  wire accum_vector_operator_1_for_not_44_nl;
  wire[22:0] ProductSum_for_mux_8_nl;
  wire accum_vector_operator_1_for_not_65_nl;
  wire[22:0] ProductSum_for_mux_9_nl;
  wire accum_vector_operator_1_for_not_46_nl;
  wire[22:0] ProductSum_for_mux_10_nl;
  wire accum_vector_operator_1_for_not_66_nl;
  wire[22:0] ProductSum_for_mux_11_nl;
  wire accum_vector_operator_1_for_not_67_nl;
  wire[22:0] ProductSum_for_mux_12_nl;
  wire accum_vector_operator_1_for_not_48_nl;
  wire[22:0] ProductSum_for_mux_13_nl;
  wire accum_vector_operator_1_for_not_68_nl;
  wire[22:0] ProductSum_for_mux_14_nl;
  wire accum_vector_operator_1_for_not_50_nl;
  wire[22:0] ProductSum_for_mux_15_nl;
  wire accum_vector_operator_1_for_not_69_nl;
  wire[22:0] ProductSum_for_mux_16_nl;
  wire accum_vector_operator_1_for_not_52_nl;
  wire[22:0] ProductSum_for_mux_24_nl;
  wire accum_vector_operator_1_for_not_54_nl;
  wire[22:0] ProductSum_for_mux_25_nl;
  wire accum_vector_operator_1_for_not_24_nl;
  wire[22:0] ProductSum_for_mux_26_nl;
  wire accum_vector_operator_1_for_not_55_nl;
  wire[22:0] ProductSum_for_mux_27_nl;
  wire accum_vector_operator_1_for_not_26_nl;
  wire[22:0] ProductSum_for_mux_28_nl;
  wire accum_vector_operator_1_for_not_56_nl;
  wire[22:0] ProductSum_for_mux_29_nl;
  wire accum_vector_operator_1_for_not_28_nl;
  wire[22:0] ProductSum_for_mux_30_nl;
  wire accum_vector_operator_1_for_not_57_nl;
  wire[22:0] ProductSum_for_mux_31_nl;
  wire accum_vector_operator_1_for_not_30_nl;
  wire[22:0] ProductSum_for_mux_32_nl;
  wire accum_vector_operator_1_for_not_58_nl;
  wire[22:0] ProductSum_for_mux_33_nl;
  wire accum_vector_operator_1_for_not_32_nl;
  wire[22:0] ProductSum_for_mux_34_nl;
  wire accum_vector_operator_1_for_not_59_nl;
  wire[22:0] ProductSum_for_mux_35_nl;
  wire accum_vector_operator_1_for_not_34_nl;
  wire[22:0] ProductSum_for_mux_36_nl;
  wire accum_vector_operator_1_for_not_60_nl;
  wire[22:0] ProductSum_for_mux_37_nl;
  wire accum_vector_operator_1_for_not_36_nl;
  wire PECore_PushAxiRsp_mux_23_nl;
  wire mux1h_3_nl;
  wire[6:0] mux1h_10_nl;
  wire not_2545_nl;
  wire mux1h_4_nl;
  wire[6:0] mux1h_11_nl;
  wire not_2546_nl;
  wire mux1h_5_nl;
  wire mux1h_12_nl;
  wire[5:0] mux1h_13_nl;
  wire not_2547_nl;
  wire mux1h_6_nl;
  wire[2:0] mux1h_14_nl;
  wire not_2549_nl;
  wire[3:0] mux1h_15_nl;
  wire not_2550_nl;
  wire input_mem_banks_bank_a_nand_nl;
  wire while_and_100_nl;
  wire while_and_101_nl;
  wire input_mem_banks_bank_a_nand_1_nl;
  wire while_and_104_nl;
  wire while_and_105_nl;
  wire input_mem_banks_bank_a_nand_2_nl;
  wire while_and_108_nl;
  wire while_and_109_nl;
  wire input_mem_banks_bank_a_nand_3_nl;
  wire while_and_112_nl;
  wire while_and_113_nl;
  wire input_mem_banks_bank_a_nand_4_nl;
  wire while_and_116_nl;
  wire while_and_117_nl;
  wire input_mem_banks_bank_a_nand_5_nl;
  wire while_and_120_nl;
  wire while_and_121_nl;
  wire input_mem_banks_bank_a_nand_6_nl;
  wire while_and_124_nl;
  wire while_and_125_nl;
  wire input_mem_banks_bank_a_nand_7_nl;
  wire while_and_128_nl;
  wire while_and_129_nl;
  wire input_mem_banks_bank_a_nand_8_nl;
  wire while_and_132_nl;
  wire while_and_133_nl;
  wire input_mem_banks_bank_a_nand_9_nl;
  wire while_and_136_nl;
  wire while_and_137_nl;
  wire input_mem_banks_bank_a_nand_10_nl;
  wire while_and_140_nl;
  wire while_and_141_nl;
  wire input_mem_banks_bank_a_nand_11_nl;
  wire while_and_144_nl;
  wire while_and_145_nl;
  wire input_mem_banks_bank_a_nand_12_nl;
  wire while_and_148_nl;
  wire while_and_149_nl;
  wire input_mem_banks_bank_a_nand_13_nl;
  wire while_and_152_nl;
  wire while_and_153_nl;
  wire input_mem_banks_bank_a_nand_14_nl;
  wire while_and_156_nl;
  wire while_and_157_nl;
  wire input_mem_banks_bank_a_nand_15_nl;
  wire while_and_160_nl;
  wire while_and_161_nl;
  wire input_mem_banks_bank_a_nand_16_nl;
  wire while_and_164_nl;
  wire while_and_165_nl;
  wire input_mem_banks_bank_a_nand_17_nl;
  wire while_and_168_nl;
  wire while_and_169_nl;
  wire input_mem_banks_bank_a_nand_18_nl;
  wire while_and_172_nl;
  wire while_and_173_nl;
  wire input_mem_banks_bank_a_nand_19_nl;
  wire while_and_176_nl;
  wire while_and_177_nl;
  wire input_mem_banks_bank_a_nand_20_nl;
  wire while_and_180_nl;
  wire while_and_181_nl;
  wire input_mem_banks_bank_a_nand_21_nl;
  wire while_and_184_nl;
  wire while_and_185_nl;
  wire input_mem_banks_bank_a_nand_22_nl;
  wire while_and_188_nl;
  wire while_and_189_nl;
  wire input_mem_banks_bank_a_nand_23_nl;
  wire while_and_192_nl;
  wire while_and_193_nl;
  wire input_mem_banks_bank_a_nand_24_nl;
  wire while_and_196_nl;
  wire while_and_197_nl;
  wire input_mem_banks_bank_a_nand_25_nl;
  wire while_and_200_nl;
  wire while_and_201_nl;
  wire input_mem_banks_bank_a_nand_26_nl;
  wire while_and_204_nl;
  wire while_and_205_nl;
  wire input_mem_banks_bank_a_nand_27_nl;
  wire while_and_208_nl;
  wire while_and_209_nl;
  wire input_mem_banks_bank_a_nand_28_nl;
  wire while_and_212_nl;
  wire while_and_213_nl;
  wire input_mem_banks_bank_a_nand_29_nl;
  wire while_and_216_nl;
  wire while_and_217_nl;
  wire input_mem_banks_bank_a_nand_30_nl;
  wire while_and_220_nl;
  wire while_and_221_nl;
  wire input_mem_banks_bank_a_nand_31_nl;
  wire while_and_224_nl;
  wire while_and_225_nl;
  wire input_mem_banks_bank_a_nand_32_nl;
  wire while_and_228_nl;
  wire while_and_229_nl;
  wire input_mem_banks_bank_a_nand_33_nl;
  wire while_and_232_nl;
  wire while_and_233_nl;
  wire input_mem_banks_bank_a_nand_34_nl;
  wire while_and_236_nl;
  wire while_and_237_nl;
  wire input_mem_banks_bank_a_nand_35_nl;
  wire while_and_240_nl;
  wire while_and_241_nl;
  wire input_mem_banks_bank_a_nand_36_nl;
  wire while_and_244_nl;
  wire while_and_245_nl;
  wire input_mem_banks_bank_a_nand_37_nl;
  wire while_and_248_nl;
  wire while_and_249_nl;
  wire input_mem_banks_bank_a_nand_38_nl;
  wire while_and_252_nl;
  wire while_and_253_nl;
  wire input_mem_banks_bank_a_nand_39_nl;
  wire while_and_256_nl;
  wire while_and_257_nl;
  wire input_mem_banks_bank_a_nand_40_nl;
  wire while_and_260_nl;
  wire while_and_261_nl;
  wire input_mem_banks_bank_a_nand_41_nl;
  wire while_and_264_nl;
  wire while_and_265_nl;
  wire input_mem_banks_bank_a_nand_42_nl;
  wire while_and_268_nl;
  wire while_and_269_nl;
  wire input_mem_banks_bank_a_nand_43_nl;
  wire while_and_272_nl;
  wire while_and_273_nl;
  wire input_mem_banks_bank_a_nand_44_nl;
  wire while_and_276_nl;
  wire while_and_277_nl;
  wire input_mem_banks_bank_a_nand_45_nl;
  wire while_and_280_nl;
  wire while_and_281_nl;
  wire input_mem_banks_bank_a_nand_46_nl;
  wire while_and_284_nl;
  wire while_and_285_nl;
  wire input_mem_banks_bank_a_nand_47_nl;
  wire while_and_288_nl;
  wire while_and_289_nl;
  wire input_mem_banks_bank_a_nand_48_nl;
  wire while_and_292_nl;
  wire while_and_293_nl;
  wire input_mem_banks_bank_a_nand_49_nl;
  wire while_and_296_nl;
  wire while_and_297_nl;
  wire input_mem_banks_bank_a_nand_50_nl;
  wire while_and_300_nl;
  wire while_and_301_nl;
  wire input_mem_banks_bank_a_nand_51_nl;
  wire while_and_304_nl;
  wire while_and_305_nl;
  wire input_mem_banks_bank_a_nand_52_nl;
  wire while_and_308_nl;
  wire while_and_309_nl;
  wire input_mem_banks_bank_a_nand_53_nl;
  wire while_and_312_nl;
  wire while_and_313_nl;
  wire input_mem_banks_bank_a_nand_54_nl;
  wire while_and_316_nl;
  wire while_and_317_nl;
  wire input_mem_banks_bank_a_nand_55_nl;
  wire while_and_320_nl;
  wire while_and_321_nl;
  wire input_mem_banks_bank_a_nand_56_nl;
  wire while_and_324_nl;
  wire while_and_325_nl;
  wire input_mem_banks_bank_a_nand_57_nl;
  wire while_and_328_nl;
  wire while_and_329_nl;
  wire input_mem_banks_bank_a_nand_58_nl;
  wire while_and_332_nl;
  wire while_and_333_nl;
  wire input_mem_banks_bank_a_nand_59_nl;
  wire while_and_336_nl;
  wire while_and_337_nl;
  wire input_mem_banks_bank_a_nand_60_nl;
  wire while_and_340_nl;
  wire while_and_341_nl;
  wire input_mem_banks_bank_a_nand_61_nl;
  wire while_and_344_nl;
  wire while_and_345_nl;
  wire input_mem_banks_bank_a_nand_62_nl;
  wire while_and_348_nl;
  wire while_and_349_nl;
  wire input_mem_banks_bank_a_nand_63_nl;
  wire while_and_352_nl;
  wire while_and_353_nl;
  wire input_mem_banks_bank_a_nand_64_nl;
  wire while_and_356_nl;
  wire while_and_357_nl;
  wire input_mem_banks_bank_a_nand_65_nl;
  wire while_and_360_nl;
  wire while_and_361_nl;
  wire input_mem_banks_bank_a_nand_66_nl;
  wire while_and_364_nl;
  wire while_and_365_nl;
  wire input_mem_banks_bank_a_nand_67_nl;
  wire while_and_368_nl;
  wire while_and_369_nl;
  wire input_mem_banks_bank_a_nand_68_nl;
  wire while_and_372_nl;
  wire while_and_373_nl;
  wire input_mem_banks_bank_a_nand_69_nl;
  wire while_and_376_nl;
  wire while_and_377_nl;
  wire input_mem_banks_bank_a_nand_70_nl;
  wire while_and_380_nl;
  wire while_and_381_nl;
  wire input_mem_banks_bank_a_nand_71_nl;
  wire while_and_384_nl;
  wire while_and_385_nl;
  wire input_mem_banks_bank_a_nand_72_nl;
  wire while_and_388_nl;
  wire while_and_389_nl;
  wire input_mem_banks_bank_a_nand_73_nl;
  wire while_and_392_nl;
  wire while_and_393_nl;
  wire input_mem_banks_bank_a_nand_74_nl;
  wire while_and_396_nl;
  wire while_and_397_nl;
  wire input_mem_banks_bank_a_nand_75_nl;
  wire while_and_400_nl;
  wire while_and_401_nl;
  wire input_mem_banks_bank_a_nand_76_nl;
  wire while_and_404_nl;
  wire while_and_405_nl;
  wire input_mem_banks_bank_a_nand_77_nl;
  wire while_and_408_nl;
  wire while_and_409_nl;
  wire input_mem_banks_bank_a_nand_78_nl;
  wire while_and_412_nl;
  wire while_and_413_nl;
  wire input_mem_banks_bank_a_nand_79_nl;
  wire while_and_416_nl;
  wire while_and_417_nl;
  wire input_mem_banks_bank_a_nand_80_nl;
  wire while_and_420_nl;
  wire while_and_421_nl;
  wire input_mem_banks_bank_a_nand_81_nl;
  wire while_and_424_nl;
  wire while_and_425_nl;
  wire input_mem_banks_bank_a_nand_82_nl;
  wire while_and_428_nl;
  wire while_and_429_nl;
  wire input_mem_banks_bank_a_nand_83_nl;
  wire while_and_432_nl;
  wire while_and_433_nl;
  wire input_mem_banks_bank_a_nand_84_nl;
  wire while_and_436_nl;
  wire while_and_437_nl;
  wire input_mem_banks_bank_a_nand_85_nl;
  wire while_and_440_nl;
  wire while_and_441_nl;
  wire input_mem_banks_bank_a_nand_86_nl;
  wire while_and_444_nl;
  wire while_and_445_nl;
  wire input_mem_banks_bank_a_nand_87_nl;
  wire while_and_448_nl;
  wire while_and_449_nl;
  wire input_mem_banks_bank_a_nand_88_nl;
  wire while_and_452_nl;
  wire while_and_453_nl;
  wire input_mem_banks_bank_a_nand_89_nl;
  wire while_and_456_nl;
  wire while_and_457_nl;
  wire input_mem_banks_bank_a_nand_90_nl;
  wire while_and_460_nl;
  wire while_and_461_nl;
  wire input_mem_banks_bank_a_nand_91_nl;
  wire while_and_464_nl;
  wire while_and_465_nl;
  wire input_mem_banks_bank_a_nand_92_nl;
  wire while_and_468_nl;
  wire while_and_469_nl;
  wire input_mem_banks_bank_a_nand_93_nl;
  wire while_and_472_nl;
  wire while_and_473_nl;
  wire input_mem_banks_bank_a_nand_94_nl;
  wire while_and_476_nl;
  wire while_and_477_nl;
  wire input_mem_banks_bank_a_nand_95_nl;
  wire while_and_480_nl;
  wire while_and_481_nl;
  wire input_mem_banks_bank_a_nand_96_nl;
  wire while_and_484_nl;
  wire while_and_485_nl;
  wire input_mem_banks_bank_a_nand_97_nl;
  wire while_and_488_nl;
  wire while_and_489_nl;
  wire input_mem_banks_bank_a_nand_98_nl;
  wire while_and_492_nl;
  wire while_and_493_nl;
  wire input_mem_banks_bank_a_nand_99_nl;
  wire while_and_496_nl;
  wire while_and_497_nl;
  wire input_mem_banks_bank_a_nand_100_nl;
  wire while_and_500_nl;
  wire while_and_501_nl;
  wire input_mem_banks_bank_a_nand_101_nl;
  wire while_and_504_nl;
  wire while_and_505_nl;
  wire input_mem_banks_bank_a_nand_102_nl;
  wire while_and_508_nl;
  wire while_and_509_nl;
  wire input_mem_banks_bank_a_nand_103_nl;
  wire while_and_512_nl;
  wire while_and_513_nl;
  wire input_mem_banks_bank_a_nand_104_nl;
  wire while_and_516_nl;
  wire while_and_517_nl;
  wire input_mem_banks_bank_a_nand_105_nl;
  wire while_and_520_nl;
  wire while_and_521_nl;
  wire input_mem_banks_bank_a_nand_106_nl;
  wire while_and_524_nl;
  wire while_and_525_nl;
  wire input_mem_banks_bank_a_nand_107_nl;
  wire while_and_528_nl;
  wire while_and_529_nl;
  wire input_mem_banks_bank_a_nand_108_nl;
  wire while_and_532_nl;
  wire while_and_533_nl;
  wire input_mem_banks_bank_a_nand_109_nl;
  wire while_and_536_nl;
  wire while_and_537_nl;
  wire input_mem_banks_bank_a_nand_110_nl;
  wire while_and_540_nl;
  wire while_and_541_nl;
  wire input_mem_banks_bank_a_nand_111_nl;
  wire while_and_544_nl;
  wire while_and_545_nl;
  wire input_mem_banks_bank_a_nand_112_nl;
  wire while_and_548_nl;
  wire while_and_549_nl;
  wire input_mem_banks_bank_a_nand_113_nl;
  wire while_and_552_nl;
  wire while_and_553_nl;
  wire input_mem_banks_bank_a_nand_114_nl;
  wire while_and_556_nl;
  wire while_and_557_nl;
  wire input_mem_banks_bank_a_nand_115_nl;
  wire while_and_560_nl;
  wire while_and_561_nl;
  wire input_mem_banks_bank_a_nand_116_nl;
  wire while_and_564_nl;
  wire while_and_565_nl;
  wire input_mem_banks_bank_a_nand_117_nl;
  wire while_and_568_nl;
  wire while_and_569_nl;
  wire input_mem_banks_bank_a_nand_118_nl;
  wire while_and_572_nl;
  wire while_and_573_nl;
  wire input_mem_banks_bank_a_nand_119_nl;
  wire while_and_576_nl;
  wire while_and_577_nl;
  wire input_mem_banks_bank_a_nand_120_nl;
  wire while_and_580_nl;
  wire while_and_581_nl;
  wire input_mem_banks_bank_a_nand_121_nl;
  wire while_and_584_nl;
  wire while_and_585_nl;
  wire input_mem_banks_bank_a_nand_122_nl;
  wire while_and_588_nl;
  wire while_and_589_nl;
  wire input_mem_banks_bank_a_nand_123_nl;
  wire while_and_592_nl;
  wire while_and_593_nl;
  wire input_mem_banks_bank_a_nand_124_nl;
  wire while_and_596_nl;
  wire while_and_597_nl;
  wire input_mem_banks_bank_a_nand_125_nl;
  wire while_and_600_nl;
  wire while_and_601_nl;
  wire input_mem_banks_bank_a_nand_126_nl;
  wire while_and_604_nl;
  wire while_and_605_nl;
  wire input_mem_banks_bank_a_nand_127_nl;
  wire while_and_608_nl;
  wire while_and_609_nl;
  wire input_mem_banks_bank_a_nand_128_nl;
  wire while_and_612_nl;
  wire while_and_613_nl;
  wire input_mem_banks_bank_a_nand_129_nl;
  wire while_and_616_nl;
  wire while_and_617_nl;
  wire input_mem_banks_bank_a_nand_130_nl;
  wire while_and_620_nl;
  wire while_and_621_nl;
  wire input_mem_banks_bank_a_nand_131_nl;
  wire while_and_624_nl;
  wire while_and_625_nl;
  wire input_mem_banks_bank_a_nand_132_nl;
  wire while_and_628_nl;
  wire while_and_629_nl;
  wire input_mem_banks_bank_a_nand_133_nl;
  wire while_and_632_nl;
  wire while_and_633_nl;
  wire input_mem_banks_bank_a_nand_134_nl;
  wire while_and_636_nl;
  wire while_and_637_nl;
  wire input_mem_banks_bank_a_nand_135_nl;
  wire while_and_640_nl;
  wire while_and_641_nl;
  wire input_mem_banks_bank_a_nand_136_nl;
  wire while_and_644_nl;
  wire while_and_645_nl;
  wire input_mem_banks_bank_a_nand_137_nl;
  wire while_and_648_nl;
  wire while_and_649_nl;
  wire input_mem_banks_bank_a_nand_138_nl;
  wire while_and_652_nl;
  wire while_and_653_nl;
  wire input_mem_banks_bank_a_nand_139_nl;
  wire while_and_656_nl;
  wire while_and_657_nl;
  wire input_mem_banks_bank_a_nand_140_nl;
  wire while_and_660_nl;
  wire while_and_661_nl;
  wire input_mem_banks_bank_a_nand_141_nl;
  wire while_and_664_nl;
  wire while_and_665_nl;
  wire input_mem_banks_bank_a_nand_142_nl;
  wire while_and_668_nl;
  wire while_and_669_nl;
  wire input_mem_banks_bank_a_nand_143_nl;
  wire while_and_672_nl;
  wire while_and_673_nl;
  wire input_mem_banks_bank_a_nand_144_nl;
  wire while_and_676_nl;
  wire while_and_677_nl;
  wire input_mem_banks_bank_a_nand_145_nl;
  wire while_and_680_nl;
  wire while_and_681_nl;
  wire input_mem_banks_bank_a_nand_146_nl;
  wire while_and_684_nl;
  wire while_and_685_nl;
  wire input_mem_banks_bank_a_nand_147_nl;
  wire while_and_688_nl;
  wire while_and_689_nl;
  wire input_mem_banks_bank_a_nand_148_nl;
  wire while_and_692_nl;
  wire while_and_693_nl;
  wire input_mem_banks_bank_a_nand_149_nl;
  wire while_and_696_nl;
  wire while_and_697_nl;
  wire input_mem_banks_bank_a_nand_150_nl;
  wire while_and_700_nl;
  wire while_and_701_nl;
  wire input_mem_banks_bank_a_nand_151_nl;
  wire while_and_704_nl;
  wire while_and_705_nl;
  wire input_mem_banks_bank_a_nand_152_nl;
  wire while_and_708_nl;
  wire while_and_709_nl;
  wire input_mem_banks_bank_a_nand_153_nl;
  wire while_and_712_nl;
  wire while_and_713_nl;
  wire input_mem_banks_bank_a_nand_154_nl;
  wire while_and_716_nl;
  wire while_and_717_nl;
  wire input_mem_banks_bank_a_nand_155_nl;
  wire while_and_720_nl;
  wire while_and_721_nl;
  wire input_mem_banks_bank_a_nand_156_nl;
  wire while_and_724_nl;
  wire while_and_725_nl;
  wire input_mem_banks_bank_a_nand_157_nl;
  wire while_and_728_nl;
  wire while_and_729_nl;
  wire input_mem_banks_bank_a_nand_158_nl;
  wire while_and_732_nl;
  wire while_and_733_nl;
  wire input_mem_banks_bank_a_nand_159_nl;
  wire while_and_736_nl;
  wire while_and_737_nl;
  wire input_mem_banks_bank_a_nand_160_nl;
  wire while_and_740_nl;
  wire while_and_741_nl;
  wire input_mem_banks_bank_a_nand_161_nl;
  wire while_and_744_nl;
  wire while_and_745_nl;
  wire input_mem_banks_bank_a_nand_162_nl;
  wire while_and_748_nl;
  wire while_and_749_nl;
  wire input_mem_banks_bank_a_nand_163_nl;
  wire while_and_752_nl;
  wire while_and_753_nl;
  wire input_mem_banks_bank_a_nand_164_nl;
  wire while_and_756_nl;
  wire while_and_757_nl;
  wire input_mem_banks_bank_a_nand_165_nl;
  wire while_and_760_nl;
  wire while_and_761_nl;
  wire input_mem_banks_bank_a_nand_166_nl;
  wire while_and_764_nl;
  wire while_and_765_nl;
  wire input_mem_banks_bank_a_nand_167_nl;
  wire while_and_768_nl;
  wire while_and_769_nl;
  wire input_mem_banks_bank_a_nand_168_nl;
  wire while_and_772_nl;
  wire while_and_773_nl;
  wire input_mem_banks_bank_a_nand_169_nl;
  wire while_and_776_nl;
  wire while_and_777_nl;
  wire input_mem_banks_bank_a_nand_170_nl;
  wire while_and_780_nl;
  wire while_and_781_nl;
  wire input_mem_banks_bank_a_nand_171_nl;
  wire while_and_784_nl;
  wire while_and_785_nl;
  wire input_mem_banks_bank_a_nand_172_nl;
  wire while_and_788_nl;
  wire while_and_789_nl;
  wire input_mem_banks_bank_a_nand_173_nl;
  wire while_and_792_nl;
  wire while_and_793_nl;
  wire input_mem_banks_bank_a_nand_174_nl;
  wire while_and_796_nl;
  wire while_and_797_nl;
  wire input_mem_banks_bank_a_nand_175_nl;
  wire while_and_800_nl;
  wire while_and_801_nl;
  wire input_mem_banks_bank_a_nand_176_nl;
  wire while_and_804_nl;
  wire while_and_805_nl;
  wire input_mem_banks_bank_a_nand_177_nl;
  wire while_and_808_nl;
  wire while_and_809_nl;
  wire input_mem_banks_bank_a_nand_178_nl;
  wire while_and_812_nl;
  wire while_and_813_nl;
  wire input_mem_banks_bank_a_nand_179_nl;
  wire while_and_816_nl;
  wire while_and_817_nl;
  wire input_mem_banks_bank_a_nand_180_nl;
  wire while_and_820_nl;
  wire while_and_821_nl;
  wire input_mem_banks_bank_a_nand_181_nl;
  wire while_and_824_nl;
  wire while_and_825_nl;
  wire input_mem_banks_bank_a_nand_182_nl;
  wire while_and_828_nl;
  wire while_and_829_nl;
  wire input_mem_banks_bank_a_nand_183_nl;
  wire while_and_832_nl;
  wire while_and_833_nl;
  wire input_mem_banks_bank_a_nand_184_nl;
  wire while_and_836_nl;
  wire while_and_837_nl;
  wire input_mem_banks_bank_a_nand_185_nl;
  wire while_and_840_nl;
  wire while_and_841_nl;
  wire input_mem_banks_bank_a_nand_186_nl;
  wire while_and_844_nl;
  wire while_and_845_nl;
  wire input_mem_banks_bank_a_nand_187_nl;
  wire while_and_848_nl;
  wire while_and_849_nl;
  wire input_mem_banks_bank_a_nand_188_nl;
  wire while_and_852_nl;
  wire while_and_853_nl;
  wire input_mem_banks_bank_a_nand_189_nl;
  wire while_and_856_nl;
  wire while_and_857_nl;
  wire input_mem_banks_bank_a_nand_190_nl;
  wire while_and_860_nl;
  wire while_and_861_nl;
  wire input_mem_banks_bank_a_nand_191_nl;
  wire while_and_864_nl;
  wire while_and_865_nl;
  wire input_mem_banks_bank_a_nand_192_nl;
  wire while_and_868_nl;
  wire while_and_869_nl;
  wire input_mem_banks_bank_a_nand_193_nl;
  wire while_and_872_nl;
  wire while_and_873_nl;
  wire input_mem_banks_bank_a_nand_194_nl;
  wire while_and_876_nl;
  wire while_and_877_nl;
  wire input_mem_banks_bank_a_nand_195_nl;
  wire while_and_880_nl;
  wire while_and_881_nl;
  wire input_mem_banks_bank_a_nand_196_nl;
  wire while_and_884_nl;
  wire while_and_885_nl;
  wire input_mem_banks_bank_a_nand_197_nl;
  wire while_and_888_nl;
  wire while_and_889_nl;
  wire input_mem_banks_bank_a_nand_198_nl;
  wire while_and_892_nl;
  wire while_and_893_nl;
  wire input_mem_banks_bank_a_nand_199_nl;
  wire while_and_896_nl;
  wire while_and_897_nl;
  wire input_mem_banks_bank_a_nand_200_nl;
  wire while_and_900_nl;
  wire while_and_901_nl;
  wire input_mem_banks_bank_a_nand_201_nl;
  wire while_and_904_nl;
  wire while_and_905_nl;
  wire input_mem_banks_bank_a_nand_202_nl;
  wire while_and_908_nl;
  wire while_and_909_nl;
  wire input_mem_banks_bank_a_nand_203_nl;
  wire while_and_912_nl;
  wire while_and_913_nl;
  wire input_mem_banks_bank_a_nand_204_nl;
  wire while_and_916_nl;
  wire while_and_917_nl;
  wire input_mem_banks_bank_a_nand_205_nl;
  wire while_and_920_nl;
  wire while_and_921_nl;
  wire input_mem_banks_bank_a_nand_206_nl;
  wire while_and_924_nl;
  wire while_and_925_nl;
  wire input_mem_banks_bank_a_nand_207_nl;
  wire while_and_928_nl;
  wire while_and_929_nl;
  wire input_mem_banks_bank_a_nand_208_nl;
  wire while_and_932_nl;
  wire while_and_933_nl;
  wire input_mem_banks_bank_a_nand_209_nl;
  wire while_and_936_nl;
  wire while_and_937_nl;
  wire input_mem_banks_bank_a_nand_210_nl;
  wire while_and_940_nl;
  wire while_and_941_nl;
  wire input_mem_banks_bank_a_nand_211_nl;
  wire while_and_944_nl;
  wire while_and_945_nl;
  wire input_mem_banks_bank_a_nand_212_nl;
  wire while_and_948_nl;
  wire while_and_949_nl;
  wire input_mem_banks_bank_a_nand_213_nl;
  wire while_and_952_nl;
  wire while_and_953_nl;
  wire input_mem_banks_bank_a_nand_214_nl;
  wire while_and_956_nl;
  wire while_and_957_nl;
  wire input_mem_banks_bank_a_nand_215_nl;
  wire while_and_960_nl;
  wire while_and_961_nl;
  wire input_mem_banks_bank_a_nand_216_nl;
  wire while_and_964_nl;
  wire while_and_965_nl;
  wire input_mem_banks_bank_a_nand_217_nl;
  wire while_and_968_nl;
  wire while_and_969_nl;
  wire input_mem_banks_bank_a_nand_218_nl;
  wire while_and_972_nl;
  wire while_and_973_nl;
  wire input_mem_banks_bank_a_nand_219_nl;
  wire while_and_976_nl;
  wire while_and_977_nl;
  wire input_mem_banks_bank_a_nand_220_nl;
  wire while_and_980_nl;
  wire while_and_981_nl;
  wire input_mem_banks_bank_a_nand_221_nl;
  wire while_and_984_nl;
  wire while_and_985_nl;
  wire input_mem_banks_bank_a_nand_222_nl;
  wire while_and_988_nl;
  wire while_and_989_nl;
  wire input_mem_banks_bank_a_nand_223_nl;
  wire while_and_992_nl;
  wire while_and_993_nl;
  wire input_mem_banks_bank_a_nand_224_nl;
  wire while_and_996_nl;
  wire while_and_997_nl;
  wire input_mem_banks_bank_a_nand_225_nl;
  wire while_and_1000_nl;
  wire while_and_1001_nl;
  wire input_mem_banks_bank_a_nand_226_nl;
  wire while_and_1004_nl;
  wire while_and_1005_nl;
  wire input_mem_banks_bank_a_nand_227_nl;
  wire while_and_1008_nl;
  wire while_and_1009_nl;
  wire input_mem_banks_bank_a_nand_228_nl;
  wire while_and_1012_nl;
  wire while_and_1013_nl;
  wire input_mem_banks_bank_a_nand_229_nl;
  wire while_and_1016_nl;
  wire while_and_1017_nl;
  wire input_mem_banks_bank_a_nand_230_nl;
  wire while_and_1020_nl;
  wire while_and_1021_nl;
  wire input_mem_banks_bank_a_nand_231_nl;
  wire while_and_1024_nl;
  wire while_and_1025_nl;
  wire input_mem_banks_bank_a_nand_232_nl;
  wire while_and_1028_nl;
  wire while_and_1029_nl;
  wire input_mem_banks_bank_a_nand_233_nl;
  wire while_and_1032_nl;
  wire while_and_1033_nl;
  wire input_mem_banks_bank_a_nand_234_nl;
  wire while_and_1036_nl;
  wire while_and_1037_nl;
  wire input_mem_banks_bank_a_nand_235_nl;
  wire while_and_1040_nl;
  wire while_and_1041_nl;
  wire input_mem_banks_bank_a_nand_236_nl;
  wire while_and_1044_nl;
  wire while_and_1045_nl;
  wire input_mem_banks_bank_a_nand_237_nl;
  wire while_and_1048_nl;
  wire while_and_1049_nl;
  wire input_mem_banks_bank_a_nand_238_nl;
  wire while_and_1052_nl;
  wire while_and_1053_nl;
  wire input_mem_banks_bank_a_nand_239_nl;
  wire while_and_1056_nl;
  wire while_and_1057_nl;
  wire input_mem_banks_bank_a_nand_240_nl;
  wire while_and_1060_nl;
  wire while_and_1061_nl;
  wire input_mem_banks_bank_a_nand_241_nl;
  wire while_and_1064_nl;
  wire while_and_1065_nl;
  wire input_mem_banks_bank_a_nand_242_nl;
  wire while_and_1068_nl;
  wire while_and_1069_nl;
  wire input_mem_banks_bank_a_nand_243_nl;
  wire while_and_1072_nl;
  wire while_and_1073_nl;
  wire input_mem_banks_bank_a_nand_244_nl;
  wire while_and_1076_nl;
  wire while_and_1077_nl;
  wire input_mem_banks_bank_a_nand_245_nl;
  wire while_and_1080_nl;
  wire while_and_1081_nl;
  wire input_mem_banks_bank_a_nand_246_nl;
  wire while_and_1084_nl;
  wire while_and_1085_nl;
  wire input_mem_banks_bank_a_nand_247_nl;
  wire while_and_1088_nl;
  wire while_and_1089_nl;
  wire input_mem_banks_bank_a_nand_248_nl;
  wire while_and_1092_nl;
  wire while_and_1093_nl;
  wire input_mem_banks_bank_a_nand_249_nl;
  wire while_and_1096_nl;
  wire while_and_1097_nl;
  wire input_mem_banks_bank_a_nand_250_nl;
  wire while_and_1100_nl;
  wire while_and_1101_nl;
  wire input_mem_banks_bank_a_nand_251_nl;
  wire while_and_1104_nl;
  wire while_and_1105_nl;
  wire input_mem_banks_bank_a_nand_252_nl;
  wire while_and_1108_nl;
  wire while_and_1109_nl;
  wire input_mem_banks_bank_a_nand_253_nl;
  wire while_and_1112_nl;
  wire while_and_1113_nl;
  wire input_mem_banks_bank_a_nand_254_nl;
  wire while_and_1116_nl;
  wire while_and_1117_nl;
  wire input_mem_banks_bank_a_nand_255_nl;
  wire while_and_1120_nl;
  wire while_and_1121_nl;
  wire weight_mem_banks_load_store_1_for_else_else_and_nl;
  wire weight_mem_banks_load_store_1_for_else_else_or_nl;
  wire weight_mem_banks_load_store_1_for_else_else_and_4_nl;
  wire weight_mem_banks_load_store_1_for_else_else_and_6_nl;
  wire weight_mem_banks_load_store_1_for_else_else_and_8_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_81_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_89_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_8_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_1_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_3_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_4_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_5_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_8_operator_4_false_2_operator_4_false_2_or_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_8_operator_3_false_1_operator_3_false_1_or_nl;
  wire mux_316_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_9_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_1_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_7_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_2_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_9_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_10_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_11_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_2_operator_4_false_2_or_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_7_operator_3_false_1_operator_3_false_1_or_nl;
  wire mux_353_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_10_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_12_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_13_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_14_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_15_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_16_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_17_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_6_operator_3_false_1_operator_3_false_1_or_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_2_operator_4_false_2_or_nl;
  wire and_667_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_11_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_3_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_19_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_4_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_21_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_22_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_23_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_2_operator_4_false_2_or_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_5_operator_3_false_1_operator_3_false_1_or_nl;
  wire mux_388_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_12_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_5_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_25_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_6_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_27_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_28_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_29_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_2_operator_4_false_2_or_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_4_operator_3_false_1_operator_3_false_1_or_nl;
  wire mux_409_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_13_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_7_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_31_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_8_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_33_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_34_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_35_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_2_operator_4_false_2_or_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_3_operator_3_false_1_operator_3_false_1_or_nl;
  wire mux_430_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_14_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_9_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_37_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_10_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_39_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_40_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_41_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_2_operator_4_false_2_or_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_2_operator_3_false_1_operator_3_false_1_or_nl;
  wire mux_455_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_15_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_3_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_11_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_43_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_44_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_45_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_46_nl;
  wire nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_47_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_1_operator_3_false_1_operator_3_false_1_or_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_2_operator_4_false_2_or_nl;
  wire and_679_nl;
  wire mux_470_nl;
  wire PECore_UpdateFSM_switch_lp_mux1h_14_nl;
  wire PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_8_nl;
  wire PECore_UpdateFSM_case_1_if_PECore_UpdateFSM_case_1_if_and_nl;
  wire PECore_UpdateFSM_switch_lp_pe_config_UpdateManagerCounter_nand_nl;
  wire[7:0] crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_mux1h_34_nl;
  wire crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_21_nl;
  wire[3:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_54_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_136_nl;
  wire[3:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_62_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_137_nl;
  wire[3:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_64_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_89_nl;
  wire[3:0] weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_65_nl;
  wire weight_mem_write_arbxbar_xbar_for_1_for_not_82_nl;
  wire mux1h_7_nl;
  wire[6:0] mux1h_16_nl;
  wire not_2551_nl;
  wire[3:0] mux1h_8_nl;
  wire not_2552_nl;
  wire[3:0] mux1h_17_nl;
  wire not_2463_nl;
  wire mux1h_9_nl;
  wire mux1h_18_nl;
  wire[5:0] mux1h_19_nl;
  wire not_2553_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_600_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_601_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_602_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_603_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_604_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_605_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_606_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_607_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_608_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_609_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_610_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_611_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_612_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_613_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_614_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_615_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_616_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_617_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_618_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_619_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_620_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_621_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_622_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_623_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_624_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_629_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_630_nl;
  wire mux_19_nl;
  wire or_120_nl;
  wire and_691_nl;
  wire or_117_nl;
  wire mux_28_nl;
  wire and_696_nl;
  wire or_187_nl;
  wire nor_288_nl;
  wire nor_289_nl;
  wire or_365_nl;
  wire nor_290_nl;
  wire mux_187_nl;
  wire nor_360_nl;
  wire nor_361_nl;
  wire mux_229_nl;
  wire mux_270_nl;
  wire or_1079_nl;
  wire mux_269_nl;
  wire or_1078_nl;
  wire nor_27_nl;
  wire mux_280_nl;
  wire mux_279_nl;
  wire or_1097_nl;
  wire mux_283_nl;
  wire mux_282_nl;
  wire or_1101_nl;
  wire or_1100_nl;
  wire mux_286_nl;
  wire mux_285_nl;
  wire nand_1_nl;
  wire nor_404_nl;
  wire nor_405_nl;
  wire mux_293_nl;
  wire mux_292_nl;
  wire mux_291_nl;
  wire mux_290_nl;
  wire mux_289_nl;
  wire nand_2_nl;
  wire mux_288_nl;
  wire or_1103_nl;
  wire mux_296_nl;
  wire or_1118_nl;
  wire mux_295_nl;
  wire or_1108_nl;
  wire or_1120_nl;
  wire or_1119_nl;
  wire mux_300_nl;
  wire or_1124_nl;
  wire or_1121_nl;
  wire mux_305_nl;
  wire mux_304_nl;
  wire mux_303_nl;
  wire mux_302_nl;
  wire or_1133_nl;
  wire mux_301_nl;
  wire or_1131_nl;
  wire or_1128_nl;
  wire or_1127_nl;
  wire mux_308_nl;
  wire mux_307_nl;
  wire or_1139_nl;
  wire or_1138_nl;
  wire or_1137_nl;
  wire or_1136_nl;
  wire mux_315_nl;
  wire mux_314_nl;
  wire mux_313_nl;
  wire mux_312_nl;
  wire mux_311_nl;
  wire mux_310_nl;
  wire or_1146_nl;
  wire or_1145_nl;
  wire or_1144_nl;
  wire or_1143_nl;
  wire or_1140_nl;
  wire or_1147_nl;
  wire or_1150_nl;
  wire mux_322_nl;
  wire mux_321_nl;
  wire mux_320_nl;
  wire or_1152_nl;
  wire mux_319_nl;
  wire or_1151_nl;
  wire or_1149_nl;
  wire or_1154_nl;
  wire or_1165_nl;
  wire mux_329_nl;
  wire mux_328_nl;
  wire mux_327_nl;
  wire or_1167_nl;
  wire mux_326_nl;
  wire or_1166_nl;
  wire or_1160_nl;
  wire or_1168_nl;
  wire or_1173_nl;
  wire or_1175_nl;
  wire mux_333_nl;
  wire or_1174_nl;
  wire or_1171_nl;
  wire mux_335_nl;
  wire or_1178_nl;
  wire or_1176_nl;
  wire mux_342_nl;
  wire mux_341_nl;
  wire mux_340_nl;
  wire mux_339_nl;
  wire mux_338_nl;
  wire or_1182_nl;
  wire or_1180_nl;
  wire or_1179_nl;
  wire mux_345_nl;
  wire mux_344_nl;
  wire or_1186_nl;
  wire or_1185_nl;
  wire or_1184_nl;
  wire or_1183_nl;
  wire mux_352_nl;
  wire mux_351_nl;
  wire mux_350_nl;
  wire mux_349_nl;
  wire mux_348_nl;
  wire mux_347_nl;
  wire or_1191_nl;
  wire or_1190_nl;
  wire or_1189_nl;
  wire or_1188_nl;
  wire or_1187_nl;
  wire mux_354_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_595_nl;
  wire or_1200_nl;
  wire mux_356_nl;
  wire or_1199_nl;
  wire or_1197_nl;
  wire mux_355_nl;
  wire or_1194_nl;
  wire mux_360_nl;
  wire mux_359_nl;
  wire mux_358_nl;
  wire nor_407_nl;
  wire nor_408_nl;
  wire or_1209_nl;
  wire mux_362_nl;
  wire or_1208_nl;
  wire or_1207_nl;
  wire mux_361_nl;
  wire or_1212_nl;
  wire or_1210_nl;
  wire mux_367_nl;
  wire nand_3_nl;
  wire or_1204_nl;
  wire mux_369_nl;
  wire mux_368_nl;
  wire or_1216_nl;
  wire or_1214_nl;
  wire mux_372_nl;
  wire mux_371_nl;
  wire or_1228_nl;
  wire or_1222_nl;
  wire or_1234_nl;
  wire or_1231_nl;
  wire mux_379_nl;
  wire mux_378_nl;
  wire mux_377_nl;
  wire or_1240_nl;
  wire or_1238_nl;
  wire mux_376_nl;
  wire or_1237_nl;
  wire or_1235_nl;
  wire mux_387_nl;
  wire mux_386_nl;
  wire mux_385_nl;
  wire mux_384_nl;
  wire nor_417_nl;
  wire nor_418_nl;
  wire nor_419_nl;
  wire nor_420_nl;
  wire mux_383_nl;
  wire mux_382_nl;
  wire mux_381_nl;
  wire nor_421_nl;
  wire nor_422_nl;
  wire nor_423_nl;
  wire nor_424_nl;
  wire mux_390_nl;
  wire mux_389_nl;
  wire or_1252_nl;
  wire or_1250_nl;
  wire mux_393_nl;
  wire mux_392_nl;
  wire or_1264_nl;
  wire or_1258_nl;
  wire or_1270_nl;
  wire or_1267_nl;
  wire mux_400_nl;
  wire mux_399_nl;
  wire mux_398_nl;
  wire or_1276_nl;
  wire or_1274_nl;
  wire mux_397_nl;
  wire or_1273_nl;
  wire or_1271_nl;
  wire mux_408_nl;
  wire mux_407_nl;
  wire mux_406_nl;
  wire mux_405_nl;
  wire nor_425_nl;
  wire nor_426_nl;
  wire nor_427_nl;
  wire nor_428_nl;
  wire mux_404_nl;
  wire mux_403_nl;
  wire mux_402_nl;
  wire nor_429_nl;
  wire nor_430_nl;
  wire nor_431_nl;
  wire nor_432_nl;
  wire mux_411_nl;
  wire mux_410_nl;
  wire or_1288_nl;
  wire or_1286_nl;
  wire mux_414_nl;
  wire mux_413_nl;
  wire or_1300_nl;
  wire or_1294_nl;
  wire or_1306_nl;
  wire or_1303_nl;
  wire mux_421_nl;
  wire mux_420_nl;
  wire mux_419_nl;
  wire or_1312_nl;
  wire or_1310_nl;
  wire mux_418_nl;
  wire or_1309_nl;
  wire or_1307_nl;
  wire mux_429_nl;
  wire mux_428_nl;
  wire mux_427_nl;
  wire mux_426_nl;
  wire nor_433_nl;
  wire nor_434_nl;
  wire nor_435_nl;
  wire nor_436_nl;
  wire mux_425_nl;
  wire mux_424_nl;
  wire mux_423_nl;
  wire nor_437_nl;
  wire nor_438_nl;
  wire nor_439_nl;
  wire nor_440_nl;
  wire mux_432_nl;
  wire mux_431_nl;
  wire or_1324_nl;
  wire or_1322_nl;
  wire mux_434_nl;
  wire or_1325_nl;
  wire mux_435_nl;
  wire or_1331_nl;
  wire mux_437_nl;
  wire mux_436_nl;
  wire or_1336_nl;
  wire or_1330_nl;
  wire or_1342_nl;
  wire or_1339_nl;
  wire mux_444_nl;
  wire mux_443_nl;
  wire mux_442_nl;
  wire or_1348_nl;
  wire or_1346_nl;
  wire mux_441_nl;
  wire or_1345_nl;
  wire or_1343_nl;
  wire mux_454_nl;
  wire mux_453_nl;
  wire mux_452_nl;
  wire mux_451_nl;
  wire nor_441_nl;
  wire nor_442_nl;
  wire mux_450_nl;
  wire nor_443_nl;
  wire nor_444_nl;
  wire mux_449_nl;
  wire nor_445_nl;
  wire nor_446_nl;
  wire mux_448_nl;
  wire mux_447_nl;
  wire nor_447_nl;
  wire nor_448_nl;
  wire mux_446_nl;
  wire nor_449_nl;
  wire nor_450_nl;
  wire mux_457_nl;
  wire mux_456_nl;
  wire or_1366_nl;
  wire or_1364_nl;
  wire while_mux_1254_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_626_nl;
  wire while_mux_1255_nl;
  wire Arbiter_8U_Roundrobin_pick_1_mux_625_nl;
  wire mux_460_nl;
  wire mux_459_nl;
  wire or_1376_nl;
  wire or_1371_nl;
  wire or_1384_nl;
  wire or_1380_nl;
  wire mux_468_nl;
  wire mux_467_nl;
  wire mux_466_nl;
  wire mux_465_nl;
  wire or_1397_nl;
  wire or_1386_nl;
  wire mux_464_nl;
  wire or_1398_nl;
  wire or_1385_nl;
  wire mux_469_nl;
  wire and_521_nl;
  wire weight_port_read_out_data_mux_8_nl;
  wire[6:0] weight_port_read_out_data_mux_22_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_5_nl;
  wire weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_5_nl;
  wire weight_mem_banks_write_if_for_if_and_35_nl;
  wire weight_mem_banks_write_if_for_if_and_36_nl;
  wire weight_mem_banks_write_if_for_if_and_37_nl;
  wire weight_mem_banks_write_if_for_if_and_38_nl;
  wire weight_mem_banks_write_if_for_if_and_39_nl;
  wire weight_mem_banks_write_if_for_if_and_40_nl;
  wire weight_mem_banks_write_if_for_if_and_41_nl;
  wire weight_mem_banks_write_if_for_if_mux_7_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_nl;
  wire mux_256_nl;
  wire nor_463_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_4_nl;
  wire weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_4_nl;
  wire weight_mem_banks_write_if_for_if_and_28_nl;
  wire weight_mem_banks_write_if_for_if_and_29_nl;
  wire weight_mem_banks_write_if_for_if_and_30_nl;
  wire weight_mem_banks_write_if_for_if_and_31_nl;
  wire weight_mem_banks_write_if_for_if_and_32_nl;
  wire weight_mem_banks_write_if_for_if_and_33_nl;
  wire weight_mem_banks_write_if_for_if_and_34_nl;
  wire weight_mem_banks_write_if_for_if_mux_6_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_1_nl;
  wire mux_255_nl;
  wire nor_462_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_3_nl;
  wire weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_3_nl;
  wire weight_mem_banks_write_if_for_if_and_21_nl;
  wire weight_mem_banks_write_if_for_if_and_22_nl;
  wire weight_mem_banks_write_if_for_if_and_23_nl;
  wire weight_mem_banks_write_if_for_if_and_24_nl;
  wire weight_mem_banks_write_if_for_if_and_25_nl;
  wire weight_mem_banks_write_if_for_if_and_26_nl;
  wire weight_mem_banks_write_if_for_if_and_27_nl;
  wire weight_mem_banks_write_if_for_if_mux_5_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_2_nl;
  wire mux_254_nl;
  wire nor_461_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_2_nl;
  wire weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_2_nl;
  wire weight_mem_banks_write_if_for_if_and_14_nl;
  wire weight_mem_banks_write_if_for_if_and_15_nl;
  wire weight_mem_banks_write_if_for_if_and_16_nl;
  wire weight_mem_banks_write_if_for_if_and_17_nl;
  wire weight_mem_banks_write_if_for_if_and_18_nl;
  wire weight_mem_banks_write_if_for_if_and_19_nl;
  wire weight_mem_banks_write_if_for_if_and_20_nl;
  wire weight_mem_banks_write_if_for_if_mux_4_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_3_nl;
  wire mux_253_nl;
  wire nor_460_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_1_nl;
  wire weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_1_nl;
  wire weight_mem_banks_write_if_for_if_and_7_nl;
  wire weight_mem_banks_write_if_for_if_and_8_nl;
  wire weight_mem_banks_write_if_for_if_and_9_nl;
  wire weight_mem_banks_write_if_for_if_and_10_nl;
  wire weight_mem_banks_write_if_for_if_and_11_nl;
  wire weight_mem_banks_write_if_for_if_and_12_nl;
  wire weight_mem_banks_write_if_for_if_and_13_nl;
  wire weight_mem_banks_write_if_for_if_mux_3_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_4_nl;
  wire mux_252_nl;
  wire nor_459_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_nl;
  wire weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_nl;
  wire weight_mem_banks_write_if_for_if_and_nl;
  wire weight_mem_banks_write_if_for_if_and_1_nl;
  wire weight_mem_banks_write_if_for_if_and_2_nl;
  wire weight_mem_banks_write_if_for_if_and_3_nl;
  wire weight_mem_banks_write_if_for_if_and_4_nl;
  wire weight_mem_banks_write_if_for_if_and_5_nl;
  wire weight_mem_banks_write_if_for_if_and_6_nl;
  wire weight_mem_banks_write_if_for_if_mux_2_nl;
  wire weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_5_nl;
  wire mux_251_nl;
  wire nor_458_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_mux_1_nl;
  wire weight_mem_banks_write_if_for_if_mux_54_nl;
  wire mux_250_nl;
  wire nor_457_nl;
  wire[10:0] weight_mem_banks_write_if_for_if_mux_nl;
  wire weight_mem_banks_write_if_for_if_mux_53_nl;
  wire mux_249_nl;
  wire nor_456_nl;
  wire rva_out_reg_data_mux_20_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_21_nl;
  wire PECore_DecodeAxiRead_switch_lp_mux_23_nl;
  wire rva_out_reg_data_mux_21_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_22_nl;
  wire PECore_DecodeAxiRead_switch_lp_mux_24_nl;
  wire rva_out_reg_data_mux_22_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_23_nl;
  wire PECore_DecodeAxiRead_switch_lp_mux_25_nl;
  wire PECore_PushAxiRsp_if_else_mux_17_nl;
  wire rva_out_reg_data_mux_24_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_25_nl;
  wire PECore_DecodeAxiRead_switch_lp_mux_26_nl;
  wire PECore_PushAxiRsp_if_else_mux_18_nl;
  wire rva_out_reg_data_mux_23_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_24_nl;
  wire mux_1255_nl;
  wire mux_1254_nl;
  wire mux_1256_nl;
  wire and_2582_nl;
  wire mux_1259_nl;
  wire or_3662_nl;
  wire or_3660_nl;
  wire mux_1258_nl;
  wire mux_1257_nl;
  wire mux_1262_nl;
  wire and_2584_nl;
  wire mux_1267_nl;
  wire mux_1266_nl;
  wire mux_1265_nl;
  wire mux_1264_nl;
  wire mux_1263_nl;
  wire mux_1269_nl;
  wire or_3670_nl;
  wire mux_1283_nl;
  wire mux_1282_nl;
  wire mux_1281_nl;
  wire mux_1280_nl;
  wire mux_1279_nl;
  wire mux_1278_nl;
  wire mux_1277_nl;
  wire or_3684_nl;
  wire mux_1290_nl;
  wire mux_1297_nl;
  wire mux_175_nl;
  wire mux_174_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_16_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_14_nl;
  wire PECore_DecodeAxiRead_switch_lp_mux_20_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_11_nl;
  wire PECore_DecodeAxiRead_switch_lp_mux_21_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_28_nl;
  wire PECore_DecodeAxiRead_switch_lp_mux_28_nl;
  wire[4:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_29_nl;
  wire[4:0] PECore_DecodeAxiRead_switch_lp_mux_29_nl;
  wire[2:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_8_nl;
  wire[2:0] PECore_DecodeAxiRead_switch_lp_mux_22_nl;
  wire[2:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_30_nl;
  wire[2:0] PECore_DecodeAxiRead_switch_lp_mux_30_nl;
  wire PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_26_nl;
  wire[4:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_31_nl;
  wire[2:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_27_nl;
  wire[2:0] PECore_DecodeAxiRead_switch_lp_mux_27_nl;
  wire[2:0] PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_32_nl;
  wire[2:0] PECore_DecodeAxiRead_switch_lp_mux_31_nl;
  wire or_1480_nl;
  wire or_1481_nl;
  wire or_1482_nl;
  wire and_2590_nl;
  wire and_2591_nl;
  wire mux_1076_nl;
  wire and_2435_nl;
  wire nor_1421_nl;
  wire mux_914_nl;
  wire and_2337_nl;
  wire nor_1193_nl;
  wire mux_1226_nl;
  wire and_2547_nl;
  wire nor_1638_nl;
  wire mux_1072_nl;
  wire nor_1414_nl;
  wire nor_1415_nl;
  wire mux_1114_nl;
  wire nand_277_nl;
  wire or_3244_nl;
  wire mux_962_nl;
  wire nand_184_nl;
  wire or_2782_nl;
  wire mux_1116_nl;
  wire nand_278_nl;
  wire or_3250_nl;
  wire mux_1234_nl;
  wire and_2560_nl;
  wire and_2561_nl;
  wire mux_1000_nl;
  wire nor_1315_nl;
  wire nor_1316_nl;
  wire mux_1092_nl;
  wire nand_259_nl;
  wire or_3180_nl;
  wire mux_1220_nl;
  wire nand_347_nl;
  wire or_3555_nl;
  wire mux_1196_nl;
  wire and_2521_nl;
  wire nor_1593_nl;
  wire mux_1018_nl;
  wire or_2952_nl;
  wire or_2948_nl;
  wire mux_1090_nl;
  wire nand_258_nl;
  wire or_3174_nl;
  wire mux_764_nl;
  wire or_2162_nl;
  wire or_2158_nl;
  wire mux_900_nl;
  wire nand_147_nl;
  wire or_2590_nl;
  wire mux_884_nl;
  wire nor_1153_nl;
  wire nor_1154_nl;
  wire mux_906_nl;
  wire nor_1181_nl;
  wire nor_1182_nl;
  wire mux_936_nl;
  wire nor_1223_nl;
  wire nor_1224_nl;
  wire mux_1118_nl;
  wire nand_279_nl;
  wire or_3255_nl;
  wire mux_1066_nl;
  wire nor_1406_nl;
  wire nor_1407_nl;
  wire mux_1152_nl;
  wire nand_299_nl;
  wire or_3360_nl;
  wire mux_928_nl;
  wire nand_164_nl;
  wire or_2678_nl;
  wire mux_850_nl;
  wire and_2306_nl;
  wire nor_1105_nl;
  wire mux_818_nl;
  wire nor_1062_nl;
  wire nor_1063_nl;
  wire mux_1126_nl;
  wire and_2469_nl;
  wire nor_1493_nl;
  wire mux_1160_nl;
  wire nor_1539_nl;
  wire nor_1540_nl;
  wire mux_1182_nl;
  wire nand_321_nl;
  wire or_3446_nl;
  wire mux_1020_nl;
  wire or_2959_nl;
  wire or_2955_nl;
  wire mux_1134_nl;
  wire and_2475_nl;
  wire nor_1505_nl;
  wire mux_1156_nl;
  wire nand_301_nl;
  wire or_3371_nl;
  wire mux_1190_nl;
  wire and_2515_nl;
  wire nor_1585_nl;
  wire mux_1150_nl;
  wire nand_298_nl;
  wire or_3354_nl;
  wire mux_844_nl;
  wire nor_1096_nl;
  wire nor_1097_nl;
  wire mux_886_nl;
  wire nand_144_nl;
  wire or_2544_nl;
  wire mux_964_nl;
  wire nand_185_nl;
  wire or_2788_nl;
  wire mux_746_nl;
  wire nor_967_nl;
  wire nor_968_nl;
  wire mux_940_nl;
  wire nor_1229_nl;
  wire nor_1230_nl;
  wire mux_872_nl;
  wire nor_1135_nl;
  wire nor_1136_nl;
  wire mux_944_nl;
  wire nor_1234_nl;
  wire nor_1235_nl;
  wire mux_846_nl;
  wire and_2303_nl;
  wire nor_1100_nl;
  wire mux_1106_nl;
  wire and_2453_nl;
  wire nor_1463_nl;
  wire mux_960_nl;
  wire nand_183_nl;
  wire or_2777_nl;
  wire mux_862_nl;
  wire nand_131_nl;
  wire or_2471_nl;
  wire mux_908_nl;
  wire nor_1184_nl;
  wire nor_1185_nl;
  wire mux_1170_nl;
  wire and_2499_nl;
  wire nor_1555_nl;
  wire mux_808_nl;
  wire nor_1047_nl;
  wire nor_1048_nl;
  wire mux_788_nl;
  wire nor_1022_nl;
  wire nor_1023_nl;
  wire mux_1088_nl;
  wire nand_257_nl;
  wire or_3169_nl;
  wire mux_1024_nl;
  wire or_2974_nl;
  wire or_2967_nl;
  wire mux_970_nl;
  wire and_2367_nl;
  wire nor_1271_nl;
  wire mux_1214_nl;
  wire nand_344_nl;
  wire or_3538_nl;
  wire mux_1218_nl;
  wire nand_346_nl;
  wire nand_486_nl;
  wire mux_1044_nl;
  wire and_2417_nl;
  wire nor_1376_nl;
  wire mux_1228_nl;
  wire and_2551_nl;
  wire nor_1641_nl;
  wire mux_1232_nl;
  wire and_2556_nl;
  wire and_2557_nl;
  wire mux_1004_nl;
  wire nor_1321_nl;
  wire nor_1322_nl;
  wire mux_930_nl;
  wire nand_165_nl;
  wire or_2683_nl;
  wire mux_1194_nl;
  wire and_2518_nl;
  wire nor_1590_nl;
  wire mux_1078_nl;
  wire nand_253_nl;
  wire or_3137_nl;
  wire mux_794_nl;
  wire or_2257_nl;
  wire or_2253_nl;
  wire mux_990_nl;
  wire nand_205_nl;
  wire or_2863_nl;
  wire mux_832_nl;
  wire or_2381_nl;
  wire or_2374_nl;
  wire mux_920_nl;
  wire or_2659_nl;
  wire or_2652_nl;
  wire mux_892_nl;
  wire or_2567_nl;
  wire or_2563_nl;
  wire mux_1068_nl;
  wire nor_1409_nl;
  wire nor_1410_nl;
  wire mux_864_nl;
  wire nand_132_nl;
  wire or_2477_nl;
  wire mux_768_nl;
  wire or_2175_nl;
  wire or_2171_nl;
  wire mux_866_nl;
  wire nand_133_nl;
  wire or_2482_nl;
  wire mux_806_nl;
  wire and_2284_nl;
  wire nor_1045_nl;
  wire mux_754_nl;
  wire nor_979_nl;
  wire nor_980_nl;
  wire mux_1162_nl;
  wire and_2490_nl;
  wire nor_1543_nl;
  wire mux_804_nl;
  wire nand_102_nl;
  wire or_2287_nl;
  wire mux_978_nl;
  wire and_2376_nl;
  wire nor_1283_nl;
  wire mux_1202_nl;
  wire and_2527_nl;
  wire nor_1602_nl;
  wire mux_1242_nl;
  wire nand_366_nl;
  wire nand_502_nl;
  wire mux_1176_nl;
  wire nand_318_nl;
  wire or_3430_nl;
  wire mux_1248_nl;
  wire nand_369_nl;
  wire nand_507_nl;
  wire mux_1166_nl;
  wire and_2495_nl;
  wire nor_1549_nl;
  wire mux_1006_nl;
  wire nor_1324_nl;
  wire nor_1325_nl;
  wire mux_828_nl;
  wire or_2366_nl;
  wire or_2362_nl;
  wire mux_1062_nl;
  wire and_2423_nl;
  wire nor_1401_nl;
  wire mux_826_nl;
  wire or_2359_nl;
  wire or_2355_nl;
  wire mux_912_nl;
  wire nor_1189_nl;
  wire nor_1190_nl;
  wire mux_750_nl;
  wire nor_973_nl;
  wire nor_974_nl;
  wire mux_774_nl;
  wire and_2271_nl;
  wire nor_1002_nl;
  wire mux_792_nl;
  wire or_2251_nl;
  wire or_2247_nl;
  wire mux_834_nl;
  wire nand_114_nl;
  wire or_2383_nl;
  wire mux_842_nl;
  wire nor_1093_nl;
  wire nor_1094_nl;
  wire mux_822_nl;
  wire nand_112_nl;
  wire or_2343_nl;
  wire mux_976_nl;
  wire and_2374_nl;
  wire nor_1280_nl;
  wire mux_1010_nl;
  wire nor_1330_nl;
  wire nor_1331_nl;
  wire mux_1052_nl;
  wire nand_236_nl;
  wire or_3059_nl;
  wire mux_1250_nl;
  wire nand_370_nl;
  wire nand_508_nl;
  wire mux_776_nl;
  wire nor_1004_nl;
  wire nor_1005_nl;
  wire mux_1158_nl;
  wire and_2487_nl;
  wire nor_1538_nl;
  wire mux_1112_nl;
  wire nand_276_nl;
  wire or_3239_nl;
  wire mux_1180_nl;
  wire nand_320_nl;
  wire or_3441_nl;
  wire mux_992_nl;
  wire nand_206_nl;
  wire nand_441_nl;
  wire mux_878_nl;
  wire nor_1144_nl;
  wire nor_1145_nl;
  wire mux_790_nl;
  wire nand_99_nl;
  wire or_2241_nl;
  wire mux_766_nl;
  wire or_2168_nl;
  wire or_2164_nl;
  wire mux_860_nl;
  wire nand_130_nl;
  wire or_2466_nl;
  wire mux_1140_nl;
  wire and_2481_nl;
  wire nor_1513_nl;
  wire mux_1054_nl;
  wire nand_237_nl;
  wire or_3064_nl;
  wire mux_896_nl;
  wire or_2582_nl;
  wire or_2575_nl;
  wire mux_1174_nl;
  wire nand_317_nl;
  wire or_3424_nl;
  wire mux_810_nl;
  wire nor_1050_nl;
  wire nor_1051_nl;
  wire mux_1244_nl;
  wire nand_367_nl;
  wire or_3621_nl;
  wire mux_1198_nl;
  wire and_2523_nl;
  wire nor_1596_nl;
  wire mux_898_nl;
  wire nand_146_nl;
  wire or_2584_nl;
  wire mux_876_nl;
  wire nor_1141_nl;
  wire nor_1142_nl;
  wire mux_780_nl;
  wire nor_1010_nl;
  wire nor_1011_nl;
  wire mux_796_nl;
  wire or_2264_nl;
  wire or_2260_nl;
  wire mux_904_nl;
  wire nor_1178_nl;
  wire nor_1179_nl;
  wire mux_1070_nl;
  wire and_2429_nl;
  wire nor_1413_nl;
  wire mux_1108_nl;
  wire and_2457_nl;
  wire nor_1466_nl;
  wire mux_1100_nl;
  wire and_2447_nl;
  wire nor_1454_nl;
  wire mux_1120_nl;
  wire nand_280_nl;
  wire nand_462_nl;
  wire mux_1168_nl;
  wire and_2497_nl;
  wire nor_1552_nl;
  wire mux_1210_nl;
  wire nand_342_nl;
  wire or_3527_nl;
  wire mux_1238_nl;
  wire nand_364_nl;
  wire or_3604_nl;
  wire mux_1240_nl;
  wire nand_365_nl;
  wire nand_501_nl;
  wire mux_966_nl;
  wire and_2364_nl;
  wire nor_1266_nl;
  wire mux_1206_nl;
  wire nand_340_nl;
  wire or_3516_nl;
  wire mux_1104_nl;
  wire and_2451_nl;
  wire nor_1460_nl;
  wire mux_778_nl;
  wire nor_1007_nl;
  wire nor_1008_nl;
  wire mux_1178_nl;
  wire nand_319_nl;
  wire or_3435_nl;
  wire mux_902_nl;
  wire and_2328_nl;
  wire nor_1176_nl;
  wire mux_984_nl;
  wire nand_202_nl;
  wire or_2847_nl;
  wire mux_772_nl;
  wire or_2188_nl;
  wire or_2184_nl;
  wire mux_926_nl;
  wire nand_163_nl;
  wire or_2672_nl;
  wire mux_1046_nl;
  wire nand_234_nl;
  wire or_3038_nl;
  wire mux_1148_nl;
  wire nand_297_nl;
  wire or_3349_nl;
  wire mux_742_nl;
  wire nor_961_nl;
  wire mux_741_nl;
  wire or_2090_nl;
  wire or_2089_nl;
  wire nor_962_nl;
  wire mux_830_nl;
  wire nand_113_nl;
  wire or_2368_nl;
  wire mux_1216_nl;
  wire nand_345_nl;
  wire nand_485_nl;
  wire mux_952_nl;
  wire or_2758_nl;
  wire or_2751_nl;
  wire mux_910_nl;
  wire and_2334_nl;
  wire nor_1188_nl;
  wire mux_1128_nl;
  wire nor_1495_nl;
  wire nor_1496_nl;
  wire mux_1192_nl;
  wire nor_1586_nl;
  wire nor_1587_nl;
  wire mux_784_nl;
  wire nor_1016_nl;
  wire nor_1017_nl;
  wire mux_1028_nl;
  wire nand_221_nl;
  wire or_2982_nl;
  wire mux_856_nl;
  wire or_2458_nl;
  wire or_2451_nl;
  wire mux_1050_nl;
  wire nand_235_nl;
  wire or_3053_nl;
  wire mux_868_nl;
  wire nand_134_nl;
  wire or_2488_nl;
  wire mux_954_nl;
  wire nand_180_nl;
  wire or_2760_nl;
  wire mux_916_nl;
  wire and_2340_nl;
  wire nor_1196_nl;
  wire mux_1096_nl;
  wire nor_1447_nl;
  wire nor_1448_nl;
  wire mux_1144_nl;
  wire or_3341_nl;
  wire or_3334_nl;
  wire mux_986_nl;
  wire nand_203_nl;
  wire or_2852_nl;
  wire mux_968_nl;
  wire nor_1267_nl;
  wire nor_1268_nl;
  wire mux_918_nl;
  wire nand_160_nl;
  wire or_2646_nl;
  wire mux_890_nl;
  wire or_2560_nl;
  wire or_2556_nl;
  wire mux_922_nl;
  wire nand_161_nl;
  wire or_2661_nl;
  wire mux_824_nl;
  wire or_2353_nl;
  wire or_2349_nl;
  wire mux_756_nl;
  wire nor_982_nl;
  wire nor_983_nl;
  wire mux_1212_nl;
  wire nand_343_nl;
  wire or_3533_nl;
  wire mux_994_nl;
  wire nand_207_nl;
  wire nand_442_nl;
  wire mux_1034_nl;
  wire nor_1361_nl;
  wire nor_1362_nl;
  wire mux_1200_nl;
  wire and_2525_nl;
  wire nor_1599_nl;
  wire mux_1188_nl;
  wire nand_324_nl;
  wire or_3463_nl;
  wire mux_1064_nl;
  wire nor_1403_nl;
  wire nor_1404_nl;
  wire mux_1154_nl;
  wire nand_300_nl;
  wire or_3365_nl;
  wire mux_1002_nl;
  wire nor_1318_nl;
  wire nor_1319_nl;
  wire mux_1132_nl;
  wire nor_1501_nl;
  wire nor_1502_nl;
  wire mux_948_nl;
  wire and_2358_nl;
  wire nor_1241_nl;
  wire mux_942_nl;
  wire and_2352_nl;
  wire nor_1233_nl;
  wire mux_1056_nl;
  wire nand_238_nl;
  wire or_3070_nl;
  wire mux_996_nl;
  wire nand_208_nl;
  wire or_2880_nl;
  wire mux_840_nl;
  wire nor_1090_nl;
  wire nor_1091_nl;
  wire mux_836_nl;
  wire nand_115_nl;
  wire or_2389_nl;
  wire mux_1222_nl;
  wire and_2543_nl;
  wire nor_1632_nl;
  wire mux_1186_nl;
  wire nand_323_nl;
  wire nand_476_nl;
  wire mux_982_nl;
  wire nand_201_nl;
  wire or_2841_nl;
  wire mux_874_nl;
  wire nor_1138_nl;
  wire nor_1139_nl;
  wire mux_812_nl;
  wire nor_1053_nl;
  wire nor_1054_nl;
  wire mux_1008_nl;
  wire nor_1327_nl;
  wire nor_1328_nl;
  wire mux_1086_nl;
  wire nand_256_nl;
  wire or_3163_nl;
  wire mux_880_nl;
  wire nor_1147_nl;
  wire nor_1148_nl;
  wire mux_958_nl;
  wire nand_182_nl;
  wire or_2771_nl;
  wire mux_770_nl;
  wire or_2181_nl;
  wire or_2177_nl;
  wire mux_1060_nl;
  wire nand_240_nl;
  wire or_3081_nl;
  wire mux_894_nl;
  wire nand_145_nl;
  wire or_2569_nl;
  wire mux_1224_nl;
  wire and_2545_nl;
  wire nor_1635_nl;
  wire mux_1084_nl;
  wire nand_255_nl;
  wire or_3158_nl;
  wire mux_1142_nl;
  wire nand_295_nl;
  wire or_3328_nl;
  wire mux_938_nl;
  wire nor_1226_nl;
  wire nor_1227_nl;
  wire mux_1208_nl;
  wire nand_341_nl;
  wire or_3522_nl;
  wire mux_1038_nl;
  wire and_2411_nl;
  wire nor_1368_nl;
  wire mux_950_nl;
  wire nand_179_nl;
  wire or_2745_nl;
  wire mux_852_nl;
  wire and_2309_nl;
  wire nor_1108_nl;
  wire mux_988_nl;
  wire nand_204_nl;
  wire or_2858_nl;
  wire mux_980_nl;
  wire and_2380_nl;
  wire nor_1286_nl;
  wire mux_1012_nl;
  wire nor_1333_nl;
  wire nor_1334_nl;
  wire mux_974_nl;
  wire and_2372_nl;
  wire nor_1277_nl;
  wire mux_998_nl;
  wire and_2392_nl;
  wire nor_1313_nl;
  wire mux_1130_nl;
  wire nor_1498_nl;
  wire nor_1499_nl;
  wire mux_802_nl;
  wire nand_101_nl;
  wire or_2281_nl;
  wire mux_1014_nl;
  wire nand_218_nl;
  wire or_2936_nl;
  wire mux_1253_nl;
  wire and_2581_nl;
  wire nand_511_nl;
  wire mux_1184_nl;
  wire nand_322_nl;
  wire nand_475_nl;
  wire mux_1230_nl;
  wire and_2553_nl;
  wire nor_1644_nl;
  wire mux_798_nl;
  wire nand_100_nl;
  wire or_2266_nl;
  wire mux_1204_nl;
  wire and_2531_nl;
  wire nor_1605_nl;
  wire mux_1102_nl;
  wire and_2449_nl;
  wire nor_1457_nl;
  wire mux_1032_nl;
  wire nor_1358_nl;
  wire nor_1359_nl;
  wire mux_1042_nl;
  wire and_2414_nl;
  wire nor_1373_nl;
  wire mux_934_nl;
  wire and_2346_nl;
  wire nor_1221_nl;
  wire mux_1022_nl;
  wire nand_219_nl;
  wire or_2961_nl;
  wire mux_758_nl;
  wire or_2142_nl;
  wire or_2138_nl;
  wire mux_924_nl;
  wire nand_162_nl;
  wire or_2667_nl;
  wire mux_1146_nl;
  wire nand_296_nl;
  wire or_3343_nl;
  wire mux_782_nl;
  wire nor_1013_nl;
  wire nor_1014_nl;
  wire mux_1080_nl;
  wire or_3150_nl;
  wire or_3143_nl;
  wire mux_1094_nl;
  wire and_2441_nl;
  wire nor_1446_nl;
  wire mux_1058_nl;
  wire nand_239_nl;
  wire or_3075_nl;
  wire mux_1040_nl;
  wire nor_1369_nl;
  wire nor_1370_nl;
  wire mux_1036_nl;
  wire nor_1364_nl;
  wire nor_1365_nl;
  wire mux_848_nl;
  wire nor_1101_nl;
  wire nor_1102_nl;
  wire mux_800_nl;
  wire or_2279_nl;
  wire or_2272_nl;
  wire mux_1048_nl;
  wire or_3051_nl;
  wire or_3044_nl;
  wire mux_1246_nl;
  wire nand_368_nl;
  wire nand_505_nl;
  wire mux_748_nl;
  wire nor_970_nl;
  wire nor_971_nl;
  wire mux_946_nl;
  wire and_2355_nl;
  wire nor_1238_nl;
  wire mux_956_nl;
  wire nand_181_nl;
  wire or_2766_nl;
  wire mux_760_nl;
  wire or_2149_nl;
  wire or_2145_nl;
  wire mux_1016_nl;
  wire or_2946_nl;
  wire or_2942_nl;
  wire mux_972_nl;
  wire and_2370_nl;
  wire nor_1274_nl;
  wire mux_1082_nl;
  wire nand_254_nl;
  wire or_3152_nl;
  wire mux_1164_nl;
  wire and_2493_nl;
  wire nor_1546_nl;
  wire mux_762_nl;
  wire or_2155_nl;
  wire or_2151_nl;
  wire mux_1136_nl;
  wire nor_1506_nl;
  wire nor_1507_nl;
  wire mux_870_nl;
  wire and_2315_nl;
  wire nor_1133_nl;
  wire mux_1074_nl;
  wire and_2432_nl;
  wire nor_1418_nl;
  wire mux_1124_nl;
  wire nand_282_nl;
  wire or_3272_nl;
  wire mux_1138_nl;
  wire and_2478_nl;
  wire nor_1510_nl;
  wire mux_1122_nl;
  wire nand_281_nl;
  wire nand_463_nl;
  wire mux_752_nl;
  wire nor_976_nl;
  wire nor_977_nl;
  wire mux_1110_nl;
  wire nand_275_nl;
  wire or_3233_nl;
  wire mux_1172_nl;
  wire and_2503_nl;
  wire nor_1558_nl;
  wire mux_816_nl;
  wire nor_1059_nl;
  wire nor_1060_nl;
  wire mux_1236_nl;
  wire and_2565_nl;
  wire nor_1651_nl;
  wire mux_814_nl;
  wire nor_1056_nl;
  wire nor_1057_nl;
  wire mux_1026_nl;
  wire nand_220_nl;
  wire or_2976_nl;
  wire mux_1098_nl;
  wire and_2444_nl;
  wire nor_1451_nl;
  wire mux_888_nl;
  wire or_2554_nl;
  wire or_2550_nl;
  wire mux_1030_nl;
  wire and_2405_nl;
  wire nor_1356_nl;
  wire mux_786_nl;
  wire nor_1019_nl;
  wire nor_1020_nl;
  wire mux_838_nl;
  wire and_2297_nl;
  wire nor_1088_nl;
  wire mux_854_nl;
  wire nand_128_nl;
  wire or_2445_nl;
  wire mux_820_nl;
  wire nor_1065_nl;
  wire nor_1066_nl;
  wire mux_858_nl;
  wire nand_129_nl;
  wire or_2460_nl;
  wire mux_744_nl;
  wire nor_964_nl;
  wire nor_965_nl;
  wire mux_932_nl;
  wire nand_166_nl;
  wire or_2689_nl;
  wire mux_882_nl;
  wire nor_1150_nl;
  wire nor_1151_nl;
  wire mux_530_nl;
  wire or_1590_nl;
  wire mux_529_nl;
  wire nor_927_nl;
  wire or_1587_nl;

  // Interconnect Declarations for Component Instantiations 
  wire  nl_weight_mem_read_arbxbar_xbar_for_1_lshift_rg_a;
  assign nl_weight_mem_read_arbxbar_xbar_for_1_lshift_rg_a = PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2
      & (~ reg_rva_in_reg_rw_sva_2_cse);
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_for_1_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_for_1_lshift_rg_s = weight_read_addrs_0_3_0_lpi_1_dfm_1_2[2:0];
  wire  nl_weight_mem_write_arbxbar_xbar_for_lshift_rg_a;
  assign nl_weight_mem_write_arbxbar_xbar_for_lshift_rg_a = PECore_DecodeAxiWrite_switch_lp_equal_tmp_1_2
      & reg_rva_in_reg_rw_sva_2_cse;
  wire [2:0] nl_weight_mem_write_arbxbar_xbar_for_lshift_rg_s;
  assign nl_weight_mem_write_arbxbar_xbar_for_lshift_rg_s = weight_write_addrs_lpi_1_dfm_1_2[2:0];
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_7_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_7_lshift_rg_s = {(weight_read_addrs_6_14_1_lpi_1_dfm_1_1[1:0])
      , (weight_read_addrs_0_3_0_lpi_1_dfm_4[0])};
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_1_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_1_lshift_rg_s = weight_read_addrs_0_3_0_lpi_1_dfm_4[2:0];
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_8_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_8_lshift_rg_s = weight_read_addrs_7_lpi_1_dfm_1_1[2:0];
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_3_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_3_lshift_rg_s = {(weight_read_addrs_2_14_1_lpi_1_dfm_1_1[1:0])
      , (weight_read_addrs_0_3_0_lpi_1_dfm_4[0])};
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_5_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_5_lshift_rg_s = {(weight_read_addrs_4_14_2_lpi_1_dfm_1_1[0])
      , (weight_read_addrs_0_3_0_lpi_1_dfm_4[1:0])};
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_4_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_4_lshift_rg_s = weight_read_addrs_3_lpi_1_dfm_1_1[2:0];
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_6_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_6_lshift_rg_s = weight_read_addrs_5_lpi_1_dfm_1_1[2:0];
  wire [2:0] nl_weight_mem_read_arbxbar_xbar_1_for_2_lshift_rg_s;
  assign nl_weight_mem_read_arbxbar_xbar_1_for_2_lshift_rg_s = weight_read_addrs_1_lpi_1_dfm_1_1[2:0];
  wire [255:0] nl_PECore_PECoreRun_act_port_Push_mioi_inst_act_port_Push_mioi_m_data_rsc_dat_PECoreRun;
  assign nl_PECore_PECoreRun_act_port_Push_mioi_inst_act_port_Push_mioi_m_data_rsc_dat_PECoreRun
      = signext_256_244({act_port_reg_data_243_224_sva_dfm_1_1 , ({{12{act_port_reg_data_211_192_sva_dfm_1_1[19]}},
      act_port_reg_data_211_192_sva_dfm_1_1}) , ({{12{act_port_reg_data_179_160_sva_dfm_1_1[19]}},
      act_port_reg_data_179_160_sva_dfm_1_1}) , ({{12{act_port_reg_data_147_128_sva_dfm_1_1[19]}},
      act_port_reg_data_147_128_sva_dfm_1_1}) , ({{12{act_port_reg_data_115_96_sva_dfm_1_1[19]}},
      act_port_reg_data_115_96_sva_dfm_1_1}) , ({{12{act_port_reg_data_83_64_sva_dfm_1_1[19]}},
      act_port_reg_data_83_64_sva_dfm_1_1}) , ({{12{act_port_reg_data_51_32_sva_dfm_1_1[19]}},
      act_port_reg_data_51_32_sva_dfm_1_1}) , ({{12{act_port_reg_data_19_0_sva_dfm_1_1[19]}},
      act_port_reg_data_19_0_sva_dfm_1_1})});
  wire weight_port_read_out_data_mux_4_nl;
  wire weight_port_read_out_data_mux_25_nl;
  wire weight_port_read_out_data_mux_2_nl;
  wire weight_port_read_out_data_mux_24_nl;
  wire weight_port_read_out_data_mux_nl;
  wire weight_port_read_out_data_mux_23_nl;
  wire [63:0] nl_PECore_PECoreRun_rva_out_Push_mioi_inst_rva_out_Push_mioi_m_data_rsc_dat_PECoreRun;
  assign weight_port_read_out_data_mux_25_nl = MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_16_itm,
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_0_itm_1, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7);
  assign weight_port_read_out_data_mux_4_nl = MUX_s_1_2_2(weight_port_read_out_data_slc_weight_port_read_out_data_0_2_0_itm_1,
      weight_port_read_out_data_mux_25_nl, fsm_output);
  assign weight_port_read_out_data_mux_24_nl = MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_15_itm,
      weight_port_read_out_data_slc_weight_port_read_out_data_0_1_0_itm_1, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7);
  assign weight_port_read_out_data_mux_2_nl = MUX_s_1_2_2(weight_port_read_out_data_slc_weight_port_read_out_data_0_1_0_itm_1,
      weight_port_read_out_data_mux_24_nl, fsm_output);
  assign weight_port_read_out_data_mux_23_nl = MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_14_itm,
      weight_port_read_out_data_slc_weight_port_read_out_data_0_0_0_itm_1, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7);
  assign weight_port_read_out_data_mux_nl = MUX_s_1_2_2(weight_port_read_out_data_slc_weight_port_read_out_data_0_0_0_itm_1,
      weight_port_read_out_data_mux_23_nl, fsm_output);
  assign nl_PECore_PECoreRun_rva_out_Push_mioi_inst_rva_out_Push_mioi_m_data_rsc_dat_PECoreRun
      = {rva_out_reg_data_63_sva_dfm_4_4 , rva_out_reg_data_62_56_sva_dfm_4_4 , reg_rva_out_reg_data_55_48_sva_dfm_4_4_ftd
      , reg_rva_out_reg_data_55_48_sva_dfm_4_4_ftd_1 , rva_out_reg_data_47_sva_dfm_4_4
      , reg_rva_out_reg_data_46_40_sva_dfm_4_4_ftd , reg_rva_out_reg_data_46_40_sva_dfm_4_4_ftd_1
      , reg_rva_out_reg_data_39_36_sva_dfm_4_4_ftd , reg_rva_out_reg_data_39_36_sva_dfm_4_4_ftd_1
      , reg_rva_out_reg_data_39_36_sva_dfm_4_4_ftd_2 , rva_out_reg_data_35_32_sva_dfm_4_4
      , PECore_PushAxiRsp_if_mux1h_17 , PECore_PushAxiRsp_if_mux1h_16_5_3 , PECore_PushAxiRsp_if_mux1h_16_2_0
      , PECore_PushAxiRsp_if_mux1h_15 , PECore_PushAxiRsp_if_mux1h_14_6 , PECore_PushAxiRsp_if_mux1h_14_5
      , PECore_PushAxiRsp_if_mux1h_14_4_0 , weight_port_read_out_data_mux_4_nl ,
      PECore_PushAxiRsp_if_mux1h_12_6 , PECore_PushAxiRsp_if_mux1h_12_5_3 , PECore_PushAxiRsp_if_mux1h_12_2_0
      , weight_port_read_out_data_mux_2_nl , PECore_PushAxiRsp_if_mux1h_10_6 , PECore_PushAxiRsp_if_mux1h_10_5
      , PECore_PushAxiRsp_if_mux1h_10_4_0 , weight_port_read_out_data_mux_nl};
  PECore_mgc_muladd1 #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd8),
  .signd_c(32'sd0),
  .width_cst(32'sd1),
  .signd_cst(32'sd0),
  .width_d(32'sd0),
  .signd_d(32'sd1),
  .width_z(32'sd11),
  .add_axb(32'sd1),
  .add_c(32'sd1),
  .add_d(32'sd1),
  .use_const(32'sd1)) PEManager_15U_GetWeightAddr_else_acc_4_cmp (
      .a(pe_config_output_counter_sva),
      .b(pe_manager_num_input_sva),
      .c(pe_config_input_counter_sva),
      .cst(1'b0),
      .z(PEManager_15U_GetWeightAddr_else_acc_4_cmp_z),
      .d(2'b0)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_for_1_lshift_rg (
      .a(nl_weight_mem_read_arbxbar_xbar_for_1_lshift_rg_a),
      .s(nl_weight_mem_read_arbxbar_xbar_for_1_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_for_1_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_write_arbxbar_xbar_for_lshift_rg (
      .a(nl_weight_mem_write_arbxbar_xbar_for_lshift_rg_a),
      .s(nl_weight_mem_write_arbxbar_xbar_for_lshift_rg_s[2:0]),
      .z(weight_mem_write_arbxbar_xbar_for_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_7_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_7_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_1_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_1_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_8_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_8_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_3_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_3_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_5_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_5_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_4_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_4_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_6_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_6_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp)
    );
  PECore_mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) weight_mem_read_arbxbar_xbar_1_for_2_lshift_rg (
      .a(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2),
      .s(nl_weight_mem_read_arbxbar_xbar_1_for_2_lshift_rg_s[2:0]),
      .z(weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp)
    );
  PECore_PECore_PECoreRun_rva_in_PopNB_mioi PECore_PECoreRun_rva_in_PopNB_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_in_vld(rva_in_vld),
      .rva_in_rdy(rva_in_rdy),
      .rva_in_dat(rva_in_dat),
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .rva_in_PopNB_mioi_oswt(reg_rva_in_PopNB_mioi_iswt0_cse),
      .rva_in_PopNB_mioi_data_data_rsc_z_mxwt(rva_in_PopNB_mioi_data_data_rsc_z_mxwt),
      .rva_in_PopNB_mioi_data_addr_rsc_z_mxwt(rva_in_PopNB_mioi_data_addr_rsc_z_mxwt),
      .rva_in_PopNB_mioi_data_rw_rsc_z_mxwt(rva_in_PopNB_mioi_data_rw_rsc_z_mxwt),
      .rva_in_PopNB_mioi_return_rsc_z_mxwt(rva_in_PopNB_mioi_return_rsc_z_mxwt),
      .rva_in_PopNB_mioi_oswt_pff(fsm_output)
    );
  PECore_PECore_PECoreRun_input_port_PopNB_mioi PECore_PECoreRun_input_port_PopNB_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .input_port_vld(input_port_vld),
      .input_port_rdy(input_port_rdy),
      .input_port_dat(input_port_dat),
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .input_port_PopNB_mioi_oswt(reg_start_PopNB_mioi_iswt0_cse),
      .input_port_PopNB_mioi_data_data_data_rsc_z_mxwt(input_port_PopNB_mioi_data_data_data_rsc_z_mxwt),
      .input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt(input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt),
      .input_port_PopNB_mioi_return_rsc_z_mxwt(input_port_PopNB_mioi_return_rsc_z_mxwt),
      .input_port_PopNB_mioi_oswt_pff(and_518_rmff)
    );
  PECore_PECore_PECoreRun_act_port_Push_mioi PECore_PECoreRun_act_port_Push_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .act_port_vld(act_port_vld),
      .act_port_rdy(act_port_rdy),
      .act_port_dat(act_port_dat),
      .PECoreRun_wen(PECoreRun_wen),
      .act_port_Push_mioi_oswt(reg_act_port_Push_mioi_iswt0_cse),
      .act_port_Push_mioi_wen_comp(act_port_Push_mioi_wen_comp),
      .act_port_Push_mioi_m_data_rsc_dat_PECoreRun(nl_PECore_PECoreRun_act_port_Push_mioi_inst_act_port_Push_mioi_m_data_rsc_dat_PECoreRun[255:0]),
      .act_port_Push_mioi_oswt_pff(and_520_rmff)
    );
  PECore_PECore_PECoreRun_start_PopNB_mioi PECore_PECoreRun_start_PopNB_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .start_vld(start_vld),
      .start_rdy(start_rdy),
      .start_dat(start_dat),
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .start_PopNB_mioi_oswt(reg_start_PopNB_mioi_iswt0_cse),
      .start_PopNB_mioi_data_rsc_z_mxwt(start_PopNB_mioi_data_rsc_z_mxwt),
      .start_PopNB_mioi_return_rsc_z_mxwt(start_PopNB_mioi_return_rsc_z_mxwt),
      .start_PopNB_mioi_oswt_pff(and_518_rmff)
    );
  PECore_PECore_PECoreRun_rva_out_Push_mioi PECore_PECoreRun_rva_out_Push_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_out_vld(rva_out_vld),
      .rva_out_rdy(rva_out_rdy),
      .rva_out_dat(rva_out_dat),
      .PECoreRun_wen(PECoreRun_wen),
      .rva_out_Push_mioi_oswt(reg_rva_out_Push_mioi_iswt0_cse),
      .rva_out_Push_mioi_wen_comp(rva_out_Push_mioi_wen_comp),
      .rva_out_Push_mioi_m_data_rsc_dat_PECoreRun(nl_PECore_PECoreRun_rva_out_Push_mioi_inst_rva_out_Push_mioi_m_data_rsc_dat_PECoreRun[63:0]),
      .rva_out_Push_mioi_oswt_pff(and_516_cse)
    );
  PECore_PECore_PECoreRun_wait_dp PECore_PECoreRun_wait_dp_inst (
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d),
      .ProductSum_for_acc_11_cmp_en(ProductSum_for_acc_11_cmp_en),
      .ProductSum_for_acc_9_cmp_en(ProductSum_for_acc_9_cmp_en),
      .PECoreRun_wen(PECoreRun_wen),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo(reg_weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_unreg(and_514_rmff),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo(reg_weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_unreg(and_510_rmff),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo(reg_weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_unreg(and_506_rmff),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo(reg_weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_unreg(and_502_rmff),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo(reg_weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_unreg(and_498_rmff),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo(reg_weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_unreg(and_494_rmff),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo(reg_weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_unreg(and_490_rmff),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo(reg_weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_cse),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_unreg(and_487_rmff),
      .ProductSum_for_acc_11_cmp_cgo(reg_PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_cgo_ir_cse),
      .ProductSum_for_acc_11_cmp_cgo_ir_unreg(and_483_rmff),
      .ProductSum_for_acc_9_cmp_cgo(reg_PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_cgo_ir_cse),
      .ProductSum_for_acc_9_cmp_cgo_ir_unreg(and_480_rmff)
    );
  PECore_PECore_PECoreRun_staller PECore_PECoreRun_staller_inst (
      .clk(clk),
      .rst(rst),
      .PECoreRun_wen(PECoreRun_wen),
      .PECoreRun_wten(PECoreRun_wten),
      .act_port_Push_mioi_wen_comp(act_port_Push_mioi_wen_comp),
      .rva_out_Push_mioi_wen_comp(rva_out_Push_mioi_wen_comp)
    );
  PECore_PECore_PECoreRun_PECoreRun_fsm PECore_PECoreRun_PECoreRun_fsm_inst (
      .clk(clk),
      .rst(rst),
      .PECoreRun_wen(PECoreRun_wen),
      .fsm_output(fsm_output)
    );
  assign weight_mem_banks_read_1_for_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_82);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb = weight_mem_banks_read_1_for_mux_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl default clock = (posedge clk);
  // psl weight_mem_banks_load_store_1_for_1_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb );
  assign weight_mem_banks_read_1_for_mux_1_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_82);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb = weight_mem_banks_read_1_for_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb = weight_mem_banks_read_1_for_mux_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_1_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb = weight_mem_banks_read_1_for_mux_1_cse;
  assign weight_mem_banks_read_1_for_mux_4_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_84);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_1 = weight_mem_banks_read_1_for_mux_4_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_1_for_2_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_1  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_1 );
  assign weight_mem_banks_read_1_for_mux_5_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_84);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_1 = weight_mem_banks_read_1_for_mux_5_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_1 = weight_mem_banks_read_1_for_mux_4_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_2_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_1  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_1 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_1 = weight_mem_banks_read_1_for_mux_5_cse;
  assign weight_mem_banks_read_1_for_mux_8_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_86);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_2 = weight_mem_banks_read_1_for_mux_8_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_1_for_3_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_2  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_2 );
  assign weight_mem_banks_read_1_for_mux_9_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_86);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_2 = weight_mem_banks_read_1_for_mux_9_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_2 = weight_mem_banks_read_1_for_mux_8_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_3_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_2  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_2 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_2 = weight_mem_banks_read_1_for_mux_9_cse;
  assign weight_mem_banks_read_1_for_mux_12_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_88);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_3 = weight_mem_banks_read_1_for_mux_12_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_1_for_4_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_3  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_3 );
  assign weight_mem_banks_read_1_for_mux_13_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_88);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_3 = weight_mem_banks_read_1_for_mux_13_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_3 = weight_mem_banks_read_1_for_mux_12_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_4_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_3  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_3 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_3 = weight_mem_banks_read_1_for_mux_13_cse;
  assign weight_mem_banks_read_1_for_mux_16_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_90);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_4 = weight_mem_banks_read_1_for_mux_16_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_1_for_5_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_4  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_4 );
  assign weight_mem_banks_read_1_for_mux_17_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_90);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_4 = weight_mem_banks_read_1_for_mux_17_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_4 = weight_mem_banks_read_1_for_mux_16_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_5_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_4  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_4 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_4 = weight_mem_banks_read_1_for_mux_17_cse;
  assign weight_mem_banks_read_1_for_mux_20_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_92);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_5 = weight_mem_banks_read_1_for_mux_20_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_1_for_6_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_5  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_5 );
  assign weight_mem_banks_read_1_for_mux_21_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_92);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_5 = weight_mem_banks_read_1_for_mux_21_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_5 = weight_mem_banks_read_1_for_mux_20_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_6_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_5  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_5 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_5 = weight_mem_banks_read_1_for_mux_21_cse;
  assign weight_mem_banks_read_1_for_mux_24_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_79);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_6 = weight_mem_banks_read_1_for_mux_24_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_1_for_7_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_6  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_6 );
  assign weight_mem_banks_read_1_for_mux_25_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_79);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_6 = weight_mem_banks_read_1_for_mux_25_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_6 = weight_mem_banks_read_1_for_mux_24_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_7_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_6  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_6 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_6 = weight_mem_banks_read_1_for_mux_25_cse;
  assign weight_mem_banks_read_1_for_mux_28_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_80);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_7 = weight_mem_banks_read_1_for_mux_28_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_1_for_8_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_2 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_7  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_7 );
  assign weight_mem_banks_read_1_for_mux_29_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_80);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_7 = weight_mem_banks_read_1_for_mux_29_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_7 = weight_mem_banks_read_1_for_mux_28_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_1_for_8_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_2 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_7  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_7 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_7 = weight_mem_banks_read_1_for_mux_29_cse;
  assign weight_mem_banks_write_if_for_if_mux_8_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_178);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_8 = weight_mem_banks_write_if_for_if_mux_8_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_1_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_8  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_8 );
  assign weight_mem_banks_write_if_for_if_mux_9_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_178);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_8 = weight_mem_banks_write_if_for_if_mux_9_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_8 = weight_mem_banks_write_if_for_if_mux_8_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_1_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_8  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_8 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_8 = weight_mem_banks_write_if_for_if_mux_9_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb
      = weight_mem_banks_write_if_for_if_mux_8_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_1_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb
      = weight_mem_banks_write_if_for_if_mux_9_cse;
  assign weight_mem_banks_read_for_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_179);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_9 = weight_mem_banks_read_for_mux_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_1_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_9  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_9 );
  assign weight_mem_banks_read_for_mux_1_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_179);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_9 = weight_mem_banks_read_for_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_9 = weight_mem_banks_read_for_mux_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_1_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_9  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_9 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_9 = weight_mem_banks_read_for_mux_1_cse;
  assign weight_mem_banks_write_if_for_if_mux_12_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_181);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_10 = weight_mem_banks_write_if_for_if_mux_12_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_2_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_10  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_10 );
  assign weight_mem_banks_write_if_for_if_mux_13_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_181);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_10 = weight_mem_banks_write_if_for_if_mux_13_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_10 = weight_mem_banks_write_if_for_if_mux_12_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_2_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_10  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_10 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_10 = weight_mem_banks_write_if_for_if_mux_13_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_1
      = weight_mem_banks_write_if_for_if_mux_12_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_2_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_1  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_1 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_1
      = weight_mem_banks_write_if_for_if_mux_13_cse;
  assign weight_mem_banks_read_for_mux_4_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_182);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_11 = weight_mem_banks_read_for_mux_4_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_2_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_11  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_11 );
  assign weight_mem_banks_read_for_mux_5_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_182);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_11 = weight_mem_banks_read_for_mux_5_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_11 = weight_mem_banks_read_for_mux_4_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_2_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_11  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_11 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_11 = weight_mem_banks_read_for_mux_5_cse;
  assign weight_mem_banks_write_if_for_if_mux_16_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_184);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_12 = weight_mem_banks_write_if_for_if_mux_16_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_3_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_12  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_12 );
  assign weight_mem_banks_write_if_for_if_mux_17_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_184);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_12 = weight_mem_banks_write_if_for_if_mux_17_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_12 = weight_mem_banks_write_if_for_if_mux_16_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_3_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_12  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_12 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_12 = weight_mem_banks_write_if_for_if_mux_17_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_2
      = weight_mem_banks_write_if_for_if_mux_16_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_3_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_2  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_2 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_2
      = weight_mem_banks_write_if_for_if_mux_17_cse;
  assign weight_mem_banks_read_for_mux_8_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_185);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_13 = weight_mem_banks_read_for_mux_8_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_3_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_13  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_13 );
  assign weight_mem_banks_read_for_mux_9_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_185);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_13 = weight_mem_banks_read_for_mux_9_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_13 = weight_mem_banks_read_for_mux_8_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_3_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_13  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_13 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_13 = weight_mem_banks_read_for_mux_9_cse;
  assign weight_mem_banks_write_if_for_if_mux_20_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_187);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_14 = weight_mem_banks_write_if_for_if_mux_20_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_4_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_14  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_14 );
  assign weight_mem_banks_write_if_for_if_mux_21_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_187);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_14 = weight_mem_banks_write_if_for_if_mux_21_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_14 = weight_mem_banks_write_if_for_if_mux_20_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_4_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_14  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_14 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_14 = weight_mem_banks_write_if_for_if_mux_21_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_3
      = weight_mem_banks_write_if_for_if_mux_20_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_4_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_3  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_3 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_3
      = weight_mem_banks_write_if_for_if_mux_21_cse;
  assign weight_mem_banks_read_for_mux_12_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_188);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_15 = weight_mem_banks_read_for_mux_12_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_4_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_15  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_15 );
  assign weight_mem_banks_read_for_mux_13_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_188);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_15 = weight_mem_banks_read_for_mux_13_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_15 = weight_mem_banks_read_for_mux_12_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_4_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_15  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_15 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_15 = weight_mem_banks_read_for_mux_13_cse;
  assign weight_mem_banks_write_if_for_if_mux_24_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_190);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_16 = weight_mem_banks_write_if_for_if_mux_24_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_5_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_16  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_16 );
  assign weight_mem_banks_write_if_for_if_mux_25_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_190);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_16 = weight_mem_banks_write_if_for_if_mux_25_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_16 = weight_mem_banks_write_if_for_if_mux_24_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_5_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_16  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_16 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_16 = weight_mem_banks_write_if_for_if_mux_25_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_4
      = weight_mem_banks_write_if_for_if_mux_24_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_5_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_4  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_4 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_4
      = weight_mem_banks_write_if_for_if_mux_25_cse;
  assign weight_mem_banks_read_for_mux_16_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_191);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_17 = weight_mem_banks_read_for_mux_16_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_5_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_17  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_17 );
  assign weight_mem_banks_read_for_mux_17_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_191);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_17 = weight_mem_banks_read_for_mux_17_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_17 = weight_mem_banks_read_for_mux_16_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_5_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_17  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_17 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_17 = weight_mem_banks_read_for_mux_17_cse;
  assign weight_mem_banks_write_if_for_if_mux_28_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_193);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_18 = weight_mem_banks_write_if_for_if_mux_28_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_6_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_18  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_18 );
  assign weight_mem_banks_write_if_for_if_mux_29_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_193);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_18 = weight_mem_banks_write_if_for_if_mux_29_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_18 = weight_mem_banks_write_if_for_if_mux_28_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_6_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_18  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_18 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_18 = weight_mem_banks_write_if_for_if_mux_29_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_5
      = weight_mem_banks_write_if_for_if_mux_28_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_6_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_5  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_5 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_5
      = weight_mem_banks_write_if_for_if_mux_29_cse;
  assign weight_mem_banks_read_for_mux_20_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_194);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_19 = weight_mem_banks_read_for_mux_20_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_6_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_19  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_19 );
  assign weight_mem_banks_read_for_mux_21_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_194);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_19 = weight_mem_banks_read_for_mux_21_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_19 = weight_mem_banks_read_for_mux_20_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_6_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_19  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_19 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_19 = weight_mem_banks_read_for_mux_21_cse;
  assign weight_mem_banks_write_if_for_if_mux_32_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_196);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_20 = weight_mem_banks_write_if_for_if_mux_32_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_7_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_20  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_20 );
  assign weight_mem_banks_write_if_for_if_mux_33_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_196);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_20 = weight_mem_banks_write_if_for_if_mux_33_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_20 = weight_mem_banks_write_if_for_if_mux_32_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_7_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_20  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_20 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_20 = weight_mem_banks_write_if_for_if_mux_33_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_6
      = weight_mem_banks_write_if_for_if_mux_32_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_7_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_6  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_6 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_6
      = weight_mem_banks_write_if_for_if_mux_33_cse;
  assign weight_mem_banks_read_for_mux_24_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_197);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_21 = weight_mem_banks_read_for_mux_24_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_7_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_21  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_21 );
  assign weight_mem_banks_read_for_mux_25_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_197);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_21 = weight_mem_banks_read_for_mux_25_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_21 = weight_mem_banks_read_for_mux_24_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_7_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_21  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_21 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_21 = weight_mem_banks_read_for_mux_25_cse;
  assign weight_mem_banks_write_if_for_if_mux_36_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_199);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_22 = weight_mem_banks_write_if_for_if_mux_36_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl weight_mem_banks_load_store_for_8_PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_22  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_22 );
  assign weight_mem_banks_write_if_for_if_mux_37_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_199);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_22 = weight_mem_banks_write_if_for_if_mux_37_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_22 = weight_mem_banks_write_if_for_if_mux_36_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl weight_mem_banks_load_store_for_8_PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_22  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_22 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_22 = weight_mem_banks_write_if_for_if_mux_37_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_7
      = weight_mem_banks_write_if_for_if_mux_36_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl weight_mem_banks_load_store_for_8_PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_7  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_7 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_7
      = weight_mem_banks_write_if_for_if_mux_37_cse;
  assign weight_mem_banks_read_for_mux_28_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_200);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_23 = weight_mem_banks_read_for_mux_28_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl weight_mem_banks_load_store_for_8_PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_23  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_23 );
  assign weight_mem_banks_read_for_mux_29_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_200);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_23 = weight_mem_banks_read_for_mux_29_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_23 = weight_mem_banks_read_for_mux_28_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl weight_mem_banks_load_store_for_8_PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_23  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_23 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_23 = weight_mem_banks_read_for_mux_29_cse;
  assign input_mem_banks_write_1_if_for_if_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_209);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_24 = input_mem_banks_write_1_if_for_if_mux_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_3 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_24  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_24 );
  assign input_mem_banks_write_1_if_for_if_mux_1_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_209);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_24 = input_mem_banks_write_1_if_for_if_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_24 = input_mem_banks_write_1_if_for_if_mux_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_3 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_24  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_24 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_24 = input_mem_banks_write_1_if_for_if_mux_1_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_8
      = input_mem_banks_write_1_if_for_if_mux_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM_3 : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_8  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_8 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_8
      = input_mem_banks_write_1_if_for_if_mux_1_cse;
  assign input_mem_banks_read_1_for_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_207);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_25 = input_mem_banks_read_1_for_mux_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_3 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_25  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_25 );
  assign input_mem_banks_read_1_for_mux_1_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_207);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_25 = input_mem_banks_read_1_for_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_25 = input_mem_banks_read_1_for_mux_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_3 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_25  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_25 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_25 = input_mem_banks_read_1_for_mux_1_cse;
  assign input_mem_banks_write_if_for_if_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_216);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_26 = input_mem_banks_write_if_for_if_mux_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl PECore_PECoreRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_1 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_26  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_26 );
  assign input_mem_banks_write_if_for_if_mux_1_cse = MUX1HOT_s_1_1_2(PECoreRun_wen,
      and_dcpl_216);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_26 = input_mem_banks_write_if_for_if_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_26 = input_mem_banks_write_if_for_if_mux_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl PECore_PECoreRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_1 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_26  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_26 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_26 = input_mem_banks_write_if_for_if_mux_1_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_9
      = input_mem_banks_write_if_for_if_mux_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl PECore_PECoreRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM_1 : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_9  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb_9 );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb_9
      = input_mem_banks_write_if_for_if_mux_1_cse;
  assign input_mem_banks_read_for_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_219);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_27 = input_mem_banks_read_for_mux_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl PECore_PECoreRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds_1 : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_27  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_27 );
  assign input_mem_banks_read_for_mux_1_cse = MUX1HOT_s_1_1_2(PECoreRun_wen, and_dcpl_219);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_27 = input_mem_banks_read_for_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_27 = input_mem_banks_read_for_mux_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl PECore_PECoreRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds_1 : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_27  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_27 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_27 = input_mem_banks_read_for_mux_1_cse;
  assign and_480_rmff = ((PECore_RunMac_PECore_RunMac_if_and_svs_st_7 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7)
      & while_stage_0_9) | and_dcpl_459) & fsm_output;
  assign and_483_rmff = (and_dcpl_31 | and_dcpl_459) & fsm_output;
  assign mux_191_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1,
      or_tmp_341, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign and_486_nl = while_stage_0_6 & mux_191_nl;
  assign or_945_nl = weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | (~ mux_188_itm);
  assign or_944_nl = or_tmp_341 | (~ mux_188_itm);
  assign mux_189_nl = MUX_s_1_2_2(or_945_nl, or_944_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_190_nl = MUX_s_1_2_2((~ mux_188_itm), mux_189_nl, while_stage_0_6);
  assign mux_192_nl = MUX_s_1_2_2(and_486_nl, mux_190_nl, while_stage_0_7);
  assign and_487_rmff = (mux_192_nl | and_dcpl_467) & fsm_output;
  assign mux_196_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1,
      or_tmp_347, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign and_489_nl = while_stage_0_6 & mux_196_nl;
  assign or_951_nl = weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | not_tmp_312;
  assign or_950_nl = or_tmp_347 | not_tmp_312;
  assign mux_194_nl = MUX_s_1_2_2(or_951_nl, or_950_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_195_nl = MUX_s_1_2_2(not_tmp_312, mux_194_nl, while_stage_0_6);
  assign mux_197_nl = MUX_s_1_2_2(and_489_nl, mux_195_nl, while_stage_0_7);
  assign and_490_rmff = (mux_197_nl | and_dcpl_469) & fsm_output;
  assign or_959_nl = weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_1
      | ProductSum_for_asn_51_itm_3;
  assign mux_202_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp,
      or_959_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_493_nl = while_stage_0_5 & mux_202_nl;
  assign or_958_nl = weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp
      | not_tmp_314;
  assign or_956_nl = weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_1
      | ProductSum_for_asn_51_itm_3;
  assign or_955_nl = (~ or_tmp_352) | weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_1
      | ProductSum_for_asn_51_itm_3;
  assign mux_198_nl = MUX_s_1_2_2(or_956_nl, or_955_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_200_nl = MUX_s_1_2_2(or_958_nl, mux_198_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_201_nl = MUX_s_1_2_2(not_tmp_314, mux_200_nl, while_stage_0_5);
  assign mux_203_nl = MUX_s_1_2_2(and_493_nl, mux_201_nl, while_stage_0_6);
  assign and_494_rmff = (mux_203_nl | and_dcpl_193) & fsm_output;
  assign or_966_nl = weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_1
      | ProductSum_for_asn_42_itm_3;
  assign mux_208_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp,
      or_966_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_497_nl = while_stage_0_5 & mux_208_nl;
  assign or_965_nl = weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp
      | not_tmp_316;
  assign or_963_nl = weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_1
      | ProductSum_for_asn_42_itm_3;
  assign or_962_nl = (~ or_tmp_358) | weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_1
      | ProductSum_for_asn_42_itm_3;
  assign mux_204_nl = MUX_s_1_2_2(or_963_nl, or_962_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_206_nl = MUX_s_1_2_2(or_965_nl, mux_204_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_207_nl = MUX_s_1_2_2(not_tmp_316, mux_206_nl, while_stage_0_5);
  assign mux_209_nl = MUX_s_1_2_2(and_497_nl, mux_207_nl, while_stage_0_6);
  assign and_498_rmff = (mux_209_nl | and_dcpl_190) & fsm_output;
  assign mux_214_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp,
      or_tmp_364, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_501_nl = while_stage_0_5 & mux_214_nl;
  assign or_972_nl = weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp
      | not_tmp_319;
  assign or_971_nl = weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | PECore_RunScale_PECore_RunScale_if_and_1_svs_st_3 | ProductSum_for_asn_25_itm_3;
  assign or_970_nl = or_tmp_364 | (~ or_tmp_365);
  assign mux_210_nl = MUX_s_1_2_2(or_971_nl, or_970_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_212_nl = MUX_s_1_2_2(or_972_nl, mux_210_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_213_nl = MUX_s_1_2_2(not_tmp_319, mux_212_nl, while_stage_0_5);
  assign mux_215_nl = MUX_s_1_2_2(and_501_nl, mux_213_nl, while_stage_0_6);
  assign and_502_rmff = (mux_215_nl | and_dcpl_187) & fsm_output;
  assign or_979_nl = PECore_RunScale_PECore_RunScale_if_and_1_svs_3 | ProductSum_for_asn_16_itm_3;
  assign mux_220_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp,
      or_979_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_505_nl = while_stage_0_5 & mux_220_nl;
  assign or_978_nl = weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp
      | not_tmp_322;
  assign or_976_nl = weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | PECore_RunScale_PECore_RunScale_if_and_1_svs_3 | ProductSum_for_asn_16_itm_3;
  assign or_975_nl = nor_17_cse | PECore_RunScale_PECore_RunScale_if_and_1_svs_3
      | ProductSum_for_asn_16_itm_3;
  assign mux_216_nl = MUX_s_1_2_2(or_976_nl, or_975_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_218_nl = MUX_s_1_2_2(or_978_nl, mux_216_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_219_nl = MUX_s_1_2_2(not_tmp_322, mux_218_nl, while_stage_0_5);
  assign mux_221_nl = MUX_s_1_2_2(and_505_nl, mux_219_nl, while_stage_0_6);
  assign and_506_rmff = (mux_221_nl | and_dcpl_184) & fsm_output;
  assign or_985_nl = PECore_UpdateFSM_switch_lp_equal_tmp_2_3 | PECore_RunMac_PECore_RunMac_if_and_svs_st_3;
  assign mux_226_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp,
      or_985_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_509_nl = while_stage_0_5 & mux_226_nl;
  assign or_984_nl = weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp
      | not_tmp_325;
  assign or_982_nl = weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | PECore_UpdateFSM_switch_lp_equal_tmp_2_3 | PECore_RunMac_PECore_RunMac_if_and_svs_st_3;
  assign or_981_nl = nor_18_cse | PECore_UpdateFSM_switch_lp_equal_tmp_2_3 | PECore_RunMac_PECore_RunMac_if_and_svs_st_3;
  assign mux_222_nl = MUX_s_1_2_2(or_982_nl, or_981_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign mux_224_nl = MUX_s_1_2_2(or_984_nl, mux_222_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_225_nl = MUX_s_1_2_2(not_tmp_325, mux_224_nl, while_stage_0_5);
  assign mux_227_nl = MUX_s_1_2_2(and_509_nl, mux_225_nl, while_stage_0_6);
  assign and_510_rmff = (mux_227_nl | and_dcpl_181) & fsm_output;
  assign or_992_nl = PECore_PushOutput_PECore_PushOutput_if_and_svs_st_3 | PECore_RunFSM_switch_lp_equal_tmp_1_2;
  assign mux_233_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp,
      or_992_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_513_nl = while_stage_0_5 & mux_233_nl;
  assign or_991_nl = weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp
      | (~ mux_230_itm);
  assign or_988_nl = (~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | (~ weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1)))
      | PECore_PushOutput_PECore_PushOutput_if_and_svs_st_3 | PECore_RunFSM_switch_lp_equal_tmp_1_2;
  assign or_987_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | PECore_PushOutput_PECore_PushOutput_if_and_svs_st_3 | PECore_RunFSM_switch_lp_equal_tmp_1_2;
  assign nor_19_nl = ~(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_19_itm_1
      | (~ reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_0_1_itm_2_cse));
  assign mux_228_nl = MUX_s_1_2_2(or_988_nl, or_987_nl, nor_19_nl);
  assign mux_231_nl = MUX_s_1_2_2(or_991_nl, mux_228_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_232_nl = MUX_s_1_2_2((~ mux_230_itm), mux_231_nl, while_stage_0_5);
  assign mux_234_nl = MUX_s_1_2_2(and_513_nl, mux_232_nl, while_stage_0_6);
  assign and_514_rmff = (mux_234_nl | and_dcpl_178) & fsm_output;
  assign and_985_nl = PECore_UpdateFSM_switch_lp_nor_7_itm_1 & PECore_UpdateFSM_switch_lp_equal_tmp_3_1
      & pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_nor_mdf_sva_st_1;
  assign and_705_nl = pe_config_is_zero_first_sva & PECore_UpdateFSM_switch_lp_equal_tmp_2_1
      & pe_manager_zero_active_sva;
  assign mux_498_itm = MUX_s_1_2_2(and_985_nl, PECore_UpdateFSM_switch_lp_nor_7_itm_1,
      and_705_nl);
  assign and_709_nl = start_PopNB_mioi_data_rsc_z_mxwt & start_PopNB_mioi_return_rsc_z_mxwt
      & PECore_UpdateFSM_switch_lp_and_7_itm_1 & pe_config_is_valid_sva;
  assign mux_243_nl = MUX_s_1_2_2(mux_498_itm, PECore_UpdateFSM_switch_lp_nor_7_itm_1,
      and_709_nl);
  assign mux_239_nl = MUX_s_1_2_2(mux_498_itm, PECore_UpdateFSM_switch_lp_nor_7_itm_1,
      and_704_cse);
  assign mux_244_nl = MUX_s_1_2_2(mux_243_nl, mux_239_nl, or_999_cse);
  assign mux_493_nl = MUX_s_1_2_2(mux_498_itm, PECore_UpdateFSM_switch_lp_nor_7_itm_1,
      and_704_cse);
  assign or_997_nl = pe_config_UpdateManagerCounter_if_if_unequal_tmp | (operator_8_false_acc_sdt_sva_1[8]);
  assign mux_240_nl = MUX_s_1_2_2(mux_493_nl, PECore_UpdateFSM_switch_lp_nor_7_itm_1,
      or_997_nl);
  assign or_996_nl = (state_2_1_sva!=2'b10) | state_0_sva;
  assign mux_241_nl = MUX_s_1_2_2(mux_240_nl, PECore_UpdateFSM_switch_lp_nor_7_itm_1,
      or_996_nl);
  assign mux_242_nl = MUX_s_1_2_2(PECore_UpdateFSM_switch_lp_nor_7_itm_1, mux_241_nl,
      pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1);
  assign mux_245_nl = MUX_s_1_2_2(mux_244_nl, mux_242_nl, PECore_UpdateFSM_switch_lp_equal_tmp_5_1);
  assign mux_246_cse = MUX_s_1_2_2(mux_245_nl, state_0_sva, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign mux_247_nl = MUX_s_1_2_2(or_999_cse, mux_246_cse, while_stage_0_3);
  assign or_995_nl = while_stage_0_3 | (state_2_1_sva!=2'b00) | state_0_sva;
  assign or_994_nl = (state_2_1_sva_dfm_1!=2'b00);
  assign mux_248_nl = MUX_s_1_2_2(mux_247_nl, or_995_nl, or_994_nl);
  assign and_518_rmff = (~ mux_248_nl) & and_dcpl_210;
  assign and_520_rmff = while_stage_0_11 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_9)
      & PECore_PushOutput_PECore_PushOutput_if_and_svs_st_9;
  assign PECore_DecodeAxiRead_switch_lp_and_2_cse = PECoreRun_wen & and_dcpl_6;
  assign rva_out_reg_data_and_14_cse = PECoreRun_wen & and_dcpl_6 & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_7
      & (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_3_8) & (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_2_8)
      & (~(PECore_DecodeAxiRead_switch_lp_nor_tmp_8 | rva_in_reg_rw_sva_st_8));
  assign rva_out_reg_data_and_78_enex5 = rva_out_reg_data_and_14_cse & reg_rva_out_reg_data_15_9_sva_dfm_8_enexo;
  assign rva_out_reg_data_and_79_enex5 = rva_out_reg_data_and_14_cse & reg_rva_out_reg_data_23_17_sva_dfm_6_enexo;
  assign rva_out_reg_data_and_80_enex5 = rva_out_reg_data_and_14_cse & reg_rva_out_reg_data_30_25_sva_dfm_6_enexo;
  assign rva_out_reg_data_and_17_cse = PECoreRun_wen & and_dcpl_5;
  assign rva_out_reg_data_and_81_enex5 = rva_out_reg_data_and_17_cse & reg_rva_out_reg_data_62_56_sva_dfm_4_3_enexo;
  assign rva_out_reg_data_and_82_enex5 = rva_out_reg_data_and_17_cse & reg_rva_out_reg_data_55_48_sva_dfm_4_3_enexo;
  assign rva_out_reg_data_and_83_enex5 = rva_out_reg_data_and_17_cse & reg_rva_out_reg_data_55_48_sva_dfm_4_3_1_enexo;
  assign rva_out_reg_data_and_84_enex5 = rva_out_reg_data_and_17_cse & reg_rva_out_reg_data_46_40_sva_dfm_4_3_1_enexo;
  assign rva_out_reg_data_and_85_enex5 = rva_out_reg_data_and_17_cse & reg_rva_out_reg_data_35_32_sva_dfm_4_3_enexo;
  assign input_mem_banks_read_read_data_and_cse = PECoreRun_wen & and_dcpl_5 & (~
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6) & input_read_req_valid_lpi_1_dfm_1_8;
  assign weight_port_read_out_data_and_68_cse = PECoreRun_wen & and_dcpl_4 & (~ rva_in_reg_rw_sva_st_1_8)
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6;
  assign rva_out_reg_data_and_cse = PECoreRun_wen & (~((~(while_stage_0_11 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_9))
      | rva_in_reg_rw_sva_9 | (~ fsm_output)));
  assign input_mem_banks_read_read_data_and_22_enex5 = input_mem_banks_read_read_data_and_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_1_enexo;
  assign input_mem_banks_read_read_data_and_23_enex5 = input_mem_banks_read_read_data_and_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_1_enexo;
  assign input_mem_banks_read_read_data_and_24_enex5 = input_mem_banks_read_read_data_and_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_1_enexo;
  assign weight_port_read_out_data_and_104_enex5 = weight_port_read_out_data_and_68_cse
      & reg_weight_port_read_out_data_0_2_sva_dfm_3_2_enexo;
  assign weight_port_read_out_data_and_105_enex5 = weight_port_read_out_data_and_68_cse
      & reg_weight_port_read_out_data_0_3_sva_dfm_3_2_enexo;
  assign input_mem_banks_read_read_data_and_25_enex5 = input_mem_banks_read_read_data_and_cse
      & reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_1_enexo;
  assign rva_in_reg_rw_and_cse = PECoreRun_wen & while_stage_0_10;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_cse = PECoreRun_wen & and_dcpl_4
      & (~(rva_in_reg_rw_sva_st_1_8 | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6))
      & (~(rva_in_reg_rw_sva_8 | input_read_req_valid_lpi_1_dfm_1_8)) & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_7;
  assign and_1002_cse = (PECore_UpdateFSM_switch_lp_equal_tmp_2_9 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_9
      | (~ while_stage_0_11) | (PECore_RunScale_PECore_RunScale_if_and_1_svs_8 &
      (~ reg_PECore_RunMac_PECore_RunMac_if_and_svs_st_8_cse))) & rva_in_reg_rw_and_cse
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8)
      & (PECore_PushOutput_PECore_PushOutput_if_and_svs_st_8 | (~ PECore_UpdateFSM_switch_lp_equal_tmp_2_8));
  assign PECore_PushOutput_if_and_cse = PECoreRun_wen & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8)
      & while_stage_0_10;
  assign rva_in_reg_rw_and_2_cse = PECoreRun_wen & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7
      & while_stage_0_9;
  assign PECore_RunMac_if_and_cse = PECoreRun_wen & (and_dcpl_27 | and_dcpl_281);
  assign while_if_and_6_cse = PECoreRun_wen & while_stage_0_9;
  assign rva_in_reg_rw_and_3_cse = PECoreRun_wen & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6
      & while_stage_0_8;
  assign PECore_RunMac_if_and_1_cse = PECoreRun_wen & (~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6
      & rva_in_reg_rw_sva_st_1_6)) & while_stage_0_8;
  assign while_if_and_7_cse = PECoreRun_wen & while_stage_0_8;
  assign ProductSum_for_and_cse = PECoreRun_wen & and_dcpl_31;
  assign input_mem_banks_read_1_read_data_and_enex5 = ProductSum_for_and_cse & reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_4_enexo;
  assign input_mem_banks_read_1_read_data_and_6_enex5 = ProductSum_for_and_cse &
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_4_enexo_1;
  assign weight_port_read_out_data_and_enex5 = PECoreRun_wen & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6)
      & while_stage_0_8 & weight_mem_run_3_for_land_3_lpi_1_dfm_3 & fsm_output &
      (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      | (~ while_stage_0_7) | (~ weight_mem_run_3_for_land_3_lpi_1_dfm_2)) & reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_000000;
  assign weight_mem_run_3_for_aelse_and_cse = PECoreRun_wen & while_stage_0_7;
  assign mux_4_nl = MUX_s_1_2_2(or_tmp_3, while_and_24_cse, PECore_RunMac_PECore_RunMac_if_and_svs_st_5);
  assign or_14_nl = (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4) | rva_in_reg_rw_sva_5
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_11_itm_1
      | rva_in_reg_rw_sva_st_1_5 | rva_in_reg_rw_sva_st_5 | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_5
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_5 | PECore_DecodeAxiRead_switch_lp_nor_tmp_5;
  assign mux_5_nl = MUX_s_1_2_2(mux_4_nl, or_tmp_2, or_14_nl);
  assign weight_mem_run_3_for_5_and_209_ssc = PECoreRun_wen & (~ mux_5_nl) & while_stage_0_7;
  assign PECore_RunMac_if_and_2_cse = PECoreRun_wen & (~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      & rva_in_reg_rw_sva_st_1_5)) & while_stage_0_7;
  assign rva_in_reg_rw_and_4_cse = PECoreRun_wen & and_dcpl_40;
  assign weight_mem_banks_read_1_read_data_and_8_cse = PECoreRun_wen & and_dcpl_41;
  assign ProductSum_for_and_8_cse = PECoreRun_wen & reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      & while_stage_0_6;
  assign input_mem_banks_read_1_read_data_and_7_enex5 = ProductSum_for_and_8_cse
      & reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_3_enexo;
  assign weight_port_read_out_data_and_1_cse = PECoreRun_wen & (~(or_dcpl_606 | (~
      weight_mem_run_3_for_land_7_lpi_1_dfm_2)));
  assign weight_mem_run_3_for_aelse_and_1_cse = PECoreRun_wen & while_stage_0_6;
  assign weight_port_read_out_data_and_3_cse = PECoreRun_wen & (~(or_dcpl_606 | (~
      weight_mem_run_3_for_land_5_lpi_1_dfm_2)));
  assign weight_port_read_out_data_and_5_cse = PECoreRun_wen & (~(or_dcpl_606 | (~
      weight_mem_run_3_for_land_4_lpi_1_dfm_2)));
  assign weight_port_read_out_data_and_7_cse = PECoreRun_wen & (~(or_dcpl_606 | (~
      weight_mem_run_3_for_land_3_lpi_1_dfm_2)));
  assign weight_port_read_out_data_and_8_cse = PECoreRun_wen & (~((~ weight_mem_run_3_for_land_2_lpi_1_dfm_2)
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      | (~ while_stage_0_7)));
  assign nor_894_cse = ~((weight_read_addrs_7_lpi_1_dfm_3_2_0[1:0]!=2'b00));
  assign mux_500_nl = MUX_s_1_2_2((weight_read_addrs_7_lpi_1_dfm_3_2_0[1]), (~ (weight_read_addrs_7_lpi_1_dfm_3_2_0[1])),
      weight_read_addrs_7_lpi_1_dfm_3_2_0[0]);
  assign mux_501_cse = MUX_s_1_2_2(mux_500_nl, nor_894_cse, weight_read_addrs_7_lpi_1_dfm_3_2_0[2]);
  assign and_1040_cse = (mux_501_cse | weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_13_itm_2)
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign and_1044_cse = (mux_501_cse | weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_12_itm_1)
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign nor_896_cse = ~((weight_read_addrs_5_lpi_1_dfm_3_2_0[1:0]!=2'b00));
  assign mux_504_nl = MUX_s_1_2_2((weight_read_addrs_5_lpi_1_dfm_3_2_0[1]), (~ (weight_read_addrs_5_lpi_1_dfm_3_2_0[1])),
      weight_read_addrs_5_lpi_1_dfm_3_2_0[0]);
  assign mux_505_nl = MUX_s_1_2_2(mux_504_nl, nor_896_cse, weight_read_addrs_5_lpi_1_dfm_3_2_0[2]);
  assign and_1048_cse = (mux_505_nl | weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_5_itm_2)
      & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign weight_port_read_out_data_and_14_cse = PECoreRun_wen & (and_dcpl_241 | and_dcpl_32);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_101_cse = PECoreRun_wen
      & weight_mem_run_3_for_land_4_lpi_1_dfm_1 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      & while_stage_0_6;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_cse = PECoreRun_wen
      & (weight_mem_run_3_for_land_4_lpi_1_dfm_1 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      & while_stage_0_6;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_105_cse = PECoreRun_wen
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | weight_mem_run_3_for_land_2_lpi_1_dfm_1) & while_stage_0_6;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_108_cse = PECoreRun_wen
      & and_dcpl_41 & weight_mem_run_3_for_land_2_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_cse = PECoreRun_wen & (~
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      & weight_mem_run_3_for_land_1_lpi_1_dfm_2 & while_stage_0_6;
  assign weight_read_addrs_and_7_enex5 = PECoreRun_wen & ((weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_1
      & (~ ProductSum_for_asn_73_itm_3)) | (weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_1
      & (~ ProductSum_for_asn_64_itm_3))) & and_dcpl_69 & reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo;
  assign weight_mem_read_arbxbar_xbar_1_for_3_and_8_cse = PECoreRun_wen & and_dcpl_79;
  assign weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 = weight_mem_read_arbxbar_xbar_1_for_3_and_8_cse
      & (reg_Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1_enexo | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_3_enexo
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_3_enexo
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_3_enexo
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1_enexo
      | reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_1 | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0_enexo
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0_enexo);
  assign weight_mem_read_arbxbar_xbar_1_for_3_and_10_cse = PECoreRun_wen & and_dcpl_80;
  assign weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 = weight_mem_read_arbxbar_xbar_1_for_3_and_10_cse
      & (reg_Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1_enexo_1 | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0_enexo_1
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_3_enexo_1
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_0_enexo
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0_enexo_1
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_3_enexo_1
      | reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_2 | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_3_enexo_1
      | reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1_enexo_1
      | reg_weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs_enexo);
  assign while_if_and_10_cse = PECoreRun_wen & while_stage_0_5;
  assign weight_mem_read_arbxbar_arbiters_next_and_cse = PECoreRun_wen & fsm_output;
  assign weight_mem_read_arbxbar_arbiters_next_and_50_cse = weight_mem_read_arbxbar_arbiters_next_and_cse
      & (and_100_cse | or_dcpl_13);
  assign weight_mem_read_arbxbar_arbiters_next_and_56_cse = weight_mem_read_arbxbar_arbiters_next_and_cse
      & ((nor_228_cse & nor_229_cse & nor_230_cse & nor_231_cse) | or_dcpl_13);
  assign weight_mem_read_arbxbar_arbiters_next_and_62_cse = weight_mem_read_arbxbar_arbiters_next_and_cse
      & or_dcpl_16;
  assign weight_mem_read_arbxbar_arbiters_next_and_67_cse = weight_mem_read_arbxbar_arbiters_next_and_cse
      & ((nor_236_cse & nor_237_cse & nor_238_cse & nor_239_cse) | or_dcpl_13);
  assign weight_mem_read_arbxbar_arbiters_next_and_73_cse = weight_mem_read_arbxbar_arbiters_next_and_cse
      & ((nor_240_cse & nor_241_cse & nor_242_cse & nor_243_cse) | or_dcpl_13);
  assign weight_mem_read_arbxbar_arbiters_next_and_79_cse = weight_mem_read_arbxbar_arbiters_next_and_cse
      & ((nor_244_cse & nor_245_cse & nor_246_cse & nor_247_cse) | or_dcpl_13);
  assign weight_mem_read_arbxbar_arbiters_next_and_85_cse = weight_mem_read_arbxbar_arbiters_next_and_cse
      & ((nor_248_cse & nor_249_cse & nor_250_cse & nor_251_cse) | or_dcpl_13);
  assign weight_mem_read_arbxbar_arbiters_next_and_91_cse = weight_mem_read_arbxbar_arbiters_next_and_cse
      & or_dcpl_21;
  assign nand_372_cse = ~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & reg_rva_in_reg_rw_sva_st_1_1_cse);
  assign weight_read_addrs_and_9_cse = PECoreRun_wen & (and_dcpl_156 | and_dcpl_155
      | and_dcpl_154 | and_dcpl_153 | and_dcpl_152 | and_dcpl_151 | and_dcpl_150
      | and_dcpl_149 | (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2))
      & while_stage_0_4;
  assign weight_write_data_data_and_cse = PECoreRun_wen & ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[7:6]!=2'b00))
      & and_dcpl_162;
  assign weight_write_data_data_and_24_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_7_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_25_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_6_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_26_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_5_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_27_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_4_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_28_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_3_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_29_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_2_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_30_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_1_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_data_data_and_31_enex5 = weight_write_data_data_and_cse & reg_weight_write_data_data_0_0_lpi_1_dfm_1_2_6_enexo;
  assign weight_write_addrs_and_enex5 = weight_write_data_data_and_cse & reg_weight_write_addrs_lpi_1_dfm_1_2_enexo;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_cse
      = PECoreRun_wen & and_dcpl_168;
  assign PECore_RunFSM_switch_lp_and_cse = PECoreRun_wen & while_stage_0_4;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_13_cse
      = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_10 & and_dcpl_168;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_14_cse
      = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11 & and_dcpl_168;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_18_cse
      = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_12 & and_dcpl_168;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_22_cse
      = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_13 & and_dcpl_168;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_26_cse
      = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_14 & and_dcpl_168;
  assign Arbiter_8U_Roundrobin_pick_1_and_15_cse = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8
      & and_dcpl_168;
  assign weight_mem_read_arbxbar_xbar_requests_transpose_and_14_cse = PECoreRun_wen
      & and_dcpl_162;
  assign Arbiter_8U_Roundrobin_pick_and_cse = PECoreRun_wen & (while_stage_0_4 |
      and_dcpl_525) & fsm_output & or_dcpl_13;
  assign Arbiter_8U_Roundrobin_pick_1_and_22_cse = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9
      & and_dcpl_168;
  assign Arbiter_8U_Roundrobin_pick_1_and_64_cse = PECoreRun_wen & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_15
      & and_dcpl_168;
  assign weight_write_data_data_and_8_cse = PECoreRun_wen & and_dcpl_203;
  assign weight_write_data_data_and_32_enex5 = weight_write_data_data_and_8_cse &
      reg_weight_write_data_data_0_7_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_33_enex5 = weight_write_data_data_and_8_cse &
      reg_weight_write_data_data_0_6_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_34_enex5 = weight_write_data_data_and_8_cse &
      reg_weight_write_data_data_0_5_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_35_enex5 = weight_write_data_data_and_8_cse &
      reg_weight_write_data_data_0_4_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_36_enex5 = weight_write_data_data_and_8_cse &
      reg_weight_write_data_data_0_3_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_37_enex5 = weight_write_data_data_and_8_cse &
      reg_weight_write_data_data_0_2_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_38_enex5 = weight_write_data_data_and_8_cse &
      reg_weight_write_data_data_0_1_lpi_1_dfm_1_1_enexo;
  assign weight_write_data_data_and_39_enex5 = weight_write_data_data_and_8_cse &
      reg_weight_write_data_data_0_0_lpi_1_dfm_1_1_enexo;
  assign weight_write_addrs_and_2_enex5 = weight_write_data_data_and_8_cse & reg_pe_manager_base_input_enexo;
  assign PECore_DecodeAxiWrite_switch_lp_and_2_cse = PECoreRun_wen & while_stage_0_3;
  assign weight_read_addrs_and_28_enex5 = weight_write_data_data_and_8_cse & reg_weight_read_addrs_0_3_0_lpi_1_dfm_1_1_enexo;
  assign state_and_cse = weight_mem_read_arbxbar_arbiters_next_and_cse & or_dcpl_87;
  assign nor_910_cse = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[15:14]!=2'b00));
  assign nor_907_cse = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[10:8]!=3'b000));
  assign nor_909_cse = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[13:11]!=3'b000));
  assign and_1065_cse = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & PECore_UpdateFSM_switch_lp_equal_tmp_5_1 & while_stage_0_3;
  assign pe_config_num_manager_and_cse = PECoreRun_wen & (~(or_dcpl_628 | or_dcpl_627
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) | (~(PECore_DecodeAxiRead_case_4_switch_lp_nor_8_tmp
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])))));
  assign rva_in_reg_rw_and_6_cse = PECoreRun_wen & reg_rva_in_PopNB_mioi_iswt0_cse;
  assign PECore_UpdateFSM_switch_lp_and_9_cse = PECoreRun_wen & and_dcpl_210;
  assign or_1491_cse = (~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17:16]!=2'b00) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:18]!=2'b01);
  assign nor_912_cse = ~((~ reg_rva_in_reg_rw_sva_st_1_1_cse) | PECore_DecodeAxiWrite_switch_lp_nor_tmp_1
      | PECore_DecodeAxiWrite_switch_lp_equal_tmp_2 | PECore_DecodeAxiWrite_switch_lp_equal_tmp_1);
  assign and_2257_cse = PECore_UpdateFSM_switch_lp_equal_tmp_5_1 & pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1;
  assign pe_config_UpdateManagerCounter_if_if_and_enex5 = PECoreRun_wen & reg_pe_config_num_output_enexo;
  assign PECore_DecodeAxiRead_switch_lp_and_cse = PECoreRun_wen & (~(or_dcpl_87 |
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt));
  assign PECore_DecodeAxiWrite_switch_lp_and_cse = PECoreRun_wen & (~ or_dcpl_627);
  assign and_1098_cse = ((~ while_stage_0_10) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8)
      & while_stage_0_11 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_9)
      & fsm_output & PECoreRun_wen;
  assign weight_port_read_out_data_and_92_cse = PECoreRun_wen & and_dcpl_221 & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5
      & while_stage_0_9;
  assign nor_259_nl = ~(and_692_cse | (state_2_1_sva[1]) | (~((state_2_1_sva[0])
      & state_0_sva)));
  assign nor_260_nl = ~(PECore_UpdateFSM_switch_lp_equal_tmp_3_1 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      | (~ PECore_RunScale_PECore_RunScale_if_and_1_svs_1_1));
  assign mux_20_nl = MUX_s_1_2_2(nor_259_nl, nor_260_nl, while_stage_0_3);
  assign nor_261_nl = ~(or_tmp_33 | (~ PECore_RunScale_PECore_RunScale_if_and_1_svs_st_2));
  assign mux_21_nl = MUX_s_1_2_2(mux_20_nl, nor_261_nl, while_stage_0_4);
  assign nor_262_nl = ~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | PECore_RunMac_PECore_RunMac_if_and_svs_st_3 | (~(PECore_RunScale_PECore_RunScale_if_and_1_svs_st_3
      & PECore_RunScale_PECore_RunScale_if_and_1_svs_3)));
  assign mux_22_nl = MUX_s_1_2_2(mux_21_nl, nor_262_nl, while_stage_0_5);
  assign nor_263_nl = ~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | (~ reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_3_1_itm_2_cse)
      | (~ reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_2_1_itm_2_cse)
      | reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse);
  assign mux_23_nl = MUX_s_1_2_2(mux_22_nl, nor_263_nl, while_stage_0_6);
  assign nor_264_nl = ~((~ PECore_RunScale_PECore_RunScale_if_and_1_svs_st_5) | (~
      PECore_RunScale_PECore_RunScale_if_and_1_svs_5) | PECore_RunMac_PECore_RunMac_if_and_svs_st_5
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign mux_24_nl = MUX_s_1_2_2(mux_23_nl, nor_264_nl, while_stage_0_7);
  assign nor_265_nl = ~((~ PECore_RunScale_PECore_RunScale_if_and_1_svs_st_6) | (~
      PECore_RunScale_PECore_RunScale_if_and_1_svs_6) | PECore_RunMac_PECore_RunMac_if_and_svs_st_6
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6);
  assign mux_25_nl = MUX_s_1_2_2(mux_24_nl, nor_265_nl, while_stage_0_8);
  assign nor_266_nl = ~((~ PECore_RunScale_PECore_RunScale_if_and_1_svs_7) | (~ PECore_RunScale_PECore_RunScale_if_and_1_svs_st_7)
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7
      | PECore_RunMac_PECore_RunMac_if_and_svs_st_7);
  assign mux_26_nl = MUX_s_1_2_2(mux_25_nl, nor_266_nl, while_stage_0_9);
  assign accum_vector_data_and_40_cse = rva_in_reg_rw_and_cse & mux_26_nl;
  assign PECore_RunScale_if_and_cse = PECoreRun_wen & and_dcpl_27;
  assign weight_mem_banks_load_store_for_else_and_cse = PECoreRun_wen & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_44_itm_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & while_stage_0_6;
  assign weight_mem_banks_load_store_for_else_and_1_cse = PECoreRun_wen & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_46_itm_1 & while_stage_0_6;
  assign weight_mem_banks_load_store_for_else_and_2_cse = PECoreRun_wen & and_dcpl_228
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_tmp
      & while_stage_0_6;
  assign and_1129_cse = (((weight_read_addrs_7_lpi_1_dfm_3_2_0[1]) ^ (weight_read_addrs_7_lpi_1_dfm_3_2_0[0])
      ^ (weight_read_addrs_7_lpi_1_dfm_3_2_0[2])) | weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_12_itm_1)
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign and_1138_cse = (and_1040_cse | or_dcpl_751 | weight_mem_run_3_for_5_and_156_itm_2
      | weight_mem_run_3_for_5_and_112_itm_1) & while_stage_0_7 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
      & PECoreRun_wen;
  assign xor_7_cse = (weight_read_addrs_5_lpi_1_dfm_3_2_0[1]) ^ (weight_read_addrs_5_lpi_1_dfm_3_2_0[0])
      ^ (weight_read_addrs_5_lpi_1_dfm_3_2_0[2]);
  assign and_1162_cse = (and_1048_cse | weight_mem_run_3_for_5_and_47_itm_1 | weight_mem_run_3_for_5_and_38_itm_1
      | or_dcpl_727) & while_stage_0_7 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
      & PECoreRun_wen;
  assign and_1166_cse = (((xor_7_cse | weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_5_itm_2)
      & weight_mem_run_3_for_land_6_lpi_1_dfm_2) | or_dcpl_779 | weight_mem_run_3_for_5_and_44_itm_2)
      & while_stage_0_7 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
      & PECoreRun_wen;
  assign xor_13_cse = (weight_read_addrs_3_lpi_1_dfm_3_2_0[1]) ^ (weight_read_addrs_3_lpi_1_dfm_3_2_0[0])
      ^ (weight_read_addrs_3_lpi_1_dfm_3_2_0[2]);
  assign and_1177_cse = (xor_13_cse | weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_3_itm_1)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign weight_port_read_out_data_and_60_cse = PECoreRun_wen & ((weight_mem_run_3_for_land_1_lpi_1_dfm_3
      & while_stage_0_7) | and_dcpl_241);
  assign weight_read_addrs_and_19_cse = PECoreRun_wen & and_dcpl_78;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_30_cse
      = weight_mem_read_arbxbar_arbiters_next_and_cse & or_dcpl_13;
  assign weight_read_addrs_and_29_enex5 = weight_write_data_data_and_8_cse & reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_1_enexo;
  assign operator_15_false_1_and_cse = PECoreRun_wen & (~(and_100_cse | or_dcpl_13));
  assign PEManager_15U_PEManagerWrite_and_enex5 = PECoreRun_wen & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & reg_rva_in_reg_rw_sva_st_1_1_cse & (~(PECore_DecodeAxiWrite_switch_lp_equal_tmp_2
      | PECore_DecodeAxiWrite_switch_lp_nor_tmp_1)) & (~ PECore_DecodeAxiWrite_switch_lp_equal_tmp_1)
      & PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_1_1 & while_stage_0_3 &
      reg_rva_in_reg_data_sva_1_enexo;
  assign pe_manager_num_input_and_cse = PECoreRun_wen & (~(or_dcpl_628 | or_dcpl_87
      | or_dcpl_658));
  assign pe_config_is_valid_and_cse = PECoreRun_wen & (~(PECore_DecodeAxiWrite_case_4_switch_lp_or_cse_1
      | PECore_DecodeAxiWrite_switch_lp_or_5_cse_1)) & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (~ or_dcpl_87);
  assign nor_922_cse = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7:6]!=2'b00));
  assign nor_536_cse = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])));
  assign while_if_and_14_cse = PECoreRun_wen & and_692_cse;
  assign rva_in_reg_rw_and_7_cse = PECoreRun_wen & and_dcpl_69;
  assign rva_in_reg_rw_and_8_cse = PECoreRun_wen & and_dcpl_241;
  assign ProductSum_for_and_16_cse = PECoreRun_wen & and_dcpl_246;
  assign or_162_cse = Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_30_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_2_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_18_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_6_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_10_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_14_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_26_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_22_tmp;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_122_cse = PECoreRun_wen
      & (weight_mem_run_3_for_land_4_lpi_1_dfm_1_1 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_cse = PECoreRun_wen
      & (weight_mem_run_3_for_land_2_lpi_1_dfm_1_1 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_72_cse = PECoreRun_wen
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_73_cse = PECoreRun_wen
      & (weight_mem_run_3_for_land_1_lpi_1_dfm_1 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign input_mem_banks_read_read_data_and_9_cse = PECoreRun_wen & and_dcpl_266
      & input_read_req_valid_lpi_1_dfm_1_7 & while_stage_0_9;
  assign input_mem_banks_read_read_data_and_26_enex5 = input_mem_banks_read_read_data_and_9_cse
      & reg_input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0_enexo;
  assign input_mem_banks_read_read_data_and_27_enex5 = input_mem_banks_read_read_data_and_9_cse
      & reg_input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0_enexo_1;
  assign input_mem_banks_read_read_data_and_28_enex5 = input_mem_banks_read_read_data_and_9_cse
      & reg_input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0_enexo_2;
  assign input_mem_banks_read_read_data_and_29_enex5 = input_mem_banks_read_read_data_and_9_cse
      & reg_input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0_enexo_3;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_4_cse = PECoreRun_wen & and_dcpl_221
      & (~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5 | rva_in_reg_rw_sva_7))
      & (~ input_read_req_valid_lpi_1_dfm_1_7) & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_6
      & while_stage_0_9;
  assign input_mem_banks_read_1_read_data_and_3_enex5 = PECoreRun_wen & (and_dcpl_246
      | (and_dcpl_376 & input_read_req_valid_lpi_1_dfm_1_3 & and_dcpl_69)) & reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_2_enexo;
  assign or_186_cse = Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_113_tmp
      | and_702_cse | and_703_cse | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_101_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_77_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_65_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_53_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_89_tmp;
  assign or_196_cse = Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_124_tmp
      | and_700_cse | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_100_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_112_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_64_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_88_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_52_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_76_tmp;
  assign input_read_req_valid_and_1_cse = PECoreRun_wen & and_dcpl_281;
  assign PECore_DecodeAxiRead_switch_lp_and_7_cse = PECoreRun_wen & and_dcpl_266
      & and_dcpl_282 & while_stage_0_9;
  assign rva_out_reg_data_and_24_cse = PECoreRun_wen & and_dcpl_266 & and_dcpl_282
      & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_6 & (~(rva_in_reg_rw_sva_st_7
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_7 | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_7))
      & (~ PECore_DecodeAxiRead_switch_lp_nor_tmp_7) & while_stage_0_9;
  assign rva_out_reg_data_and_86_enex5 = rva_out_reg_data_and_24_cse & reg_rva_out_reg_data_30_25_sva_dfm_5_enexo;
  assign rva_out_reg_data_and_87_enex5 = rva_out_reg_data_and_24_cse & reg_rva_out_reg_data_23_17_sva_dfm_5_enexo;
  assign rva_out_reg_data_and_88_enex5 = rva_out_reg_data_and_24_cse & reg_rva_out_reg_data_15_9_sva_dfm_7_enexo;
  assign rva_out_reg_data_and_89_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_35_32_sva_dfm_4_2_enexo;
  assign rva_out_reg_data_and_90_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_62_56_sva_dfm_4_2_enexo;
  assign nor_340_cse = ~(state_0_sva | (state_2_1_sva[1]));
  assign mux_531_nl = MUX_s_1_2_2((~ state_0_sva), state_0_sva, state_2_1_sva[0]);
  assign nor_929_cse = ~((state_2_1_sva[1]) | mux_531_nl);
  assign or_1608_nl = rva_in_PopNB_mioi_return_rsc_z_mxwt | (~(reg_rva_in_PopNB_mioi_iswt0_cse
      & (accum_vector_data_7_sva_1_load | nor_929_cse)));
  assign or_1605_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      | (~(accum_vector_data_7_sva_1_load | PECore_UpdateFSM_switch_lp_equal_tmp_3_1
      | PECore_UpdateFSM_switch_lp_equal_tmp_2_1));
  assign mux_532_nl = MUX_s_1_2_2(or_1608_nl, or_1605_nl, while_stage_0_3);
  assign or_1603_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      | (~(accum_vector_operator_1_for_asn_70_itm_1 | PECore_RunMac_PECore_RunMac_if_and_svs_st_2));
  assign mux_533_nl = MUX_s_1_2_2(mux_532_nl, or_1603_nl, while_stage_0_4);
  assign or_1601_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(accum_vector_operator_1_for_asn_70_itm_2 | PECore_RunMac_PECore_RunMac_if_and_svs_st_3));
  assign mux_534_nl = MUX_s_1_2_2(mux_533_nl, or_1601_nl, while_stage_0_5);
  assign or_1599_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | (~(accum_vector_operator_1_for_asn_70_itm_3 | reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse));
  assign mux_535_nl = MUX_s_1_2_2(mux_534_nl, or_1599_nl, while_stage_0_6);
  assign or_1597_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      | (~(PECore_RunMac_PECore_RunMac_if_and_svs_st_5 | accum_vector_operator_1_for_asn_70_itm_4));
  assign mux_536_nl = MUX_s_1_2_2(mux_535_nl, or_1597_nl, while_stage_0_7);
  assign or_1595_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6
      | (~(PECore_RunMac_PECore_RunMac_if_and_svs_st_6 | accum_vector_operator_1_for_asn_70_itm_5));
  assign mux_537_cse = MUX_s_1_2_2(mux_536_nl, or_1595_nl, while_stage_0_8);
  assign or_1627_nl = rva_in_PopNB_mioi_return_rsc_z_mxwt | (~(reg_rva_in_PopNB_mioi_iswt0_cse
      & (accum_vector_data_6_sva_1_load | nor_929_cse)));
  assign or_1624_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      | (~(accum_vector_data_6_sva_1_load | PECore_UpdateFSM_switch_lp_equal_tmp_3_1
      | PECore_UpdateFSM_switch_lp_equal_tmp_2_1));
  assign mux_540_nl = MUX_s_1_2_2(or_1627_nl, or_1624_nl, while_stage_0_3);
  assign or_1622_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      | (~(PECore_DecodeAxiWrite_switch_lp_equal_tmp_1_2 | PECore_RunMac_PECore_RunMac_if_and_svs_st_2));
  assign mux_541_nl = MUX_s_1_2_2(mux_540_nl, or_1622_nl, while_stage_0_4);
  assign or_1620_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(accum_vector_operator_1_for_asn_61_itm_2 | PECore_RunMac_PECore_RunMac_if_and_svs_st_3));
  assign mux_542_nl = MUX_s_1_2_2(mux_541_nl, or_1620_nl, while_stage_0_5);
  assign or_1618_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | (~(accum_vector_operator_1_for_asn_61_itm_3 | reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse));
  assign mux_543_nl = MUX_s_1_2_2(mux_542_nl, or_1618_nl, while_stage_0_6);
  assign or_1616_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      | (~(PECore_RunMac_PECore_RunMac_if_and_svs_st_5 | accum_vector_operator_1_for_asn_61_itm_4));
  assign mux_544_nl = MUX_s_1_2_2(mux_543_nl, or_1616_nl, while_stage_0_7);
  assign or_1614_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6
      | (~(PECore_RunMac_PECore_RunMac_if_and_svs_st_6 | accum_vector_operator_1_for_asn_61_itm_5));
  assign mux_545_cse = MUX_s_1_2_2(mux_544_nl, or_1614_nl, while_stage_0_8);
  assign or_1647_nl = rva_in_PopNB_mioi_return_rsc_z_mxwt | (~(reg_rva_in_PopNB_mioi_iswt0_cse
      & (accum_vector_data_5_sva_1_load | nor_929_cse)));
  assign or_1644_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      | (~(accum_vector_data_5_sva_1_load | PECore_UpdateFSM_switch_lp_equal_tmp_3_1
      | PECore_UpdateFSM_switch_lp_equal_tmp_2_1));
  assign mux_548_nl = MUX_s_1_2_2(or_1647_nl, or_1644_nl, while_stage_0_3);
  assign or_1642_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      | (~(PECore_DecodeAxiRead_switch_lp_nor_tmp_2 | PECore_RunMac_PECore_RunMac_if_and_svs_st_2));
  assign mux_549_nl = MUX_s_1_2_2(mux_548_nl, or_1642_nl, while_stage_0_4);
  assign or_1640_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(PECore_DecodeAxiRead_switch_lp_nor_tmp_3 | PECore_RunMac_PECore_RunMac_if_and_svs_st_3));
  assign mux_550_nl = MUX_s_1_2_2(mux_549_nl, or_1640_nl, while_stage_0_5);
  assign or_1638_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | (~(accum_vector_operator_1_for_asn_52_itm_3 | reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse));
  assign mux_551_nl = MUX_s_1_2_2(mux_550_nl, or_1638_nl, while_stage_0_6);
  assign or_1636_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      | (~(PECore_RunMac_PECore_RunMac_if_and_svs_st_5 | accum_vector_operator_1_for_asn_52_itm_4));
  assign mux_552_nl = MUX_s_1_2_2(mux_551_nl, or_1636_nl, while_stage_0_7);
  assign or_1634_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6
      | (~(PECore_RunMac_PECore_RunMac_if_and_svs_st_6 | accum_vector_operator_1_for_asn_52_itm_5));
  assign mux_553_cse = MUX_s_1_2_2(mux_552_nl, or_1634_nl, while_stage_0_8);
  assign or_1665_nl = rva_in_PopNB_mioi_return_rsc_z_mxwt | (~(reg_rva_in_PopNB_mioi_iswt0_cse
      & (accum_vector_data_4_sva_1_load | nor_929_cse)));
  assign or_1662_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      | (~(accum_vector_data_4_sva_1_load | PECore_UpdateFSM_switch_lp_equal_tmp_3_1
      | PECore_UpdateFSM_switch_lp_equal_tmp_2_1));
  assign mux_556_nl = MUX_s_1_2_2(or_1665_nl, or_1662_nl, while_stage_0_3);
  assign or_1660_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      | (~(PECore_DecodeAxiRead_switch_lp_equal_tmp_3_2 | PECore_RunMac_PECore_RunMac_if_and_svs_st_2));
  assign mux_557_nl = MUX_s_1_2_2(mux_556_nl, or_1660_nl, while_stage_0_4);
  assign or_1658_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(PECore_DecodeAxiRead_switch_lp_equal_tmp_3_3 | PECore_RunMac_PECore_RunMac_if_and_svs_st_3));
  assign mux_558_nl = MUX_s_1_2_2(mux_557_nl, or_1658_nl, while_stage_0_5);
  assign or_1656_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | (~(accum_vector_operator_1_for_asn_43_itm_3 | reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse));
  assign mux_559_nl = MUX_s_1_2_2(mux_558_nl, or_1656_nl, while_stage_0_6);
  assign or_1654_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      | (~(PECore_RunMac_PECore_RunMac_if_and_svs_st_5 | accum_vector_operator_1_for_asn_43_itm_4));
  assign mux_560_nl = MUX_s_1_2_2(mux_559_nl, or_1654_nl, while_stage_0_7);
  assign or_1652_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6
      | (~(PECore_RunMac_PECore_RunMac_if_and_svs_st_6 | accum_vector_operator_1_for_asn_43_itm_5));
  assign mux_561_cse = MUX_s_1_2_2(mux_560_nl, or_1652_nl, while_stage_0_8);
  assign or_1650_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7
      | (~ or_tmp_796);
  assign mux_562_nl = MUX_s_1_2_2(mux_561_cse, or_1650_nl, while_stage_0_9);
  assign and_1250_cse = mux_562_nl & and_dcpl_885 & PECoreRun_wen & (accum_vector_operator_1_for_asn_37_itm_7
      | reg_PECore_RunMac_PECore_RunMac_if_and_svs_st_8_cse) & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign or_1701_nl = rva_in_PopNB_mioi_return_rsc_z_mxwt | (~(reg_rva_in_PopNB_mioi_iswt0_cse
      & (accum_vector_data_3_sva_1_load | nor_929_cse)));
  assign or_1698_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      | (~(accum_vector_data_3_sva_1_load | PECore_UpdateFSM_switch_lp_equal_tmp_3_1
      | PECore_UpdateFSM_switch_lp_equal_tmp_2_1));
  assign mux_572_nl = MUX_s_1_2_2(or_1701_nl, or_1698_nl, while_stage_0_3);
  assign or_1696_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      | (~(PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_2 | PECore_RunMac_PECore_RunMac_if_and_svs_st_2));
  assign mux_573_nl = MUX_s_1_2_2(mux_572_nl, or_1696_nl, while_stage_0_4);
  assign or_1694_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(accum_vector_operator_1_for_asn_34_itm_2 | PECore_RunMac_PECore_RunMac_if_and_svs_st_3));
  assign mux_574_nl = MUX_s_1_2_2(mux_573_nl, or_1694_nl, while_stage_0_5);
  assign or_1692_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | (~(accum_vector_operator_1_for_asn_34_itm_3 | reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse));
  assign mux_575_nl = MUX_s_1_2_2(mux_574_nl, or_1692_nl, while_stage_0_6);
  assign or_1690_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      | (~(PECore_RunMac_PECore_RunMac_if_and_svs_st_5 | accum_vector_operator_1_for_asn_34_itm_4));
  assign mux_576_nl = MUX_s_1_2_2(mux_575_nl, or_1690_nl, while_stage_0_7);
  assign or_1688_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6
      | (~(PECore_RunMac_PECore_RunMac_if_and_svs_st_6 | accum_vector_operator_1_for_asn_34_itm_5));
  assign mux_577_cse = MUX_s_1_2_2(mux_576_nl, or_1688_nl, while_stage_0_8);
  assign or_1686_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7
      | (~ or_tmp_830);
  assign mux_578_nl = MUX_s_1_2_2(mux_577_cse, or_1686_nl, while_stage_0_9);
  assign and_1262_cse = mux_578_nl & and_dcpl_885 & PECoreRun_wen & (accum_vector_operator_1_for_asn_28_itm_7
      | reg_PECore_RunMac_PECore_RunMac_if_and_svs_st_8_cse) & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign or_1737_nl = rva_in_PopNB_mioi_return_rsc_z_mxwt | (~(reg_rva_in_PopNB_mioi_iswt0_cse
      & (accum_vector_data_2_sva_1_load | nor_929_cse)));
  assign or_1734_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      | (~(accum_vector_data_2_sva_1_load | PECore_UpdateFSM_switch_lp_equal_tmp_3_1
      | PECore_UpdateFSM_switch_lp_equal_tmp_2_1));
  assign mux_588_nl = MUX_s_1_2_2(or_1737_nl, or_1734_nl, while_stage_0_3);
  assign or_1732_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      | (~(PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_2 | PECore_RunMac_PECore_RunMac_if_and_svs_st_2));
  assign mux_589_nl = MUX_s_1_2_2(mux_588_nl, or_1732_nl, while_stage_0_4);
  assign or_1730_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(accum_vector_operator_1_for_asn_25_itm_2 | PECore_RunMac_PECore_RunMac_if_and_svs_st_3));
  assign mux_590_nl = MUX_s_1_2_2(mux_589_nl, or_1730_nl, while_stage_0_5);
  assign or_1728_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | (~(accum_vector_operator_1_for_asn_25_itm_3 | reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse));
  assign mux_591_nl = MUX_s_1_2_2(mux_590_nl, or_1728_nl, while_stage_0_6);
  assign or_1726_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      | (~(PECore_RunMac_PECore_RunMac_if_and_svs_st_5 | accum_vector_operator_1_for_asn_25_itm_4));
  assign mux_592_nl = MUX_s_1_2_2(mux_591_nl, or_1726_nl, while_stage_0_7);
  assign or_1724_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6
      | (~(PECore_RunMac_PECore_RunMac_if_and_svs_st_6 | accum_vector_operator_1_for_asn_25_itm_5));
  assign mux_593_nl = MUX_s_1_2_2(mux_592_nl, or_1724_nl, while_stage_0_8);
  assign or_1722_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7
      | (~ or_tmp_864);
  assign mux_594_nl = MUX_s_1_2_2(mux_593_nl, or_1722_nl, while_stage_0_9);
  assign and_1274_cse = mux_594_nl & and_dcpl_885 & PECoreRun_wen & (accum_vector_operator_1_for_asn_22_itm_7
      | reg_PECore_RunMac_PECore_RunMac_if_and_svs_st_8_cse) & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign or_1791_nl = rva_in_PopNB_mioi_return_rsc_z_mxwt | (~(reg_rva_in_PopNB_mioi_iswt0_cse
      & (accum_vector_data_1_sva_1_load | nor_929_cse)));
  assign or_1788_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      | (~(accum_vector_data_1_sva_1_load | PECore_UpdateFSM_switch_lp_equal_tmp_3_1
      | PECore_UpdateFSM_switch_lp_equal_tmp_2_1));
  assign mux_612_nl = MUX_s_1_2_2(or_1791_nl, or_1788_nl, while_stage_0_3);
  assign or_1786_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      | (~(PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_2 | PECore_RunMac_PECore_RunMac_if_and_svs_st_2));
  assign mux_613_nl = MUX_s_1_2_2(mux_612_nl, or_1786_nl, while_stage_0_4);
  assign or_1784_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(accum_vector_operator_1_for_asn_16_itm_2 | PECore_RunMac_PECore_RunMac_if_and_svs_st_3));
  assign mux_614_nl = MUX_s_1_2_2(mux_613_nl, or_1784_nl, while_stage_0_5);
  assign or_1782_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | (~(accum_vector_operator_1_for_asn_16_itm_3 | reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse));
  assign mux_615_nl = MUX_s_1_2_2(mux_614_nl, or_1782_nl, while_stage_0_6);
  assign or_1780_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      | (~(PECore_RunMac_PECore_RunMac_if_and_svs_st_5 | accum_vector_operator_1_for_asn_16_itm_4));
  assign mux_616_nl = MUX_s_1_2_2(mux_615_nl, or_1780_nl, while_stage_0_7);
  assign or_1778_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6
      | (~(PECore_RunMac_PECore_RunMac_if_and_svs_st_6 | accum_vector_operator_1_for_asn_16_itm_5));
  assign mux_617_cse = MUX_s_1_2_2(mux_616_nl, or_1778_nl, while_stage_0_8);
  assign or_1776_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7
      | (~ or_tmp_915);
  assign mux_618_nl = MUX_s_1_2_2(mux_617_cse, or_1776_nl, while_stage_0_9);
  assign and_1292_cse = mux_618_nl & and_dcpl_885 & PECoreRun_wen & (accum_vector_operator_1_for_asn_10_itm_7
      | reg_PECore_RunMac_PECore_RunMac_if_and_svs_st_8_cse) & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign or_1827_nl = rva_in_PopNB_mioi_return_rsc_z_mxwt | (~(reg_rva_in_PopNB_mioi_iswt0_cse
      & (accum_vector_data_0_sva_1_load | nor_929_cse)));
  assign or_1824_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      | (~(accum_vector_data_0_sva_1_load | PECore_UpdateFSM_switch_lp_equal_tmp_3_1
      | PECore_UpdateFSM_switch_lp_equal_tmp_2_1));
  assign mux_628_nl = MUX_s_1_2_2(or_1827_nl, or_1824_nl, while_stage_0_3);
  assign or_1822_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      | (~(accum_vector_operator_1_for_asn_7_itm_1 | PECore_RunMac_PECore_RunMac_if_and_svs_st_2));
  assign mux_629_nl = MUX_s_1_2_2(mux_628_nl, or_1822_nl, while_stage_0_4);
  assign or_1820_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(input_read_req_valid_lpi_1_dfm_1_3 | PECore_RunMac_PECore_RunMac_if_and_svs_st_3));
  assign mux_630_nl = MUX_s_1_2_2(mux_629_nl, or_1820_nl, while_stage_0_5);
  assign or_1818_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | (~(accum_vector_operator_1_for_asn_7_itm_3 | reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse));
  assign mux_631_nl = MUX_s_1_2_2(mux_630_nl, or_1818_nl, while_stage_0_6);
  assign or_1816_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      | (~(PECore_RunMac_PECore_RunMac_if_and_svs_st_5 | accum_vector_operator_1_for_asn_7_itm_4));
  assign mux_632_nl = MUX_s_1_2_2(mux_631_nl, or_1816_nl, while_stage_0_7);
  assign or_1814_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6
      | (~(PECore_RunMac_PECore_RunMac_if_and_svs_st_6 | accum_vector_operator_1_for_asn_7_itm_5));
  assign mux_633_cse = MUX_s_1_2_2(mux_632_nl, or_1814_nl, while_stage_0_8);
  assign or_1812_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7
      | (~ or_tmp_949);
  assign mux_634_nl = MUX_s_1_2_2(mux_633_cse, or_1812_nl, while_stage_0_9);
  assign and_1304_cse = mux_634_nl & and_dcpl_885 & PECoreRun_wen & (accum_vector_operator_1_for_asn_1_itm_7
      | reg_PECore_RunMac_PECore_RunMac_if_and_svs_st_8_cse) & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign input_mem_banks_read_read_data_and_18_enex5 = PECoreRun_wen & and_dcpl_294
      & input_read_req_valid_lpi_1_dfm_1_6 & while_stage_0_8 & reg_input_mem_banks_read_read_data_lpi_1_dfm_1_5_31_0_enexo;
  assign weight_mem_banks_load_store_for_else_and_3_cse = PECoreRun_wen & nor_tmp_1
      & and_dcpl_40;
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_103_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm
      = MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[55:48]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_103_nl);
  assign mux_103_nl = MUX_s_1_2_2((~ or_tmp_4), or_tmp_206, crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_95_itm_1);
  assign weight_mem_banks_load_store_for_else_and_4_ssc = PECoreRun_wen & mux_103_nl
      & and_dcpl_40;
  assign weight_mem_banks_load_store_for_else_and_9_cse = PECoreRun_wen & and_dcpl_228
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_86_itm_1 & while_stage_0_6;
  assign mux_106_nl = MUX_s_1_2_2(or_tmp_4, (~ or_tmp_206), crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2]);
  assign mux_105_nl = MUX_s_1_2_2((~ or_tmp_206), or_tmp_4, crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2]);
  assign mux_107_nl = MUX_s_1_2_2(mux_106_nl, mux_105_nl, crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1]);
  assign mux_104_nl = MUX_s_1_2_2((~ or_tmp_206), or_tmp_4, or_362_cse);
  assign mux_108_nl = MUX_s_1_2_2(mux_107_nl, mux_104_nl, crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0]);
  assign weight_mem_banks_load_store_for_else_and_10_ssc = PECoreRun_wen & (~ mux_108_nl)
      & and_dcpl_40;
  assign nor_464_cse = ~((crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1:0]!=2'b00));
  assign mux_474_nl = MUX_s_1_2_2(nor_tmp, (weight_mem_write_arbxbar_xbar_for_empty_sva_2[2]),
      crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1]);
  assign or_1401_tmp = mux_474_nl | ((weight_mem_write_arbxbar_xbar_for_empty_sva_2[4])
      & nor_464_cse);
  assign or_362_cse = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2:1]!=2'b00);
  assign weight_mem_banks_load_store_for_else_and_17_cse = PECoreRun_wen & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & while_stage_0_6;
  assign nor_291_nl = ~(rva_in_reg_rw_sva_st_1_4 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_17_itm_1
      | rva_in_reg_rw_sva_st_4 | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_4 | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_4
      | rva_in_reg_rw_sva_4 | (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3) |
      PECore_DecodeAxiRead_switch_lp_nor_tmp_4);
  assign mux_118_nl = MUX_s_1_2_2((crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0]),
      (~ (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0])), crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1]);
  assign mux_119_nl = MUX_s_1_2_2(mux_118_nl, nor_464_cse, crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2]);
  assign mux_120_nl = MUX_s_1_2_2(nor_291_nl, mux_119_nl, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
  assign weight_mem_banks_load_store_for_else_and_20_ssc = PECoreRun_wen & mux_120_nl
      & and_dcpl_40;
  assign weight_mem_banks_load_store_for_else_and_22_cse = PECoreRun_wen & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_76_itm_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & while_stage_0_6;
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_78_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm
      = MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[23:16]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_78_nl);
  assign mux_121_nl = MUX_s_1_2_2((~ or_tmp_4), or_tmp_206, crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_86_itm_1);
  assign weight_mem_banks_load_store_for_else_and_27_ssc = PECoreRun_wen & mux_121_nl
      & and_dcpl_40;
  assign weight_mem_write_arbxbar_xbar_for_empty_and_enex5 = rva_in_reg_rw_and_7_cse
      & reg_weight_mem_write_arbxbar_xbar_for_empty_sva_1_enexo;
  assign and_321_cse = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]) & PECore_DecodeAxiRead_case_4_switch_lp_nor_6_tmp;
  assign ProductSum_for_and_24_cse = PECoreRun_wen & or_tmp_33 & while_stage_0_4;
  assign ProductSum_for_and_30_cse = PECoreRun_wen & PECore_RunMac_PECore_RunMac_if_and_svs_st_2
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2)
      & while_stage_0_4;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_8_cse = PECoreRun_wen & and_dcpl_293
      & (~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_4 | input_read_req_valid_lpi_1_dfm_1_6))
      & (~ rva_in_reg_rw_sva_6) & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_5 &
      while_stage_0_8;
  assign and_698_nl = accum_vector_operator_1_for_asn_7_itm_1 & not_tmp_217;
  assign mux_123_nl = MUX_s_1_2_2(PECore_RunMac_PECore_RunMac_if_and_svs_st_2, and_698_nl,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
  assign input_mem_banks_read_1_read_data_and_4_enex5 = PECoreRun_wen & mux_123_nl
      & while_stage_0_4 & reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_1_enexo;
  assign input_read_req_valid_and_2_cse = PECoreRun_wen & and_dcpl_293 & while_stage_0_8;
  assign PECore_DecodeAxiRead_switch_lp_and_11_cse = PECoreRun_wen & and_dcpl_294
      & and_dcpl_329 & while_stage_0_8;
  assign rva_out_reg_data_and_32_cse = PECoreRun_wen & and_dcpl_294 & and_dcpl_329
      & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_5 & (~(PECore_DecodeAxiRead_switch_lp_equal_tmp_3_6
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_6 | PECore_DecodeAxiRead_switch_lp_nor_tmp_6))
      & while_stage_0_8 & (~ rva_in_reg_rw_sva_st_6);
  assign rva_out_reg_data_and_91_enex5 = rva_out_reg_data_and_32_cse & reg_weight_mem_run_3_for_5_mux_12_itm_1_1_enexo;
  assign rva_out_reg_data_and_92_enex5 = rva_out_reg_data_and_32_cse & reg_weight_mem_run_3_for_5_mux_11_itm_1_1_enexo;
  assign rva_out_reg_data_and_93_enex5 = rva_out_reg_data_and_32_cse & reg_weight_mem_run_3_for_5_mux_10_itm_1_1_enexo;
  assign rva_out_reg_data_and_94_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_35_32_sva_dfm_4_1_enexo;
  assign rva_out_reg_data_and_95_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_62_56_sva_dfm_4_1_enexo;
  assign PECore_RunScale_if_and_3_cse = PECoreRun_wen & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6)
      & while_stage_0_8;
  assign and_1320_cse = mux_537_cse & and_dcpl_964 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7)
      & or_tmp_745 & PECoreRun_wen;
  assign and_1332_cse = mux_545_cse & and_dcpl_964 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7)
      & or_tmp_762 & PECoreRun_wen;
  assign and_1344_cse = mux_553_cse & and_dcpl_964 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7)
      & or_tmp_779 & PECoreRun_wen;
  assign and_1356_cse = mux_561_cse & and_dcpl_964 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7)
      & or_tmp_796 & PECoreRun_wen;
  assign and_1368_cse = mux_577_cse & and_dcpl_964 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7)
      & or_tmp_830 & PECoreRun_wen;
  assign and_1380_cse = mux_617_cse & and_dcpl_964 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7)
      & or_tmp_915 & PECoreRun_wen;
  assign and_1392_cse = mux_633_cse & and_dcpl_964 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7)
      & or_tmp_949 & PECoreRun_wen;
  assign PECore_RunMac_if_and_5_cse = PECoreRun_wen & and_dcpl_204;
  assign ProductSum_for_and_32_cse = PECoreRun_wen & while_and_4_cse;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_12_cse = PECoreRun_wen & while_and_23_cse
      & while_stage_0_7 & (~ rva_in_reg_rw_sva_st_1_5) & (~(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_11_itm_1
      | rva_in_reg_rw_sva_5)) & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4;
  assign nor_353_nl = ~((~ ProductSum_for_asn_64_itm_1) | reg_rva_in_reg_rw_sva_st_1_1_cse);
  assign mux_173_nl = MUX_s_1_2_2(PECore_UpdateFSM_switch_lp_equal_tmp_3_1, nor_353_nl,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign input_mem_banks_read_1_read_data_and_5_enex5 = PECoreRun_wen & mux_173_nl
      & while_stage_0_3 & (reg_input_mem_banks_bank_a_56_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_229_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_160_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_92_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_100_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_43_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_118_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_201_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_99_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_4_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_230_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_128_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_191_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_40_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_244_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_219_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_106_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_120_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_52_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_16_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_149_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_142_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_104_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_170_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_23_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_222_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_147_sva_dfm_2_enexo | reg_input_read_addrs_sva_1_1_enexo
      | reg_input_mem_banks_bank_a_156_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_113_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_32_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_196_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_44_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_175_sva_dfm_2_enexo
      | reg_input_mem_banks_read_read_data_sva_1_enexo | reg_input_mem_banks_bank_a_6_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_83_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_19_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_197_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_181_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_254_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_95_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_105_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_242_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_28_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_218_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_236_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_24_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_88_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_210_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_3_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_178_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_68_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_162_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_192_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_233_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_37_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_125_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_203_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_111_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_55_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_112_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_208_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_146_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_85_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_78_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_221_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_194_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_186_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_150_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_70_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_79_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_110_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_71_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_108_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_90_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_212_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_202_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_198_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_60_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_15_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_93_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_5_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_165_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_58_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_187_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_42_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_47_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_190_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_225_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_158_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_80_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_129_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_234_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_65_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_45_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_207_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_2_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_167_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_89_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_238_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_217_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_204_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_74_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_127_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_220_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_166_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_164_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_54_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_139_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_98_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_25_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_0_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_53_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_141_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_29_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_86_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_14_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_248_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_67_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_184_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_82_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_143_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_240_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_136_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_61_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_109_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_228_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_63_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_241_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_26_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_34_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_94_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_159_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_62_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_30_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_144_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_209_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_215_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_51_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_119_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_173_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_8_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_12_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_116_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_132_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_35_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_84_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_134_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_18_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_11_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_39_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_124_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_224_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_161_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_235_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_73_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_232_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_239_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_253_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_205_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_133_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_223_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_249_sva_dfm_2_enexo
      | reg_input_write_req_valid_lpi_1_dfm_1_1_enexo | reg_input_mem_banks_bank_a_75_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_251_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_20_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_182_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_153_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_172_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_176_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_252_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_185_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_211_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_57_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_123_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_66_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_231_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_126_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_81_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_1_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_206_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_237_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_64_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_213_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_97_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_36_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_155_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_107_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_130_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_189_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_115_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_49_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_245_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_114_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_169_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_17_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_22_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_9_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_87_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_59_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_180_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_200_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_255_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_195_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_246_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_27_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_21_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_157_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_168_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_243_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_131_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_214_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_33_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_77_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_174_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_193_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_38_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_216_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_151_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_152_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_171_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_163_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_227_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_103_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_69_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_117_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_140_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_122_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_91_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_135_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_96_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_50_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_148_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_48_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_179_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_7_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_10_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_31_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_145_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_199_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_226_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_102_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_72_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_247_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_76_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_46_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_250_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_101_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_137_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_121_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_188_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_13_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_138_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_154_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_41_sva_dfm_2_enexo | reg_input_mem_banks_bank_a_183_sva_dfm_2_enexo
      | reg_input_mem_banks_bank_a_177_sva_dfm_2_enexo);
  assign input_mem_banks_read_read_data_and_19_enex5 = PECoreRun_wen & and_dcpl_355
      & (~ rva_in_reg_rw_sva_st_1_5) & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_11_itm_1
      & reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo;
  assign input_read_req_valid_and_3_cse = PECoreRun_wen & and_dcpl_241 & (~ rva_in_reg_rw_sva_st_1_5);
  assign PECore_DecodeAxiRead_switch_lp_and_15_cse = PECoreRun_wen & and_dcpl_355
      & (~(rva_in_reg_rw_sva_st_1_5 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_11_itm_1
      | rva_in_reg_rw_sva_5));
  assign rva_out_reg_data_and_40_cse = PECoreRun_wen & and_dcpl_241 & (~(rva_in_reg_rw_sva_st_1_5
      & rva_in_reg_rw_sva_5));
  assign and_1402_cse = (~(((~((~ while_stage_0_8) | rva_in_reg_rw_sva_6 | (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6)
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_11_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3)) | rva_in_reg_rw_sva_st_1_5)
      & rva_in_reg_rw_sva_5)) & weight_mem_run_3_for_aelse_and_cse & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
  assign PECore_RunScale_if_and_5_cse = PECoreRun_wen & and_dcpl_32;
  assign rva_out_reg_data_and_45_cse = weight_mem_read_arbxbar_arbiters_next_and_cse
      & (nand_27_cse | rva_in_reg_rw_sva_5);
  assign and_1411_cse = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6
      & (~ rva_in_reg_rw_sva_6) & while_stage_0_8 & fsm_output & (rva_in_reg_rw_sva_5
      | (~ while_stage_0_7) | (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5))
      & PECoreRun_wen;
  assign nor_469_cse = ~(weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign or_2088_cse = state_0_sva | (state_2_1_sva[1]);
  assign nor_963_nl = ~((state_2_1_sva[0]) | (~ input_port_PopNB_mioi_return_rsc_z_mxwt));
  assign mux_743_cse = MUX_s_1_2_2(nor_963_nl, PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva,
      or_2088_cse);
  assign nand_407_cse = ~((while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[1:0]==2'b11));
  assign nand_408_cse = ~((while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2:0]==3'b111));
  assign nand_410_cse = ~((while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3:0]==4'b1111));
  assign nor_1000_nl = ~((state_2_1_sva[0]) | (~ input_port_PopNB_mioi_return_rsc_z_mxwt)
      | PECore_RunFSM_switch_lp_nor_tmp_1);
  assign nor_1001_nl = ~((~ PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva)
      | PECore_RunFSM_switch_lp_nor_tmp_1);
  assign mux_773_cse = MUX_s_1_2_2(nor_1000_nl, nor_1001_nl, or_2088_cse);
  assign or_2278_nl = (state_2_1_sva[0]) | (~ input_port_PopNB_mioi_return_rsc_z_mxwt)
      | PECore_RunFSM_switch_lp_nor_tmp_1 | (~ (PEManager_15U_GetInputAddr_acc_tmp[0]));
  assign or_2276_nl = (~ PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva)
      | PECore_RunFSM_switch_lp_nor_tmp_1 | (~ (PEManager_15U_GetInputAddr_acc_tmp[0]));
  assign mux_799_cse = MUX_s_1_2_2(or_2278_nl, or_2276_nl, or_2088_cse);
  assign nand_414_cse = ~((while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4:0]==5'b11111));
  assign nand_422_cse = ~((while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5:0]==6'b111111));
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_16_cse = PECoreRun_wen & (~ or_tmp_4)
      & and_dcpl_40 & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3;
  assign mux_176_nl = MUX_s_1_2_2(weight_mem_run_3_for_land_4_lpi_1_dfm_1, (~ or_tmp_4),
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign PECore_DecodeAxiRead_switch_lp_and_19_cse = PECoreRun_wen & mux_176_nl &
      while_stage_0_6;
  assign or_1095_nl = (~ (state_2_1_sva[0])) | state_0_sva | (state_2_1_sva[1]) |
      (~ reg_rva_in_PopNB_mioi_iswt0_cse) | rva_in_PopNB_mioi_return_rsc_z_mxwt;
  assign and_649_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & (state_0_sva | (state_2_1_sva_dfm_1[1]) | (~ reg_rva_in_PopNB_mioi_iswt0_cse)
      | rva_in_PopNB_mioi_return_rsc_z_mxwt);
  assign mux_277_nl = MUX_s_1_2_2(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1,
      and_649_nl, state_2_1_sva_dfm_1[0]);
  assign mux_278_nl = MUX_s_1_2_2(or_1095_nl, mux_277_nl, while_stage_0_3);
  assign and_680_cse = PECoreRun_wen & (~ mux_278_nl);
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_19_cse = PECoreRun_wen & and_dcpl_376
      & (~(input_read_req_valid_lpi_1_dfm_1_3 | rva_in_reg_rw_sva_3)) & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_2
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      & while_stage_0_5;
  assign and_700_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1 & Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_1;
  assign and_703_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1 & Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_5;
  assign and_702_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1 & reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_5_cse;
  assign mux_185_nl = MUX_s_1_2_2(weight_mem_run_3_for_land_1_lpi_1_dfm_1, (~ or_tmp_334),
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign PECore_DecodeAxiRead_switch_lp_and_23_cse = PECoreRun_wen & mux_185_nl &
      while_stage_0_5;
  assign rva_out_reg_data_and_51_cse = PECoreRun_wen & and_dcpl_389 & (~(rva_in_reg_rw_sva_3
      | PECore_DecodeAxiRead_switch_lp_nor_tmp_3)) & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_2
      & (~(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_3 | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_3
      | rva_in_reg_rw_sva_st_3)) & and_dcpl_69;
  assign rva_out_reg_data_and_96_enex5 = rva_out_reg_data_and_51_cse & reg_rva_out_reg_data_30_25_sva_dfm_1_enexo;
  assign rva_out_reg_data_and_97_enex5 = rva_out_reg_data_and_51_cse & reg_rva_out_reg_data_23_17_sva_dfm_1_enexo;
  assign rva_out_reg_data_and_98_enex5 = rva_out_reg_data_and_51_cse & reg_rva_out_reg_data_15_9_sva_dfm_3_enexo;
  assign rva_out_reg_data_and_54_cse = PECoreRun_wen & and_dcpl_389 & (~ rva_in_reg_rw_sva_3)
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      & while_stage_0_5;
  assign rva_out_reg_data_and_99_enex5 = rva_out_reg_data_and_54_cse & reg_rva_out_reg_data_35_32_sva_dfm_1_3_enexo;
  assign rva_out_reg_data_and_100_enex5 = rva_out_reg_data_and_54_cse & reg_rva_out_reg_data_39_36_sva_dfm_1_3_enexo;
  assign rva_out_reg_data_and_101_enex5 = rva_out_reg_data_and_54_cse & reg_rva_out_reg_data_46_40_sva_dfm_1_3_enexo;
  assign rva_out_reg_data_and_102_enex5 = rva_out_reg_data_and_54_cse & reg_rva_out_reg_data_62_56_sva_dfm_1_3_enexo;
  assign rva_out_reg_data_and_103_enex5 = rva_out_reg_data_and_54_cse & reg_rva_out_reg_data_55_48_sva_dfm_1_3_enexo;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_24_cse = PECoreRun_wen & and_dcpl_401
      & and_dcpl_398 & while_stage_0_4 & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_1;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_25_cse = PECoreRun_wen & and_dcpl_401
      & and_dcpl_398 & while_stage_0_4;
  assign PECore_DecodeAxiRead_switch_lp_and_27_cse = PECoreRun_wen & (~((~(not_tmp_217
      & nor_320_cse)) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2))
      & while_stage_0_4;
  assign rva_out_reg_data_and_59_cse = PECoreRun_wen & not_tmp_217 & nor_320_cse
      & (~ PECore_DecodeAxiRead_switch_lp_nor_tmp_2) & (~(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_2)) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4 & PECore_DecodeAxiRead_switch_lp_equal_tmp_1_1;
  assign rva_out_reg_data_and_104_enex5 = rva_out_reg_data_and_59_cse & reg_rva_out_reg_data_15_9_sva_dfm_2_enexo;
  assign rva_out_reg_data_and_105_enex5 = PECore_DecodeAxiRead_case_4_switch_lp_and_25_cse
      & reg_rva_out_reg_data_35_32_sva_dfm_1_2_enexo;
  assign rva_out_reg_data_and_106_enex5 = PECore_DecodeAxiRead_case_4_switch_lp_and_25_cse
      & reg_rva_out_reg_data_39_36_sva_dfm_1_2_enexo;
  assign rva_out_reg_data_and_107_enex5 = PECore_DecodeAxiRead_case_4_switch_lp_and_25_cse
      & reg_rva_out_reg_data_46_40_sva_dfm_1_2_enexo;
  assign rva_out_reg_data_and_108_enex5 = PECore_DecodeAxiRead_case_4_switch_lp_and_25_cse
      & reg_rva_out_reg_data_62_56_sva_dfm_1_2_enexo;
  assign rva_out_reg_data_and_109_enex5 = PECore_DecodeAxiRead_case_4_switch_lp_and_25_cse
      & reg_rva_out_reg_data_55_48_sva_dfm_1_2_enexo;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_29_cse = PECoreRun_wen & mux_tmp_182
      & and_dcpl_420;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_30_cse = PECoreRun_wen & and_dcpl_420;
  assign PECore_DecodeAxiRead_switch_lp_and_31_cse = PECoreRun_wen & (and_dcpl_419
      | (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      & while_stage_0_3;
  assign rva_out_reg_data_and_67_enex5 = PECoreRun_wen & and_dcpl_431 & (while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1[3:1]==3'b010)
      & (~(reg_rva_in_reg_rw_sva_st_1_1_cse | PECore_DecodeAxiRead_switch_lp_nor_tmp_1
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_3)) & (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_2)
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3 & reg_rva_out_reg_data_15_9_sva_dfm_1_enexo;
  assign rva_out_reg_data_and_110_enex5 = PECore_DecodeAxiRead_case_4_switch_lp_and_30_cse
      & reg_rva_out_reg_data_35_32_sva_dfm_1_1_enexo;
  assign rva_out_reg_data_and_111_enex5 = PECore_DecodeAxiRead_case_4_switch_lp_and_30_cse
      & reg_rva_out_reg_data_39_36_sva_dfm_1_1_enexo;
  assign rva_out_reg_data_and_112_enex5 = PECore_DecodeAxiRead_case_4_switch_lp_and_30_cse
      & reg_rva_out_reg_data_46_40_sva_dfm_1_1_enexo;
  assign rva_out_reg_data_and_113_enex5 = PECore_DecodeAxiRead_case_4_switch_lp_and_30_cse
      & reg_rva_out_reg_data_62_56_sva_dfm_1_1_enexo;
  assign rva_out_reg_data_and_114_enex5 = PECore_DecodeAxiRead_case_4_switch_lp_and_30_cse
      & reg_pe_config_input_counter_sva_dfm_1_enexo;
  assign PECore_DecodeAxiRead_switch_lp_nor_2_cse = ~((while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1[3])
      | (while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1[1])
      | (while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1[0]));
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_33_cse = PECoreRun_wen & (~((~(mux_tmp_182
      & and_dcpl_419)) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      & while_stage_0_3;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_34_cse = PECoreRun_wen & mux_tmp_182
      & and_dcpl_419 & (~ PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_1) &
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_37_cse = PECoreRun_wen & and_dcpl_215
      & and_dcpl_217 & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]));
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_39_cse = PECoreRun_wen & and_dcpl_312
      & (~(rva_in_PopNB_mioi_data_rw_rsc_z_mxwt | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])))
      & nand_36_cse;
  assign PECore_DecodeAxiRead_case_4_switch_lp_and_41_cse = PECoreRun_wen & (or_dcpl_91
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17:16]!=2'b10)) & and_dcpl_242;
  assign nor_17_cse = ~(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_itm_1
      | (~ reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_2_1_itm_2_cse));
  assign nor_18_cse = ~(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_20_itm_1
      | (~ reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse));
  assign and_516_cse = while_stage_0_11 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_9
      & (~ rva_in_reg_rw_sva_st_1_9);
  assign or_999_cse = (state_2_1_sva!=2'b00) | state_0_sva;
  assign weight_mem_run_3_for_5_and_161_cse = reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_20_itm_2_cse
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_175_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_54_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_176_cse = reg_weight_mem_run_3_for_5_and_163_itm_2_cse
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_177_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_56_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_178_cse = reg_weight_mem_run_3_for_5_and_165_itm_2_cse
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_180_cse = reg_weight_mem_run_3_for_5_and_167_itm_2_cse
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_181_cse = reg_weight_mem_run_3_for_5_and_168_itm_2_cse
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_port_read_out_data_5_0_sva_dfm_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[7:0]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[7:0]),
      BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9, weight_port_read_out_data_5_0_sva_dfm_1,
      {weight_mem_run_3_for_5_and_172 , weight_mem_run_3_for_5_asn_315 , weight_mem_run_3_for_5_asn_317
      , weight_mem_run_3_for_5_and_44_itm_2 , weight_mem_run_3_for_5_asn_319 , weight_mem_run_3_for_5_and_38_itm_1
      , weight_mem_run_3_for_5_and_39_itm_2 , weight_mem_run_3_for_5_and_48_itm_1
      , (~ weight_mem_run_3_for_land_6_lpi_1_dfm_2)});
  assign weight_port_read_out_data_5_1_sva_dfm_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:8]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:8]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[7:0]), weight_port_read_out_data_5_1_sva_dfm_1,
      {weight_mem_run_3_for_5_and_172 , weight_mem_run_3_for_5_asn_315 , weight_mem_run_3_for_5_asn_317
      , weight_mem_run_3_for_5_and_44_itm_2 , weight_mem_run_3_for_5_asn_319 , weight_mem_run_3_for_5_and_46_itm_2
      , weight_mem_run_3_for_5_and_47_itm_1 , weight_mem_run_3_for_5_and_48_itm_1
      , (~ weight_mem_run_3_for_land_6_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_0_sva_dfm_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[7:0]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[7:0]),
      BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9, weight_port_read_out_data_7_0_sva_dfm_1,
      {weight_mem_run_3_for_5_and_168 , weight_mem_run_3_for_5_asn_309 , weight_mem_run_3_for_5_asn_311
      , weight_mem_run_3_for_5_and_108_itm_1 , weight_mem_run_3_for_5_asn_313 , weight_mem_run_3_for_5_and_102_itm_2
      , weight_mem_run_3_for_5_and_103_itm_2 , weight_mem_run_3_for_5_and_112_itm_1
      , (~ weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_1_sva_dfm_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:8]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:8]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[7:0]), weight_port_read_out_data_7_1_sva_dfm_1,
      {weight_mem_run_3_for_5_and_174 , weight_mem_run_3_for_5_asn_309 , weight_mem_run_3_for_5_asn_311
      , weight_mem_run_3_for_5_and_108_itm_1 , weight_mem_run_3_for_5_asn_313 , weight_mem_run_3_for_5_and_110_itm_1
      , weight_mem_run_3_for_5_and_111_itm_1 , weight_mem_run_3_for_5_and_112_itm_1
      , (~ weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_3_sva_dfm_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:24]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31:24]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[23:16]), weight_port_read_out_data_7_3_sva_dfm_1_1,
      {weight_mem_run_3_for_5_and_174 , weight_mem_run_3_for_5_asn_309 , weight_mem_run_3_for_5_asn_311
      , weight_mem_run_3_for_5_and_156_itm_2 , weight_mem_run_3_for_5_asn_313 , weight_mem_run_3_for_5_and_102_itm_2
      , weight_mem_run_3_for_5_and_111_itm_1 , weight_mem_run_3_for_5_and_112_itm_1
      , (~ weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_2_sva_dfm_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[23:16]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[23:16]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[15:8]), weight_port_read_out_data_7_2_sva_dfm_1_1,
      {weight_mem_run_3_for_5_and_168 , weight_mem_run_3_for_5_asn_309 , weight_mem_run_3_for_5_asn_311
      , weight_mem_run_3_for_5_and_108_itm_1 , weight_mem_run_3_for_5_asn_313 , weight_mem_run_3_for_5_and_102_itm_2
      , weight_mem_run_3_for_5_and_111_itm_1 , weight_mem_run_3_for_5_and_112_itm_1
      , (~ weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_5_sva_dfm_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:40]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:40]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[39:32]), weight_port_read_out_data_7_5_sva_dfm_1_1,
      {weight_mem_run_3_for_5_and_174 , weight_mem_run_3_for_5_asn_309 , weight_mem_run_3_for_5_asn_311
      , weight_mem_run_3_for_5_and_156_itm_2 , weight_mem_run_3_for_5_asn_313 , weight_mem_run_3_for_5_and_102_itm_2
      , weight_mem_run_3_for_5_and_111_itm_1 , weight_mem_run_3_for_5_and_112_itm_1
      , (~ weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_4_sva_dfm_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[39:32]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[39:32]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[31:24]), weight_port_read_out_data_7_4_sva_dfm_1_1,
      {weight_mem_run_3_for_5_and_168 , weight_mem_run_3_for_5_asn_309 , weight_mem_run_3_for_5_asn_311
      , weight_mem_run_3_for_5_and_108_itm_1 , weight_mem_run_3_for_5_asn_313 , weight_mem_run_3_for_5_and_102_itm_2
      , weight_mem_run_3_for_5_and_111_itm_1 , weight_mem_run_3_for_5_asn_321 , (~
      weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_7_sva_dfm_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:56]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:56]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[55:48]), weight_port_read_out_data_7_7_sva_dfm_1_1,
      {weight_mem_run_3_for_5_and_168 , weight_mem_run_3_for_5_asn_309 , weight_mem_run_3_for_5_asn_311
      , weight_mem_run_3_for_5_and_156_itm_2 , weight_mem_run_3_for_5_asn_313 , weight_mem_run_3_for_5_and_110_itm_1
      , weight_mem_run_3_for_5_and_111_itm_1 , weight_mem_run_3_for_5_asn_321 , (~
      weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_7_6_sva_dfm_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[55:48]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[55:48]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[47:40]), weight_port_read_out_data_7_6_sva_dfm_1_1,
      {weight_mem_run_3_for_5_and_168 , weight_mem_run_3_for_5_asn_309 , weight_mem_run_3_for_5_asn_311
      , weight_mem_run_3_for_5_and_156_itm_2 , weight_mem_run_3_for_5_asn_313 , weight_mem_run_3_for_5_and_102_itm_2
      , weight_mem_run_3_for_5_and_111_itm_1 , weight_mem_run_3_for_5_asn_321 , (~
      weight_mem_run_3_for_land_lpi_1_dfm_2)});
  assign weight_port_read_out_data_5_3_sva_dfm_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:24]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31:24]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[23:16]), weight_port_read_out_data_5_3_sva_dfm_1_1,
      {weight_mem_run_3_for_5_and_172 , weight_mem_run_3_for_5_asn_315 , weight_mem_run_3_for_5_asn_317
      , weight_mem_run_3_for_5_and_44_itm_2 , weight_mem_run_3_for_5_asn_319 , weight_mem_run_3_for_5_and_38_itm_1
      , weight_mem_run_3_for_5_and_47_itm_1 , weight_mem_run_3_for_5_and_48_itm_1
      , (~ weight_mem_run_3_for_land_6_lpi_1_dfm_2)});
  assign weight_port_read_out_data_5_2_sva_dfm_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[23:16]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[23:16]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[15:8]), weight_port_read_out_data_5_2_sva_dfm_1_1,
      {weight_mem_run_3_for_5_and_172 , weight_mem_run_3_for_5_asn_315 , weight_mem_run_3_for_5_asn_317
      , weight_mem_run_3_for_5_and_44_itm_2 , weight_mem_run_3_for_5_asn_319 , weight_mem_run_3_for_5_and_46_itm_2
      , weight_mem_run_3_for_5_and_39_itm_2 , weight_mem_run_3_for_5_asn_323 , (~
      weight_mem_run_3_for_land_6_lpi_1_dfm_2)});
  assign weight_port_read_out_data_5_5_sva_dfm_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:40]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:40]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[39:32]), weight_port_read_out_data_5_5_sva_dfm_1_1,
      {weight_mem_run_3_for_5_and_172 , weight_mem_run_3_for_5_asn_315 , weight_mem_run_3_for_5_asn_317
      , weight_mem_run_3_for_5_and_44_itm_2 , weight_mem_run_3_for_5_asn_319 , weight_mem_run_3_for_5_and_38_itm_1
      , weight_mem_run_3_for_5_and_47_itm_1 , weight_mem_run_3_for_5_and_48_itm_1
      , (~ weight_mem_run_3_for_land_6_lpi_1_dfm_2)});
  assign weight_port_read_out_data_5_4_sva_dfm_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[39:32]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[39:32]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[31:24]), weight_port_read_out_data_5_4_sva_dfm_1_1,
      {weight_mem_run_3_for_5_and_172 , weight_mem_run_3_for_5_asn_315 , weight_mem_run_3_for_5_asn_317
      , weight_mem_run_3_for_5_and_44_itm_2 , weight_mem_run_3_for_5_asn_319 , weight_mem_run_3_for_5_and_46_itm_2
      , weight_mem_run_3_for_5_and_39_itm_2 , weight_mem_run_3_for_5_asn_323 , (~
      weight_mem_run_3_for_land_6_lpi_1_dfm_2)});
  assign weight_port_read_out_data_5_7_sva_dfm_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:56]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:56]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[55:48]), weight_port_read_out_data_5_7_sva_dfm_1_1,
      {weight_mem_run_3_for_5_and_172 , weight_mem_run_3_for_5_asn_315 , weight_mem_run_3_for_5_asn_317
      , weight_mem_run_3_for_5_and_44_itm_2 , weight_mem_run_3_for_5_asn_319 , weight_mem_run_3_for_5_and_38_itm_1
      , weight_mem_run_3_for_5_and_39_itm_2 , weight_mem_run_3_for_5_and_48_itm_1
      , (~ weight_mem_run_3_for_land_6_lpi_1_dfm_2)});
  assign weight_mem_run_3_for_5_and_81_nl = weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_10_itm_1
      & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign weight_port_read_out_data_5_6_sva_dfm_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[55:48]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[55:48]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[47:40]), weight_port_read_out_data_5_6_sva_dfm_1_1,
      {weight_mem_run_3_for_5_and_81_nl , weight_mem_run_3_for_5_asn_315 , weight_mem_run_3_for_5_asn_317
      , weight_mem_run_3_for_5_and_84_itm_1 , weight_mem_run_3_for_5_asn_319 , weight_mem_run_3_for_5_and_46_itm_2
      , weight_mem_run_3_for_5_and_39_itm_2 , weight_mem_run_3_for_5_asn_323 , (~
      weight_mem_run_3_for_land_6_lpi_1_dfm_2)});
  assign weight_port_read_out_data_3_5_sva_dfm_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:40]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:40]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[39:32]), weight_port_read_out_data_3_5_sva_dfm_1_1,
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_65_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_118
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_120 , weight_mem_run_3_for_5_and_20_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_122 , weight_mem_run_3_for_5_and_30_itm_2
      , weight_mem_run_3_for_5_and_31_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_124
      , (~ weight_mem_run_3_for_land_4_lpi_1_dfm_2)});
  assign weight_mem_run_3_for_5_and_7_nl = (weight_read_addrs_3_lpi_1_dfm_3_2_0==3'b110)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign weight_port_read_out_data_3_4_sva_dfm_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[39:32]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[39:32]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[31:24]), weight_port_read_out_data_3_4_sva_dfm_1_1,
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_65_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_118
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_120 , weight_mem_run_3_for_5_and_20_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_122 , weight_mem_run_3_for_5_and_30_itm_2
      , weight_mem_run_3_for_5_and_7_nl , weight_mem_run_3_for_5_and_8_itm_1 , (~
      weight_mem_run_3_for_land_4_lpi_1_dfm_2)});
  assign weight_port_read_out_data_3_7_sva_dfm_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:56]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:56]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[55:48]), weight_port_read_out_data_3_7_sva_dfm_1_1,
      {weight_mem_run_3_for_5_and_166 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_118
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_120 , weight_mem_run_3_for_5_and_28_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_122 , weight_mem_run_3_for_5_and_30_itm_2
      , weight_mem_run_3_for_5_and_31_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_124
      , (~ weight_mem_run_3_for_land_4_lpi_1_dfm_2)});
  assign weight_port_read_out_data_3_6_sva_dfm_2 = MUX1HOT_v_8_9_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[55:48]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[55:48]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[47:40]), weight_port_read_out_data_3_6_sva_dfm_1_1,
      {weight_mem_run_3_for_5_and_166 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_118
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_120 , weight_mem_run_3_for_5_and_20_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_122 , weight_mem_run_3_for_5_and_22_itm_1
      , weight_mem_run_3_for_5_and_23_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_124
      , (~ weight_mem_run_3_for_land_4_lpi_1_dfm_2)});
  assign PECore_PushAxiRsp_if_else_mux_13_mx0w2 = MUX_s_1_2_2(rva_out_reg_data_63_sva_dfm_7,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[63]), crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_11_itm_1);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_10_itm_mx0w0
      = ~((weight_read_addrs_3_lpi_1_dfm_2_2_0!=3'b000));
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_tmp
      = ~((crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2!=3'b000));
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_84_itm_mx0w0 = (weight_read_addrs_3_lpi_1_dfm_2_2_0==3'b011)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_1;
  assign Arbiter_8U_Roundrobin_pick_nand_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1)
      & and_dcpl_78)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_40_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1
      & and_dcpl_78;
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_56_nl = weight_mem_read_arbxbar_arbiters_next_7_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign weight_mem_read_arbxbar_arbiters_next_7_1_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_56_nl,
      weight_mem_read_arbxbar_arbiters_next_7_1_sva, Arbiter_8U_Roundrobin_pick_1_mux_542_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_nand_cse , Arbiter_8U_Roundrobin_pick_and_40_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_57_nl = weight_mem_read_arbxbar_arbiters_next_7_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign weight_mem_read_arbxbar_arbiters_next_7_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_57_nl,
      weight_mem_read_arbxbar_arbiters_next_7_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_541_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_nand_cse , Arbiter_8U_Roundrobin_pick_and_40_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_58_nl = weight_mem_read_arbxbar_arbiters_next_7_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign weight_mem_read_arbxbar_arbiters_next_7_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_58_nl,
      weight_mem_read_arbxbar_arbiters_next_7_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_540_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_nand_cse , Arbiter_8U_Roundrobin_pick_and_40_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_59_nl = weight_mem_read_arbxbar_arbiters_next_7_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign weight_mem_read_arbxbar_arbiters_next_7_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_59_nl,
      weight_mem_read_arbxbar_arbiters_next_7_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_539_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_nand_cse , Arbiter_8U_Roundrobin_pick_and_40_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_60_nl = weight_mem_read_arbxbar_arbiters_next_7_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign weight_mem_read_arbxbar_arbiters_next_7_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_60_nl,
      weight_mem_read_arbxbar_arbiters_next_7_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_538_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_nand_cse , Arbiter_8U_Roundrobin_pick_and_40_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_61_nl = weight_mem_read_arbxbar_arbiters_next_7_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign weight_mem_read_arbxbar_arbiters_next_7_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_61_nl,
      weight_mem_read_arbxbar_arbiters_next_7_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_537_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_nand_cse , Arbiter_8U_Roundrobin_pick_and_40_cse});
  assign weight_mem_read_arbxbar_arbiters_next_7_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_576_itm_1, and_dcpl_78);
  assign Arbiter_8U_Roundrobin_pick_nand_69_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1)
      & and_dcpl_78)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_52_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1
      & and_dcpl_78;
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_62_nl = weight_mem_read_arbxbar_arbiters_next_6_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[6]);
  assign weight_mem_read_arbxbar_arbiters_next_6_1_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_62_nl,
      weight_mem_read_arbxbar_arbiters_next_6_1_sva, Arbiter_8U_Roundrobin_pick_1_mux_469_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_nand_69_cse , Arbiter_8U_Roundrobin_pick_and_52_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_63_nl = weight_mem_read_arbxbar_arbiters_next_6_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[6]);
  assign weight_mem_read_arbxbar_arbiters_next_6_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_63_nl,
      weight_mem_read_arbxbar_arbiters_next_6_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_468_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_nand_69_cse , Arbiter_8U_Roundrobin_pick_and_52_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_64_nl = weight_mem_read_arbxbar_arbiters_next_6_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[6]);
  assign weight_mem_read_arbxbar_arbiters_next_6_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_64_nl,
      weight_mem_read_arbxbar_arbiters_next_6_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_467_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_nand_69_cse , Arbiter_8U_Roundrobin_pick_and_52_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_65_nl = weight_mem_read_arbxbar_arbiters_next_6_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[6]);
  assign weight_mem_read_arbxbar_arbiters_next_6_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_65_nl,
      weight_mem_read_arbxbar_arbiters_next_6_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_466_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_nand_69_cse , Arbiter_8U_Roundrobin_pick_and_52_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_66_nl = weight_mem_read_arbxbar_arbiters_next_6_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[6]);
  assign weight_mem_read_arbxbar_arbiters_next_6_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_66_nl,
      weight_mem_read_arbxbar_arbiters_next_6_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_465_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_nand_69_cse , Arbiter_8U_Roundrobin_pick_and_52_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_67_nl = weight_mem_read_arbxbar_arbiters_next_6_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[6]);
  assign weight_mem_read_arbxbar_arbiters_next_6_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_67_nl,
      weight_mem_read_arbxbar_arbiters_next_6_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_464_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_nand_69_cse , Arbiter_8U_Roundrobin_pick_and_52_cse});
  assign weight_mem_read_arbxbar_arbiters_next_6_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_496_itm_1, and_dcpl_78);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_41_mx1w0 = weight_mem_read_arbxbar_arbiters_next_5_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[5]);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_nand_cse = ~((~((~
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1) & and_dcpl_78)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_1_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1
      & and_dcpl_78;
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_69_nl = weight_mem_read_arbxbar_arbiters_next_5_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[5]);
  assign weight_mem_read_arbxbar_arbiters_next_5_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_69_nl,
      weight_mem_read_arbxbar_arbiters_next_5_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_395_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_nand_cse
      , Arbiter_8U_Roundrobin_pick_and_1_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_70_nl = weight_mem_read_arbxbar_arbiters_next_5_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[5]);
  assign weight_mem_read_arbxbar_arbiters_next_5_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_70_nl,
      weight_mem_read_arbxbar_arbiters_next_5_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_394_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_nand_cse
      , Arbiter_8U_Roundrobin_pick_and_1_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_71_nl = weight_mem_read_arbxbar_arbiters_next_5_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[5]);
  assign weight_mem_read_arbxbar_arbiters_next_5_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_71_nl,
      weight_mem_read_arbxbar_arbiters_next_5_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_393_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_nand_cse
      , Arbiter_8U_Roundrobin_pick_and_1_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_72_nl = weight_mem_read_arbxbar_arbiters_next_5_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[5]);
  assign weight_mem_read_arbxbar_arbiters_next_5_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_72_nl,
      weight_mem_read_arbxbar_arbiters_next_5_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_392_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_nand_cse
      , Arbiter_8U_Roundrobin_pick_and_1_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_36_mx1w0 = weight_mem_read_arbxbar_arbiters_next_5_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[5]);
  assign weight_mem_read_arbxbar_arbiters_next_5_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_36_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_5_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_391_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_nand_cse
      , Arbiter_8U_Roundrobin_pick_and_1_cse});
  assign weight_mem_read_arbxbar_arbiters_next_5_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_423_itm_1, and_dcpl_78);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_34_mx1w0 = weight_mem_read_arbxbar_arbiters_next_4_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[4]);
  assign Arbiter_8U_Roundrobin_pick_nand_54_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1)
      & and_dcpl_78)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_37_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1
      & and_dcpl_78;
  assign weight_mem_read_arbxbar_arbiters_next_4_1_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_34_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_4_1_sva, Arbiter_8U_Roundrobin_pick_1_mux_323_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_nand_54_cse , Arbiter_8U_Roundrobin_pick_and_37_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_33_mx1w0 = weight_mem_read_arbxbar_arbiters_next_4_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[4]);
  assign weight_mem_read_arbxbar_arbiters_next_4_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_33_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_4_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_322_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_nand_54_cse , Arbiter_8U_Roundrobin_pick_and_37_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_32_mx1w0 = weight_mem_read_arbxbar_arbiters_next_4_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[4]);
  assign weight_mem_read_arbxbar_arbiters_next_4_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_32_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_4_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_321_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_nand_54_cse , Arbiter_8U_Roundrobin_pick_and_37_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_31_mx1w0 = weight_mem_read_arbxbar_arbiters_next_4_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[4]);
  assign weight_mem_read_arbxbar_arbiters_next_4_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_31_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_4_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_320_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_nand_54_cse , Arbiter_8U_Roundrobin_pick_and_37_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_30_mx1w0 = weight_mem_read_arbxbar_arbiters_next_4_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[4]);
  assign weight_mem_read_arbxbar_arbiters_next_4_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_30_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_4_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_319_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_nand_54_cse , Arbiter_8U_Roundrobin_pick_and_37_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_29_mx1w0 = weight_mem_read_arbxbar_arbiters_next_4_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[4]);
  assign weight_mem_read_arbxbar_arbiters_next_4_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_29_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_4_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_318_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_nand_54_cse , Arbiter_8U_Roundrobin_pick_and_37_cse});
  assign weight_mem_read_arbxbar_arbiters_next_4_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_350_itm_1, and_dcpl_78);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_27_mx1w0 = weight_mem_read_arbxbar_arbiters_next_3_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[3]);
  assign Arbiter_8U_Roundrobin_pick_nand_42_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1)
      & and_dcpl_78)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_31_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1
      & and_dcpl_78;
  assign weight_mem_read_arbxbar_arbiters_next_3_1_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_27_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_3_1_sva, Arbiter_8U_Roundrobin_pick_1_mux_250_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_nand_42_cse , Arbiter_8U_Roundrobin_pick_and_31_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_26_mx1w0 = weight_mem_read_arbxbar_arbiters_next_3_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[3]);
  assign weight_mem_read_arbxbar_arbiters_next_3_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_26_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_3_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_249_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_nand_42_cse , Arbiter_8U_Roundrobin_pick_and_31_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_25_mx1w0 = weight_mem_read_arbxbar_arbiters_next_3_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[3]);
  assign weight_mem_read_arbxbar_arbiters_next_3_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_25_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_3_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_248_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_nand_42_cse , Arbiter_8U_Roundrobin_pick_and_31_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_24_mx1w0 = weight_mem_read_arbxbar_arbiters_next_3_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[3]);
  assign weight_mem_read_arbxbar_arbiters_next_3_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_24_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_3_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_247_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_nand_42_cse , Arbiter_8U_Roundrobin_pick_and_31_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_23_mx1w0 = weight_mem_read_arbxbar_arbiters_next_3_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[3]);
  assign weight_mem_read_arbxbar_arbiters_next_3_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_23_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_3_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_246_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_nand_42_cse , Arbiter_8U_Roundrobin_pick_and_31_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_22_mx1w0 = weight_mem_read_arbxbar_arbiters_next_3_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[3]);
  assign weight_mem_read_arbxbar_arbiters_next_3_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_22_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_3_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_245_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_nand_42_cse , Arbiter_8U_Roundrobin_pick_and_31_cse});
  assign weight_mem_read_arbxbar_arbiters_next_3_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_277_itm_1, and_dcpl_78);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_20_mx1w0 = weight_mem_read_arbxbar_arbiters_next_2_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2]);
  assign Arbiter_8U_Roundrobin_pick_nand_30_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1)
      & and_dcpl_78)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_25_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1
      & and_dcpl_78;
  assign weight_mem_read_arbxbar_arbiters_next_2_1_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_20_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_2_1_sva, Arbiter_8U_Roundrobin_pick_1_mux_177_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_nand_30_cse , Arbiter_8U_Roundrobin_pick_and_25_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_19_mx1w0 = weight_mem_read_arbxbar_arbiters_next_2_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2]);
  assign weight_mem_read_arbxbar_arbiters_next_2_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_19_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_2_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_176_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_nand_30_cse , Arbiter_8U_Roundrobin_pick_and_25_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_18_mx1w0 = weight_mem_read_arbxbar_arbiters_next_2_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2]);
  assign weight_mem_read_arbxbar_arbiters_next_2_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_18_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_2_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_175_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_nand_30_cse , Arbiter_8U_Roundrobin_pick_and_25_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_17_mx1w0 = weight_mem_read_arbxbar_arbiters_next_2_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2]);
  assign weight_mem_read_arbxbar_arbiters_next_2_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_17_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_2_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_174_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_nand_30_cse , Arbiter_8U_Roundrobin_pick_and_25_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_16_mx1w0 = weight_mem_read_arbxbar_arbiters_next_2_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2]);
  assign weight_mem_read_arbxbar_arbiters_next_2_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_16_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_2_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_173_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_nand_30_cse , Arbiter_8U_Roundrobin_pick_and_25_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_15_mx1w0 = weight_mem_read_arbxbar_arbiters_next_2_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[2]);
  assign weight_mem_read_arbxbar_arbiters_next_2_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_15_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_2_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_172_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_nand_30_cse , Arbiter_8U_Roundrobin_pick_and_25_cse});
  assign weight_mem_read_arbxbar_arbiters_next_2_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_204_itm_1, and_dcpl_78);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_13_mx1w0 = weight_mem_read_arbxbar_arbiters_next_1_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign Arbiter_8U_Roundrobin_pick_nand_18_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1)
      & and_dcpl_78)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_19_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1
      & and_dcpl_78;
  assign weight_mem_read_arbxbar_arbiters_next_1_1_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_13_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_1_1_sva, Arbiter_8U_Roundrobin_pick_1_mux_104_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_nand_18_cse , Arbiter_8U_Roundrobin_pick_and_19_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_12_mx1w0 = weight_mem_read_arbxbar_arbiters_next_1_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign weight_mem_read_arbxbar_arbiters_next_1_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_12_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_1_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_103_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_nand_18_cse , Arbiter_8U_Roundrobin_pick_and_19_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_11_mx1w0 = weight_mem_read_arbxbar_arbiters_next_1_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign weight_mem_read_arbxbar_arbiters_next_1_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_11_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_1_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_102_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_nand_18_cse , Arbiter_8U_Roundrobin_pick_and_19_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_10_mx1w0 = weight_mem_read_arbxbar_arbiters_next_1_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign weight_mem_read_arbxbar_arbiters_next_1_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_10_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_1_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_101_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_nand_18_cse , Arbiter_8U_Roundrobin_pick_and_19_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_9_mx1w0 = weight_mem_read_arbxbar_arbiters_next_1_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign weight_mem_read_arbxbar_arbiters_next_1_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_9_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_1_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_100_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_nand_18_cse , Arbiter_8U_Roundrobin_pick_and_19_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_8_mx1w0 = weight_mem_read_arbxbar_arbiters_next_1_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[1]);
  assign weight_mem_read_arbxbar_arbiters_next_1_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_8_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_1_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_99_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_nand_18_cse , Arbiter_8U_Roundrobin_pick_and_19_cse});
  assign weight_mem_read_arbxbar_arbiters_next_1_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_131_itm_1, and_dcpl_78);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_6_mx1w0 = weight_mem_read_arbxbar_arbiters_next_0_1_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[0]);
  assign Arbiter_8U_Roundrobin_pick_nand_6_cse = ~((~((~ Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1)
      & and_dcpl_78)) & while_stage_0_5);
  assign Arbiter_8U_Roundrobin_pick_and_13_cse = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1
      & and_dcpl_78;
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_5_mx1w0 = weight_mem_read_arbxbar_arbiters_next_0_2_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[0]);
  assign weight_mem_read_arbxbar_arbiters_next_0_2_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_5_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_0_2_sva, Arbiter_8U_Roundrobin_pick_1_mux_30_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_nand_6_cse , Arbiter_8U_Roundrobin_pick_and_13_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_100_nl = weight_mem_read_arbxbar_arbiters_next_0_3_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[0]);
  assign weight_mem_read_arbxbar_arbiters_next_0_3_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_100_nl,
      weight_mem_read_arbxbar_arbiters_next_0_3_sva, Arbiter_8U_Roundrobin_pick_1_mux_29_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_nand_6_cse , Arbiter_8U_Roundrobin_pick_and_13_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_101_nl = weight_mem_read_arbxbar_arbiters_next_0_4_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[0]);
  assign weight_mem_read_arbxbar_arbiters_next_0_4_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_101_nl,
      weight_mem_read_arbxbar_arbiters_next_0_4_sva, Arbiter_8U_Roundrobin_pick_1_mux_28_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_nand_6_cse , Arbiter_8U_Roundrobin_pick_and_13_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_2_mx1w0 = weight_mem_read_arbxbar_arbiters_next_0_5_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[0]);
  assign weight_mem_read_arbxbar_arbiters_next_0_5_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_2_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_0_5_sva, Arbiter_8U_Roundrobin_pick_1_mux_27_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_nand_6_cse , Arbiter_8U_Roundrobin_pick_and_13_cse});
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_1_mx1w0 = weight_mem_read_arbxbar_arbiters_next_0_6_sva
      | (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[0]);
  assign weight_mem_read_arbxbar_arbiters_next_0_6_sva_mx1 = MUX1HOT_s_1_3_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_1_mx1w0,
      weight_mem_read_arbxbar_arbiters_next_0_6_sva, Arbiter_8U_Roundrobin_pick_1_mux_26_itm_1,
      {and_dcpl_69 , Arbiter_8U_Roundrobin_pick_nand_6_cse , Arbiter_8U_Roundrobin_pick_and_13_cse});
  assign weight_mem_read_arbxbar_arbiters_next_0_7_sva_mx0 = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1,
      Arbiter_8U_Roundrobin_pick_1_mux_57_itm_1, and_dcpl_78);
  assign pe_manager_base_weight_sva_mx1_3_0 = MUX_v_4_2_2((pe_manager_base_weight_sva[3:0]),
      (pe_manager_base_weight_sva_dfm_3_1[3:0]), while_stage_0_5);
  assign pe_manager_base_weight_sva_mx2 = MUX_v_15_2_2(pe_manager_base_weight_sva,
      pe_manager_base_weight_sva_dfm_3_1, while_stage_0_5);
  assign nl_PECore_RunFSM_case_2_for_2_operator_15_false_acc_nl = ({PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1
      , pe_manager_base_weight_sva_mx1_3_0}) + 15'b000000000000001;
  assign PECore_RunFSM_case_2_for_2_operator_15_false_acc_nl = nl_PECore_RunFSM_case_2_for_2_operator_15_false_acc_nl[14:0];
  assign weight_read_addrs_1_lpi_1_dfm_1_1 = MUX_v_15_2_2(15'b000000000000000, PECore_RunFSM_case_2_for_2_operator_15_false_acc_nl,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign nl_operator_15_false_acc_nl = ({PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1
      , (pe_manager_base_weight_sva_mx2[3:1])}) + 14'b00000000000001;
  assign operator_15_false_acc_nl = nl_operator_15_false_acc_nl[13:0];
  assign weight_read_addrs_2_14_1_lpi_1_dfm_1_1 = MUX_v_14_2_2(14'b00000000000000,
      operator_15_false_acc_nl, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign nl_PECore_RunFSM_case_2_for_4_operator_15_false_acc_nl = ({PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1
      , pe_manager_base_weight_sva_mx1_3_0}) + 15'b000000000000011;
  assign PECore_RunFSM_case_2_for_4_operator_15_false_acc_nl = nl_PECore_RunFSM_case_2_for_4_operator_15_false_acc_nl[14:0];
  assign weight_read_addrs_3_lpi_1_dfm_1_1 = MUX_v_15_2_2(15'b000000000000000, PECore_RunFSM_case_2_for_4_operator_15_false_acc_nl,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign nl_operator_15_false_acc_1_nl = ({PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1
      , (pe_manager_base_weight_sva_mx2[3:2])}) + 13'b0000000000001;
  assign operator_15_false_acc_1_nl = nl_operator_15_false_acc_1_nl[12:0];
  assign weight_read_addrs_4_14_2_lpi_1_dfm_1_1 = MUX_v_13_2_2(13'b0000000000000,
      operator_15_false_acc_1_nl, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign nl_PECore_RunFSM_case_2_for_6_operator_15_false_acc_nl = ({PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1
      , pe_manager_base_weight_sva_mx1_3_0}) + 15'b000000000000101;
  assign PECore_RunFSM_case_2_for_6_operator_15_false_acc_nl = nl_PECore_RunFSM_case_2_for_6_operator_15_false_acc_nl[14:0];
  assign weight_read_addrs_5_lpi_1_dfm_1_1 = MUX_v_15_2_2(15'b000000000000000, PECore_RunFSM_case_2_for_6_operator_15_false_acc_nl,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign nl_operator_15_false_acc_2_nl = ({PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1
      , (pe_manager_base_weight_sva_mx2[3:1])}) + 14'b00000000000011;
  assign operator_15_false_acc_2_nl = nl_operator_15_false_acc_2_nl[13:0];
  assign weight_read_addrs_6_14_1_lpi_1_dfm_1_1 = MUX_v_14_2_2(14'b00000000000000,
      operator_15_false_acc_2_nl, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign nl_PECore_RunFSM_case_2_for_8_operator_15_false_acc_nl = ({PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1
      , pe_manager_base_weight_sva_mx1_3_0}) + 15'b000000000000111;
  assign PECore_RunFSM_case_2_for_8_operator_15_false_acc_nl = nl_PECore_RunFSM_case_2_for_8_operator_15_false_acc_nl[14:0];
  assign weight_read_addrs_7_lpi_1_dfm_1_1 = MUX_v_15_2_2(15'b000000000000000, PECore_RunFSM_case_2_for_8_operator_15_false_acc_nl,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_22_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112, and_100_cse);
  assign Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_2 = Arbiter_8U_Roundrobin_pick_1_if_1_mux_22_nl
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
  assign Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[7]);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_20_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97, and_dcpl_533);
  assign Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_2 = Arbiter_8U_Roundrobin_pick_1_if_1_mux_20_nl
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9;
  assign Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[6]);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_18_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82, and_114_cse);
  assign Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_2 = Arbiter_8U_Roundrobin_pick_1_if_1_mux_18_nl
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_10;
  assign Arbiter_8U_Roundrobin_pick_1_unequal_tmp_10 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[5]);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_13 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_13 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_13 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_13 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_13 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_13 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_13 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_16_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67, and_dcpl_547);
  assign Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_2 = Arbiter_8U_Roundrobin_pick_1_if_1_mux_16_nl
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11;
  assign Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[4]);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_12 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_12 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_12 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_12 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_12 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_12 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_12 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_14_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52, and_dcpl_554);
  assign Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_2 = Arbiter_8U_Roundrobin_pick_1_if_1_mux_14_nl
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_12;
  assign Arbiter_8U_Roundrobin_pick_1_unequal_tmp_12 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[3]);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_11 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_11 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_11 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_11 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_11 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_11 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_11 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_12_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37, and_dcpl_561);
  assign Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_2 = Arbiter_8U_Roundrobin_pick_1_if_1_mux_12_nl
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_13;
  assign Arbiter_8U_Roundrobin_pick_1_unequal_tmp_13 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[2]);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_10 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_10 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_10 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_10 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_10 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_10 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_10 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_10_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22, and_dcpl_568);
  assign Arbiter_8U_Roundrobin_pick_return_1_0_2_lpi_1_dfm_2 = Arbiter_8U_Roundrobin_pick_1_if_1_mux_10_nl
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_14;
  assign Arbiter_8U_Roundrobin_pick_1_unequal_tmp_14 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[1]);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_9 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_9 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_9 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_9 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_9 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_9 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_9 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_mux_8_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7_mx0w0,
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7, and_149_cse);
  assign Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_2 = Arbiter_8U_Roundrobin_pick_1_if_1_mux_8_nl
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_15;
  assign Arbiter_8U_Roundrobin_pick_1_unequal_tmp_15 = (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0]);
  assign accum_vector_data_6_sva_1_load_mx0w1 = PECore_UpdateFSM_switch_lp_equal_tmp_2_1
      | accum_vector_data_6_sva_1_load;
  assign PECore_RunFSM_switch_lp_equal_tmp_1_mx0w1 = (state_2_1_sva[0]) & nor_340_cse;
  assign state_mux_1_cse = MUX_v_2_2_2(state_2_1_sva, state_2_1_sva_dfm_1, while_stage_0_3);
  assign state_0_sva_mx1 = MUX_s_1_2_2(PECore_UpdateFSM_next_state_0_lpi_1_dfm_4,
      state_0_sva, or_dcpl_616);
  assign pe_config_manager_counter_sva_mx1 = MUX_v_4_2_2(pe_config_manager_counter_sva,
      pe_config_manager_counter_sva_dfm_3_1, and_1065_cse);
  assign PECore_PushOutput_PECore_PushOutput_if_and_svs_1 = (state_mux_1_cse[1])
      & (~((state_mux_1_cse[0]) | state_0_sva_mx1));
  assign PECore_DecodeAxiWrite_switch_lp_nor_tmp_1_1 = ~(PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_and_5
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0 | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0);
  assign PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva_mx1
      = MUX_s_1_2_2(input_port_PopNB_mioi_return_rsc_z_mxwt, PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva,
      or_dcpl_632);
  assign pe_config_input_counter_and_cse = while_if_and_tmp_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign while_and_4_cse = PECore_UpdateFSM_switch_lp_equal_tmp_3_1 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign nl_operator_8_false_acc_nl = pe_config_input_counter_sva + 8'b00000001;
  assign operator_8_false_acc_nl = nl_operator_8_false_acc_nl[7:0];
  assign pe_config_UpdateInputCounter_not_nl = ~ pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_nor_mdf_sva_st_1;
  assign pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_and_nl = MUX_v_8_2_2(8'b00000000,
      operator_8_false_acc_nl, pe_config_UpdateInputCounter_not_nl);
  assign pe_config_input_counter_nand_nl = ~(while_stage_0_3 & (~((~(PECore_UpdateFSM_switch_lp_equal_tmp_3_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | while_and_1129_cse_1)));
  assign pe_config_input_counter_sva_mx1 = MUX1HOT_v_8_3_2(pe_config_input_counter_sva,
      pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_and_nl, pe_config_input_counter_sva_dfm_1,
      {pe_config_input_counter_nand_nl , while_and_4_cse , pe_config_input_counter_and_cse});
  assign nl_operator_8_false_1_acc_nl = pe_config_output_counter_sva + 8'b00000001;
  assign operator_8_false_1_acc_nl = nl_operator_8_false_1_acc_nl[7:0];
  assign pe_config_UpdateManagerCounter_if_not_9_nl = ~ pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_if_nor_mdf_sva_1;
  assign pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_and_1_nl
      = MUX_v_8_2_2(8'b00000000, operator_8_false_1_acc_nl, pe_config_UpdateManagerCounter_if_not_9_nl);
  assign pe_config_output_counter_nand_nl = ~(while_stage_0_3 & (~((~(and_2257_cse
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | while_and_1129_cse_1)));
  assign while_and_63_nl = and_2257_cse & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign pe_config_output_counter_sva_mx1 = MUX1HOT_v_8_3_2(pe_config_output_counter_sva,
      pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_and_1_nl,
      pe_config_output_counter_sva_dfm_1, {pe_config_output_counter_nand_nl , while_and_63_nl
      , pe_config_input_counter_and_cse});
  assign while_if_and_2_m1c = PECore_UpdateFSM_switch_lp_equal_tmp_5_1 & and_dcpl_204;
  assign pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_and_nl
      = pe_config_is_zero_first_sva & (~ pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_if_nor_mdf_sva_1);
  assign while_if_or_nl = (~((~((~ PECore_UpdateFSM_switch_lp_equal_tmp_5_1) & and_dcpl_204))
      & while_stage_0_3)) | ((~ pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1)
      & while_if_and_2_m1c);
  assign while_if_and_4_nl = pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1
      & while_if_and_2_m1c;
  assign pe_config_is_zero_first_sva_mx1 = MUX1HOT_s_1_3_2(while_if_mux_19_itm_1,
      pe_config_is_zero_first_sva, pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_and_nl,
      {and_dcpl_203 , while_if_or_nl , while_if_and_4_nl});
  assign PECore_UpdateFSM_switch_lp_equal_tmp_6 = state_0_sva_mx1 & (state_mux_1_cse==2'b00);
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_1_cse_1 = (state_mux_1_cse[0])
      & (~((state_mux_1_cse[1]) | state_0_sva_mx1));
  assign pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1_1
      = ~((pe_config_manager_counter_sva_mx1 != (operator_4_false_acc_sdt_sva_1[3:0]))
      | (operator_4_false_acc_sdt_sva_1[4]));
  assign PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:16]==4'b0110);
  assign PECore_UpdateFSM_switch_lp_not_23_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_15_nl
      = MUX_v_20_2_2(20'b00000000000000000000, act_port_reg_data_19_0_sva_dfm_1_1,
      PECore_UpdateFSM_switch_lp_not_23_nl);
  assign act_port_reg_data_19_0_sva_mx1 = MUX_v_20_2_2(PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_15_nl,
      act_port_reg_data_19_0_sva, or_dcpl_635);
  assign PECore_UpdateFSM_switch_lp_not_24_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_14_nl
      = MUX_v_20_2_2(20'b00000000000000000000, act_port_reg_data_51_32_sva_dfm_1_1,
      PECore_UpdateFSM_switch_lp_not_24_nl);
  assign act_port_reg_data_51_32_sva_mx1 = MUX_v_20_2_2(PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_14_nl,
      act_port_reg_data_51_32_sva, or_dcpl_635);
  assign PECore_UpdateFSM_switch_lp_not_25_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_13_nl
      = MUX_v_20_2_2(20'b00000000000000000000, act_port_reg_data_83_64_sva_dfm_1_1,
      PECore_UpdateFSM_switch_lp_not_25_nl);
  assign act_port_reg_data_83_64_sva_mx1 = MUX_v_20_2_2(PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_13_nl,
      act_port_reg_data_83_64_sva, or_dcpl_635);
  assign PECore_UpdateFSM_switch_lp_not_26_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_12_nl
      = MUX_v_20_2_2(20'b00000000000000000000, act_port_reg_data_115_96_sva_dfm_1_1,
      PECore_UpdateFSM_switch_lp_not_26_nl);
  assign act_port_reg_data_115_96_sva_mx1 = MUX_v_20_2_2(PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_12_nl,
      act_port_reg_data_115_96_sva, or_dcpl_635);
  assign PECore_UpdateFSM_switch_lp_not_27_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_11_nl
      = MUX_v_20_2_2(20'b00000000000000000000, act_port_reg_data_147_128_sva_dfm_1_1,
      PECore_UpdateFSM_switch_lp_not_27_nl);
  assign act_port_reg_data_147_128_sva_mx1 = MUX_v_20_2_2(PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_11_nl,
      act_port_reg_data_147_128_sva, or_dcpl_635);
  assign PECore_UpdateFSM_switch_lp_not_28_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_10_nl
      = MUX_v_20_2_2(20'b00000000000000000000, act_port_reg_data_179_160_sva_dfm_1_1,
      PECore_UpdateFSM_switch_lp_not_28_nl);
  assign act_port_reg_data_179_160_sva_mx1 = MUX_v_20_2_2(PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_10_nl,
      act_port_reg_data_179_160_sva, or_dcpl_635);
  assign PECore_UpdateFSM_switch_lp_not_29_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_9_nl
      = MUX_v_20_2_2(20'b00000000000000000000, act_port_reg_data_211_192_sva_dfm_1_1,
      PECore_UpdateFSM_switch_lp_not_29_nl);
  assign act_port_reg_data_211_192_sva_mx1 = MUX_v_20_2_2(PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_9_nl,
      act_port_reg_data_211_192_sva, or_dcpl_635);
  assign PECore_UpdateFSM_switch_lp_not_19_nl = ~ PECore_UpdateFSM_switch_lp_equal_tmp_2_9;
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_8_nl
      = MUX_v_20_2_2(20'b00000000000000000000, act_port_reg_data_243_224_sva_dfm_1_1,
      PECore_UpdateFSM_switch_lp_not_19_nl);
  assign act_port_reg_data_243_224_sva_mx1 = MUX_v_20_2_2(PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_8_nl,
      act_port_reg_data_243_224_sva, or_dcpl_635);
  assign while_and_24_cse = crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
  assign while_and_23_cse = (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3)
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
  assign while_while_nor_259_cse = ~(weight_mem_run_3_for_land_1_lpi_1_dfm_3 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign while_and_1123_rgt = weight_mem_run_3_for_land_1_lpi_1_dfm_3 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_94_itm_1 = (weight_read_addrs_3_lpi_1_dfm_2_2_0==3'b101)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_71_itm_1_1 = (weight_read_addrs_3_lpi_1_dfm_2_2_0==3'b110)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_72_itm_1_1 = (weight_read_addrs_3_lpi_1_dfm_2_2_0==3'b111)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_and_49_tmp = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2==3'b111)
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2;
  assign weight_mem_run_3_for_land_lpi_1_dfm_1_1 = PECore_RunFSM_switch_lp_equal_tmp_1_2
      & (Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_1
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_1
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_1
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6_1);
  assign weight_mem_run_3_for_land_6_lpi_1_dfm_1_1 = PECore_RunFSM_switch_lp_equal_tmp_1_2
      & (Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_4_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_1
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_4_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_1
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_1
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4_1);
  assign weight_mem_run_3_for_land_4_lpi_1_dfm_1_1 = PECore_RunFSM_switch_lp_equal_tmp_1_2
      & (Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_38_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_50_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_62_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_74_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_86_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_98_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_110_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_122_tmp);
  assign weight_mem_read_arbxbar_xbar_1_for_3_8_for_2_or_cse = Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_42_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_54_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_66_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_78_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_90_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_102_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_114_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_126_tmp;
  assign weight_mem_run_3_for_land_2_lpi_1_dfm_1_1 = PECore_RunFSM_switch_lp_equal_tmp_1_2
      & weight_mem_read_arbxbar_xbar_1_for_3_8_for_2_or_cse;
  assign weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp
      = Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_101_tmp
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_22_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_98_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_100_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_102_tmp | Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_1_1;
  assign weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp
      = Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_89_tmp
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_18_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_86_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_88_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_90_tmp | Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_1_1;
  assign weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp
      = Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_77_tmp
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_14_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_74_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_76_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_78_tmp | Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_1_1;
  assign weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp
      = Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_65_tmp
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_4_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_10_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_62_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_64_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_66_tmp | Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_1_1;
  assign weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp
      = Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_53_tmp
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_6_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_50_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_52_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_54_tmp | Arbiter_8U_Roundrobin_pick_return_1_0_2_lpi_1_dfm_1_1;
  assign weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp
      = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_6_1 | and_703_cse |
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_4_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_2_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_38_tmp | and_700_cse
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_42_tmp | Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_1_1;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6_mx1
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_6_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6,
      or_dcpl_615);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0_mx1
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_0_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0,
      or_dcpl_615);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5_mx1
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_5_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5,
      or_dcpl_615);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1_mx1
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_1_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1,
      or_dcpl_615);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4_mx1
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_4_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4,
      or_dcpl_615);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2_mx1
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_2_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2,
      or_dcpl_615);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3_mx1
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_3_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3,
      or_dcpl_615);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_15 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_15 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_15 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_15 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_15 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_15 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_15 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_14 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_14 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_14 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_14 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_14 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_14 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_14 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_8
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_9
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_2_sva_1);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_10
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_3_sva_1);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_11
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_4_sva_1);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_12
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_5_sva_1);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_13
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_14
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_7_sva_1);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112_mx0w0 = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_15
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_sva_1);
  assign PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:16]==4'b0101);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_1 = (pe_manager_base_weight_sva[2:0]==3'b111)
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_1 = (pe_manager_base_weight_sva[2:0]==3'b110)
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_9_itm_1 = (pe_manager_base_weight_sva[2:0]==3'b100)
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_7_itm_1 = (pe_manager_base_weight_sva[2:0]==3'b010)
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_6_itm_1 = (pe_manager_base_weight_sva[2:0]==3'b001)
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_95_itm_mx0w0 = (weight_read_addrs_3_lpi_1_dfm_1[2:0]==3'b110)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_1_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_mx0w0 = (weight_read_addrs_3_lpi_1_dfm_1[2:0]==3'b101)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_1_1;
  assign weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp
      = Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6_1 | and_702_cse | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4_1
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_30_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_122_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_124_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_126_tmp
      | Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_1_1;
  assign weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp
      = Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_113_tmp
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4_1 | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_26_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_110_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_112_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_114_tmp | Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_1_1;
  assign ProductSum_for_mux_nl = MUX_v_23_2_2(accum_vector_data_7_sva_5, ProductSum_for_acc_9_cmp_z,
      reg_PECore_RunMac_PECore_RunMac_if_and_svs_st_8_cse);
  assign accum_vector_operator_1_for_not_61_nl = ~ accum_vector_operator_1_for_asn_64_itm_7;
  assign accum_vector_data_7_sva_5_mx1w0 = MUX_v_23_2_2(23'b00000000000000000000000,
      ProductSum_for_mux_nl, accum_vector_operator_1_for_not_61_nl);
  assign ProductSum_for_mux_1_nl = MUX_v_23_2_2(accum_vector_data_7_sva_4, ProductSum_for_acc_8_cmp_z,
      reg_PECore_RunMac_PECore_RunMac_if_and_svs_st_8_cse);
  assign accum_vector_operator_1_for_not_38_nl = ~ accum_vector_operator_1_for_asn_64_itm_7;
  assign accum_vector_data_7_sva_4_mx0w0 = MUX_v_23_2_2(23'b00000000000000000000000,
      ProductSum_for_mux_1_nl, accum_vector_operator_1_for_not_38_nl);
  assign ProductSum_for_mux_2_nl = MUX_v_23_2_2(accum_vector_data_6_sva_5, PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_z,
      reg_PECore_RunMac_PECore_RunMac_if_and_svs_st_8_cse);
  assign accum_vector_operator_1_for_not_62_nl = ~ accum_vector_operator_1_for_asn_55_itm_7;
  assign accum_vector_data_6_sva_5_mx1w0 = MUX_v_23_2_2(23'b00000000000000000000000,
      ProductSum_for_mux_2_nl, accum_vector_operator_1_for_not_62_nl);
  assign ProductSum_for_mux_3_nl = MUX_v_23_2_2(accum_vector_data_6_sva_4, PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_z,
      reg_PECore_RunMac_PECore_RunMac_if_and_svs_st_8_cse);
  assign accum_vector_operator_1_for_not_40_nl = ~ accum_vector_operator_1_for_asn_55_itm_7;
  assign accum_vector_data_6_sva_4_mx0w0 = MUX_v_23_2_2(23'b00000000000000000000000,
      ProductSum_for_mux_3_nl, accum_vector_operator_1_for_not_40_nl);
  assign ProductSum_for_mux_4_nl = MUX_v_23_2_2(accum_vector_data_5_sva_5, PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_z,
      reg_PECore_RunMac_PECore_RunMac_if_and_svs_st_8_cse);
  assign accum_vector_operator_1_for_not_63_nl = ~ accum_vector_operator_1_for_asn_46_itm_7;
  assign accum_vector_data_5_sva_5_mx0w0 = MUX_v_23_2_2(23'b00000000000000000000000,
      ProductSum_for_mux_4_nl, accum_vector_operator_1_for_not_63_nl);
  assign ProductSum_for_mux_5_nl = MUX_v_23_2_2(accum_vector_data_5_sva_4, PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_z,
      reg_PECore_RunMac_PECore_RunMac_if_and_svs_st_8_cse);
  assign accum_vector_operator_1_for_not_42_nl = ~ accum_vector_operator_1_for_asn_46_itm_7;
  assign accum_vector_data_5_sva_4_mx1w0 = MUX_v_23_2_2(23'b00000000000000000000000,
      ProductSum_for_mux_5_nl, accum_vector_operator_1_for_not_42_nl);
  assign ProductSum_for_mux_6_nl = MUX_v_23_2_2(accum_vector_data_4_sva_5, PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_z,
      reg_PECore_RunMac_PECore_RunMac_if_and_svs_st_8_cse);
  assign accum_vector_operator_1_for_not_64_nl = ~ accum_vector_operator_1_for_asn_37_itm_7;
  assign accum_vector_data_4_sva_5_mx1w0 = MUX_v_23_2_2(23'b00000000000000000000000,
      ProductSum_for_mux_6_nl, accum_vector_operator_1_for_not_64_nl);
  assign ProductSum_for_mux_7_nl = MUX_v_23_2_2(accum_vector_data_4_sva_4, PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_z,
      reg_PECore_RunMac_PECore_RunMac_if_and_svs_st_8_cse);
  assign accum_vector_operator_1_for_not_44_nl = ~ accum_vector_operator_1_for_asn_37_itm_7;
  assign accum_vector_data_4_sva_4_mx1w0 = MUX_v_23_2_2(23'b00000000000000000000000,
      ProductSum_for_mux_7_nl, accum_vector_operator_1_for_not_44_nl);
  assign ProductSum_for_mux_8_nl = MUX_v_23_2_2(accum_vector_data_3_sva_5, PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_z,
      reg_PECore_RunMac_PECore_RunMac_if_and_svs_st_8_cse);
  assign accum_vector_operator_1_for_not_65_nl = ~ accum_vector_operator_1_for_asn_28_itm_7;
  assign accum_vector_data_3_sva_5_mx1w0 = MUX_v_23_2_2(23'b00000000000000000000000,
      ProductSum_for_mux_8_nl, accum_vector_operator_1_for_not_65_nl);
  assign ProductSum_for_mux_9_nl = MUX_v_23_2_2(accum_vector_data_3_sva_4, PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_z,
      reg_PECore_RunMac_PECore_RunMac_if_and_svs_st_8_cse);
  assign accum_vector_operator_1_for_not_46_nl = ~ accum_vector_operator_1_for_asn_28_itm_7;
  assign accum_vector_data_3_sva_4_mx1w0 = MUX_v_23_2_2(23'b00000000000000000000000,
      ProductSum_for_mux_9_nl, accum_vector_operator_1_for_not_46_nl);
  assign ProductSum_for_mux_10_nl = MUX_v_23_2_2(accum_vector_data_2_sva_6, PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_z,
      reg_PECore_RunMac_PECore_RunMac_if_and_svs_st_8_cse);
  assign accum_vector_operator_1_for_not_66_nl = ~ accum_vector_operator_1_for_asn_22_itm_7;
  assign accum_vector_data_2_sva_6_mx1w0 = MUX_v_23_2_2(23'b00000000000000000000000,
      ProductSum_for_mux_10_nl, accum_vector_operator_1_for_not_66_nl);
  assign ProductSum_for_mux_11_nl = MUX_v_23_2_2(accum_vector_data_2_sva_5, PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_z,
      reg_PECore_RunMac_PECore_RunMac_if_and_svs_st_8_cse);
  assign accum_vector_operator_1_for_not_67_nl = ~ accum_vector_operator_1_for_asn_22_itm_7;
  assign accum_vector_data_2_sva_5_mx1w0 = MUX_v_23_2_2(23'b00000000000000000000000,
      ProductSum_for_mux_11_nl, accum_vector_operator_1_for_not_67_nl);
  assign ProductSum_for_mux_12_nl = MUX_v_23_2_2(accum_vector_data_2_sva_4, PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_z,
      reg_PECore_RunMac_PECore_RunMac_if_and_svs_st_8_cse);
  assign accum_vector_operator_1_for_not_48_nl = ~ accum_vector_operator_1_for_asn_22_itm_7;
  assign accum_vector_data_2_sva_4_mx1w0 = MUX_v_23_2_2(23'b00000000000000000000000,
      ProductSum_for_mux_12_nl, accum_vector_operator_1_for_not_48_nl);
  assign ProductSum_for_mux_13_nl = MUX_v_23_2_2(accum_vector_data_1_sva_5, PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_z,
      reg_PECore_RunMac_PECore_RunMac_if_and_svs_st_8_cse);
  assign accum_vector_operator_1_for_not_68_nl = ~ accum_vector_operator_1_for_asn_10_itm_7;
  assign accum_vector_data_1_sva_5_mx1w0 = MUX_v_23_2_2(23'b00000000000000000000000,
      ProductSum_for_mux_13_nl, accum_vector_operator_1_for_not_68_nl);
  assign ProductSum_for_mux_14_nl = MUX_v_23_2_2(accum_vector_data_1_sva_4, PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_z,
      reg_PECore_RunMac_PECore_RunMac_if_and_svs_st_8_cse);
  assign accum_vector_operator_1_for_not_50_nl = ~ accum_vector_operator_1_for_asn_10_itm_7;
  assign accum_vector_data_1_sva_4_mx1w0 = MUX_v_23_2_2(23'b00000000000000000000000,
      ProductSum_for_mux_14_nl, accum_vector_operator_1_for_not_50_nl);
  assign ProductSum_for_mux_15_nl = MUX_v_23_2_2(accum_vector_data_0_sva_5, PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_z,
      reg_PECore_RunMac_PECore_RunMac_if_and_svs_st_8_cse);
  assign accum_vector_operator_1_for_not_69_nl = ~ accum_vector_operator_1_for_asn_1_itm_7;
  assign accum_vector_data_0_sva_5_mx1w0 = MUX_v_23_2_2(23'b00000000000000000000000,
      ProductSum_for_mux_15_nl, accum_vector_operator_1_for_not_69_nl);
  assign ProductSum_for_mux_16_nl = MUX_v_23_2_2(accum_vector_data_0_sva_4, PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_z,
      reg_PECore_RunMac_PECore_RunMac_if_and_svs_st_8_cse);
  assign accum_vector_operator_1_for_not_52_nl = ~ accum_vector_operator_1_for_asn_1_itm_7;
  assign accum_vector_data_0_sva_4_mx1w0 = MUX_v_23_2_2(23'b00000000000000000000000,
      ProductSum_for_mux_16_nl, accum_vector_operator_1_for_not_52_nl);
  assign weight_mem_run_3_for_land_1_lpi_1_dfm_1_1 = PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2
      & (Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_2 | Arbiter_8U_Roundrobin_pick_return_1_0_2_lpi_1_dfm_2
      | Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_2 | Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_2
      | Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_2 | Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_2
      | Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_2 | Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_2);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_1_1 = (weight_read_addrs_3_lpi_1_dfm_1[2:0]==3'b011)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_1_1;
  assign ProductSum_for_mux_24_nl = MUX_v_23_2_2(accum_vector_data_7_sva_7, ProductSum_for_acc_11_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_7);
  assign accum_vector_operator_1_for_not_54_nl = ~ accum_vector_operator_1_for_asn_70_itm_6;
  assign accum_vector_data_7_sva_7_mx1w0 = MUX_v_23_2_2(23'b00000000000000000000000,
      ProductSum_for_mux_24_nl, accum_vector_operator_1_for_not_54_nl);
  assign ProductSum_for_mux_25_nl = MUX_v_23_2_2(accum_vector_data_7_sva_6, ProductSum_for_acc_10_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_7);
  assign accum_vector_operator_1_for_not_24_nl = ~ accum_vector_operator_1_for_asn_70_itm_6;
  assign accum_vector_data_7_sva_6_mx1w0 = MUX_v_23_2_2(23'b00000000000000000000000,
      ProductSum_for_mux_25_nl, accum_vector_operator_1_for_not_24_nl);
  assign ProductSum_for_mux_26_nl = MUX_v_23_2_2(accum_vector_data_6_sva_7, PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_7);
  assign accum_vector_operator_1_for_not_55_nl = ~ accum_vector_operator_1_for_asn_61_itm_6;
  assign accum_vector_data_6_sva_7_mx1w0 = MUX_v_23_2_2(23'b00000000000000000000000,
      ProductSum_for_mux_26_nl, accum_vector_operator_1_for_not_55_nl);
  assign ProductSum_for_mux_27_nl = MUX_v_23_2_2(accum_vector_data_6_sva_6, PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_4_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_7);
  assign accum_vector_operator_1_for_not_26_nl = ~ accum_vector_operator_1_for_asn_61_itm_6;
  assign accum_vector_data_6_sva_6_mx1w0 = MUX_v_23_2_2(23'b00000000000000000000000,
      ProductSum_for_mux_27_nl, accum_vector_operator_1_for_not_26_nl);
  assign ProductSum_for_mux_28_nl = MUX_v_23_2_2(accum_vector_data_5_sva_7, PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_7);
  assign accum_vector_operator_1_for_not_56_nl = ~ accum_vector_operator_1_for_asn_52_itm_6;
  assign accum_vector_data_5_sva_7_mx1w0 = MUX_v_23_2_2(23'b00000000000000000000000,
      ProductSum_for_mux_28_nl, accum_vector_operator_1_for_not_56_nl);
  assign ProductSum_for_mux_29_nl = MUX_v_23_2_2(accum_vector_data_5_sva_6, PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_4_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_7);
  assign accum_vector_operator_1_for_not_28_nl = ~ accum_vector_operator_1_for_asn_52_itm_6;
  assign accum_vector_data_5_sva_6_mx1w0 = MUX_v_23_2_2(23'b00000000000000000000000,
      ProductSum_for_mux_29_nl, accum_vector_operator_1_for_not_28_nl);
  assign ProductSum_for_mux_30_nl = MUX_v_23_2_2(accum_vector_data_4_sva_7, PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_7);
  assign accum_vector_operator_1_for_not_57_nl = ~ accum_vector_operator_1_for_asn_43_itm_6;
  assign accum_vector_data_4_sva_7_mx1w0 = MUX_v_23_2_2(23'b00000000000000000000000,
      ProductSum_for_mux_30_nl, accum_vector_operator_1_for_not_57_nl);
  assign ProductSum_for_mux_31_nl = MUX_v_23_2_2(accum_vector_data_4_sva_6, PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_4_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_7);
  assign accum_vector_operator_1_for_not_30_nl = ~ accum_vector_operator_1_for_asn_43_itm_6;
  assign accum_vector_data_4_sva_6_mx1w0 = MUX_v_23_2_2(23'b00000000000000000000000,
      ProductSum_for_mux_31_nl, accum_vector_operator_1_for_not_30_nl);
  assign ProductSum_for_mux_32_nl = MUX_v_23_2_2(accum_vector_data_3_sva_7, PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_7);
  assign accum_vector_operator_1_for_not_58_nl = ~ accum_vector_operator_1_for_asn_34_itm_6;
  assign accum_vector_data_3_sva_7_mx1w0 = MUX_v_23_2_2(23'b00000000000000000000000,
      ProductSum_for_mux_32_nl, accum_vector_operator_1_for_not_58_nl);
  assign ProductSum_for_mux_33_nl = MUX_v_23_2_2(accum_vector_data_3_sva_6, PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_4_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_7);
  assign accum_vector_operator_1_for_not_32_nl = ~ accum_vector_operator_1_for_asn_34_itm_6;
  assign accum_vector_data_3_sva_6_mx1w0 = MUX_v_23_2_2(23'b00000000000000000000000,
      ProductSum_for_mux_33_nl, accum_vector_operator_1_for_not_32_nl);
  assign ProductSum_for_mux_34_nl = MUX_v_23_2_2(accum_vector_data_1_sva_7, PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_7);
  assign accum_vector_operator_1_for_not_59_nl = ~ accum_vector_operator_1_for_asn_16_itm_6;
  assign accum_vector_data_1_sva_7_mx1w0 = MUX_v_23_2_2(23'b00000000000000000000000,
      ProductSum_for_mux_34_nl, accum_vector_operator_1_for_not_59_nl);
  assign ProductSum_for_mux_35_nl = MUX_v_23_2_2(accum_vector_data_1_sva_6, PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_4_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_7);
  assign accum_vector_operator_1_for_not_34_nl = ~ accum_vector_operator_1_for_asn_16_itm_6;
  assign accum_vector_data_1_sva_6_mx1w0 = MUX_v_23_2_2(23'b00000000000000000000000,
      ProductSum_for_mux_35_nl, accum_vector_operator_1_for_not_34_nl);
  assign ProductSum_for_mux_36_nl = MUX_v_23_2_2(accum_vector_data_0_sva_7, PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_7);
  assign accum_vector_operator_1_for_not_60_nl = ~ accum_vector_operator_1_for_asn_7_itm_6;
  assign accum_vector_data_0_sva_7_mx1w0 = MUX_v_23_2_2(23'b00000000000000000000000,
      ProductSum_for_mux_36_nl, accum_vector_operator_1_for_not_60_nl);
  assign ProductSum_for_mux_37_nl = MUX_v_23_2_2(accum_vector_data_0_sva_6, PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_z,
      PECore_RunMac_PECore_RunMac_if_and_svs_st_7);
  assign accum_vector_operator_1_for_not_36_nl = ~ accum_vector_operator_1_for_asn_7_itm_6;
  assign accum_vector_data_0_sva_6_mx1w0 = MUX_v_23_2_2(23'b00000000000000000000000,
      ProductSum_for_mux_37_nl, accum_vector_operator_1_for_not_36_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1_1 = MUX_v_3_2_2(3'b000,
      (weight_read_addrs_0_3_0_lpi_1_dfm_1_2[2:0]), weight_mem_run_1_if_for_weight_mem_run_1_if_for_weight_mem_run_1_if_for_nor_tmp);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_mux_1_tmp = MUX_s_1_8_2((weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[2]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5]), (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6]),
      (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7]), crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1_1);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1_1 = ~(crossbar_spec_PE_Weight_WordType_8U_8U_for_mux_1_tmp
      | (~ weight_mem_run_1_if_for_weight_mem_run_1_if_for_weight_mem_run_1_if_for_nor_tmp));
  assign PECore_PushAxiRsp_mux_23_nl = MUX_s_1_2_2(pe_manager_base_weight_slc_pe_manager_base_weight_0_12_itm_2,
      PECore_PushAxiRsp_mux_10_itm_1, rva_in_reg_rw_sva_5);
  assign PECore_PushAxiRsp_if_else_mux_10_mx0w2 = MUX_s_1_2_2(PECore_PushAxiRsp_mux_23_nl,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[47]), crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_11_itm_1);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_1_cse = ~((reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[2])
      | (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[0]));
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_2_cse = ~((reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1:0]!=2'b00));
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_or_cse = ((reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1])
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_1_cse & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3)
      | ((reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[2]) & crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_2_cse
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign and_923_cse = crossbar_spec_PE_Weight_WordType_8U_8U_for_asn_56 & (~ or_dcpl_683);
  assign and_924_cse = crossbar_spec_PE_Weight_WordType_8U_8U_for_or_cse & (~ or_dcpl_683);
  assign and_925_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_48_itm_1
      & (~ or_dcpl_683);
  assign and_926_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_72_itm_1
      & (~ or_dcpl_683);
  assign and_927_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_79_itm_1
      & (~ or_dcpl_683);
  assign and_928_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_62_itm_1
      & (~ or_dcpl_683);
  assign nor_523_cse = ~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3
      | or_dcpl_683);
  assign and_922_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_for_and_54 & (~ or_dcpl_683);
  assign mux1h_3_nl = MUX1HOT_s_1_8_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_21_itm_1[7]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_itm_1_7,
      (weight_mem_banks_load_store_1_for_3_result_val_Marshall_64U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1[7]),
      (weight_mem_banks_load_store_1_for_5_result_val_Marshall_64U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1[7]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[7]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[7]),
      weight_port_read_out_data_0_0_sva_dfm_2_7, {and_922_ssc , and_923_cse , and_924_cse
      , and_925_cse , and_926_cse , and_927_cse , and_928_cse , nor_523_cse});
  assign weight_port_read_out_data_0_0_sva_dfm_mx0w0_7 = mux1h_3_nl & (~ or_dcpl_683);
  assign mux1h_10_nl = MUX1HOT_v_7_8_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_itm_1[6:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_21_itm_1[6:0]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_itm_1_6_0,
      (weight_mem_banks_load_store_1_for_3_result_val_Marshall_64U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1[6:0]),
      (weight_mem_banks_load_store_1_for_5_result_val_Marshall_64U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1[6:0]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[6:0]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[6:0]),
      weight_port_read_out_data_0_0_sva_dfm_2_6_0, {and_922_ssc , and_923_cse , and_924_cse
      , and_925_cse , and_926_cse , and_927_cse , and_928_cse , nor_523_cse});
  assign not_2545_nl = ~ or_dcpl_683;
  assign weight_port_read_out_data_0_0_sva_dfm_mx0w0_6_0 = MUX_v_7_2_2(7'b0000000,
      mux1h_10_nl, not_2545_nl);
  assign and_931_cse = crossbar_spec_PE_Weight_WordType_8U_8U_for_and_52 & (~ or_dcpl_684);
  assign and_932_cse = crossbar_spec_PE_Weight_WordType_8U_8U_for_asn_56 & (~ or_dcpl_684);
  assign and_933_cse = crossbar_spec_PE_Weight_WordType_8U_8U_for_or_cse & (~ or_dcpl_684);
  assign and_934_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_48_itm_1
      & (~ or_dcpl_684);
  assign and_935_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_60_itm_1
      & (~ or_dcpl_684);
  assign and_936_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_47_itm_1
      & (~ or_dcpl_684);
  assign and_937_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_62_itm_1
      & (~ or_dcpl_684);
  assign nor_524_cse = ~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3
      | or_dcpl_684);
  assign mux1h_4_nl = MUX1HOT_s_1_8_2((rva_out_reg_data_55_48_sva_dfm_1_5[7]), (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_23_itm_1[7]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1_7,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_25_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_41_itm_1[7]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[15]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[15]),
      weight_port_read_out_data_0_1_sva_dfm_2_7, {and_931_cse , and_932_cse , and_933_cse
      , and_934_cse , and_935_cse , and_936_cse , and_937_cse , nor_524_cse});
  assign weight_port_read_out_data_0_1_sva_dfm_mx0w0_7 = mux1h_4_nl & (~ or_dcpl_684);
  assign mux1h_11_nl = MUX1HOT_v_7_8_2((rva_out_reg_data_55_48_sva_dfm_1_5[6:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_23_itm_1[6:0]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1_6_0,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_25_itm_1[6:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_41_itm_1[6:0]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[14:8]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[14:8]),
      weight_port_read_out_data_0_1_sva_dfm_2_6_0, {and_931_cse , and_932_cse , and_933_cse
      , and_934_cse , and_935_cse , and_936_cse , and_937_cse , nor_524_cse});
  assign not_2546_nl = ~ or_dcpl_684;
  assign weight_port_read_out_data_0_1_sva_dfm_mx0w0_6_0 = MUX_v_7_2_2(7'b0000000,
      mux1h_11_nl, not_2546_nl);
  assign and_940_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_for_and_52 & (~ or_dcpl_683);
  assign mux1h_5_nl = MUX1HOT_s_1_8_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1_7,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_itm_1_7,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_itm_1_7_6[1]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_26_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_42_itm_1[7]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[23]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[23]),
      weight_port_read_out_data_0_2_sva_dfm_2_7, {and_940_ssc , and_923_cse , and_924_cse
      , and_925_cse , and_926_cse , and_927_cse , and_928_cse , nor_523_cse});
  assign weight_port_read_out_data_0_2_sva_dfm_mx0w0_7 = mux1h_5_nl & (~ or_dcpl_683);
  assign mux1h_12_nl = MUX1HOT_s_1_8_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1_6_0[6]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_itm_1_6_0[6]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_itm_1_7_6[0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_26_itm_1[6]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_42_itm_1[6]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[22]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[22]),
      weight_port_read_out_data_0_2_sva_dfm_2_6, {and_940_ssc , and_923_cse , and_924_cse
      , and_925_cse , and_926_cse , and_927_cse , and_928_cse , nor_523_cse});
  assign weight_port_read_out_data_0_2_sva_dfm_mx0w0_6 = mux1h_12_nl & (~ or_dcpl_683);
  assign mux1h_13_nl = MUX1HOT_v_6_8_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1_6_0[5:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_itm_1_6_0[5:0]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_itm_1_5_0,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_26_itm_1[5:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_42_itm_1[5:0]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[21:16]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[21:16]),
      weight_port_read_out_data_0_2_sva_dfm_2_5_0, {and_940_ssc , and_923_cse , and_924_cse
      , and_925_cse , and_926_cse , and_927_cse , and_928_cse , nor_523_cse});
  assign not_2547_nl = ~ or_dcpl_683;
  assign weight_port_read_out_data_0_2_sva_dfm_mx0w0_5_0 = MUX_v_6_2_2(6'b000000,
      mux1h_13_nl, not_2547_nl);
  assign mux1h_6_nl = MUX1HOT_s_1_8_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_3_itm_1[7]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1_7,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1_7_4[3]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_27_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_43_itm_1[7]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[31]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[31]),
      weight_port_read_out_data_0_3_sva_dfm_2_7, {and_931_cse , and_932_cse , and_933_cse
      , and_934_cse , and_935_cse , and_936_cse , and_937_cse , nor_524_cse});
  assign weight_port_read_out_data_0_3_sva_dfm_mx0w0_7 = mux1h_6_nl & (~ or_dcpl_684);
  assign mux1h_14_nl = MUX1HOT_v_3_8_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_3_itm_1[6:4]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1_6_0[6:4]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1_7_4[2:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_27_itm_1[6:4]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_43_itm_1[6:4]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[30:28]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[30:28]),
      weight_port_read_out_data_0_3_sva_dfm_2_6_4, {and_931_cse , and_932_cse , and_933_cse
      , and_934_cse , and_935_cse , and_936_cse , and_937_cse , nor_524_cse});
  assign not_2549_nl = ~ or_dcpl_684;
  assign weight_port_read_out_data_0_3_sva_dfm_mx0w0_6_4 = MUX_v_3_2_2(3'b000, mux1h_14_nl,
      not_2549_nl);
  assign mux1h_15_nl = MUX1HOT_v_4_8_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_3_itm_1[3:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1_6_0[3:0]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1_3_0,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_27_itm_1[3:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_43_itm_1[3:0]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[27:24]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[27:24]),
      weight_port_read_out_data_0_3_sva_dfm_2_3_0, {and_931_cse , and_932_cse , and_933_cse
      , and_934_cse , and_935_cse , and_936_cse , and_937_cse , nor_524_cse});
  assign not_2550_nl = ~ or_dcpl_684;
  assign weight_port_read_out_data_0_3_sva_dfm_mx0w0_3_0 = MUX_v_4_2_2(4'b0000, mux1h_15_nl,
      not_2550_nl);
  assign rva_out_reg_data_62_56_sva_dfm_6_mx1 = MUX_v_7_2_2(rva_out_reg_data_62_56_sva_dfm_4_1,
      rva_out_reg_data_62_56_sva_dfm_6, or_dcpl_665);
  assign rva_out_reg_data_35_32_sva_dfm_6_mx1 = MUX_v_4_2_2(rva_out_reg_data_35_32_sva_dfm_4_1,
      rva_out_reg_data_35_32_sva_dfm_6, or_dcpl_665);
  assign input_mem_banks_bank_a_nand_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_2_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_100_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_2_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_101_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_tmp_1 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_0_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_0_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_nl
      , while_and_100_nl , while_and_101_nl});
  assign input_mem_banks_bank_a_nand_1_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_3_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_1_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_104_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_3_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_105_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_1_tmp_1 &
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_1_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_1_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_1_nl
      , while_and_104_nl , while_and_105_nl});
  assign input_mem_banks_bank_a_nand_2_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_4_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_2_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_108_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_4_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_109_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_2_tmp_1 &
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_2_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_2_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_2_nl
      , while_and_108_nl , while_and_109_nl});
  assign input_mem_banks_bank_a_nand_3_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_5_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_3_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_112_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_5_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_113_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_3_tmp_1 &
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_3_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_3_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_3_nl
      , while_and_112_nl , while_and_113_nl});
  assign input_mem_banks_bank_a_nand_4_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_6_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_4_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_116_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_6_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_117_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_4_tmp_1 &
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_4_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_4_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_4_nl
      , while_and_116_nl , while_and_117_nl});
  assign input_mem_banks_bank_a_nand_5_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_7_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_5_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_120_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_7_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_121_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_5_tmp_1 &
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_5_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_5_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_5_nl
      , while_and_120_nl , while_and_121_nl});
  assign input_mem_banks_bank_a_nand_6_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_8_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_6_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_124_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_8_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_125_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_6_tmp_1 &
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_6_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_6_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_6_nl
      , while_and_124_nl , while_and_125_nl});
  assign input_mem_banks_bank_a_nand_7_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_9_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_7_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_128_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_9_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_129_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_7_tmp_1 &
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_7_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_7_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_7_nl
      , while_and_128_nl , while_and_129_nl});
  assign input_mem_banks_bank_a_nand_8_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_10_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_8_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_132_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_10_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_133_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_8_tmp_1 &
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_8_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_8_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_8_nl
      , while_and_132_nl , while_and_133_nl});
  assign input_mem_banks_bank_a_nand_9_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_11_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_9_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_136_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_11_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_137_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_9_tmp_1 &
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_9_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_9_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_9_nl
      , while_and_136_nl , while_and_137_nl});
  assign input_mem_banks_bank_a_nand_10_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_12_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_10_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_140_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_12_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_141_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_10_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_10_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_10_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_10_nl
      , while_and_140_nl , while_and_141_nl});
  assign input_mem_banks_bank_a_nand_11_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_13_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_11_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_144_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_13_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_145_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_11_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_11_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_11_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_11_nl
      , while_and_144_nl , while_and_145_nl});
  assign input_mem_banks_bank_a_nand_12_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_14_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_12_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_148_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_14_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_149_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_12_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_12_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_12_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_12_nl
      , while_and_148_nl , while_and_149_nl});
  assign input_mem_banks_bank_a_nand_13_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_15_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_13_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_152_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_15_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_153_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_13_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_13_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_13_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_13_nl
      , while_and_152_nl , while_and_153_nl});
  assign input_mem_banks_bank_a_nand_14_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_16_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_14_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_156_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_16_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_157_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_14_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_14_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_14_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_14_nl
      , while_and_156_nl , while_and_157_nl});
  assign input_mem_banks_bank_a_nand_15_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_17_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_15_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_160_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_17_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_161_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_15_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_15_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_15_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_15_nl
      , while_and_160_nl , while_and_161_nl});
  assign input_mem_banks_bank_a_nand_16_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_18_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_16_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_164_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_18_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_165_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_16_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_16_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_16_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_16_nl
      , while_and_164_nl , while_and_165_nl});
  assign input_mem_banks_bank_a_nand_17_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_19_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_17_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_168_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_19_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_169_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_17_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_17_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_17_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_17_nl
      , while_and_168_nl , while_and_169_nl});
  assign input_mem_banks_bank_a_nand_18_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_20_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_18_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_172_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_20_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_173_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_18_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_18_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_18_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_18_nl
      , while_and_172_nl , while_and_173_nl});
  assign input_mem_banks_bank_a_nand_19_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_21_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_19_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_176_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_21_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_177_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_19_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_19_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_19_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_19_nl
      , while_and_176_nl , while_and_177_nl});
  assign input_mem_banks_bank_a_nand_20_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_22_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_20_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_180_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_22_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_181_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_20_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_20_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_20_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_20_nl
      , while_and_180_nl , while_and_181_nl});
  assign input_mem_banks_bank_a_nand_21_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_23_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_21_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_184_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_23_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_185_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_21_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_21_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_21_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_21_nl
      , while_and_184_nl , while_and_185_nl});
  assign input_mem_banks_bank_a_nand_22_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_24_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_22_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_188_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_24_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_189_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_22_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_22_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_22_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_22_nl
      , while_and_188_nl , while_and_189_nl});
  assign input_mem_banks_bank_a_nand_23_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_25_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_23_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_192_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_25_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_193_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_23_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_23_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_23_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_23_nl
      , while_and_192_nl , while_and_193_nl});
  assign input_mem_banks_bank_a_nand_24_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_26_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_24_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_196_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_26_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_197_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_24_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_24_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_24_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_24_nl
      , while_and_196_nl , while_and_197_nl});
  assign input_mem_banks_bank_a_nand_25_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_27_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_25_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_200_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_27_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_201_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_25_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_25_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_25_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_25_nl
      , while_and_200_nl , while_and_201_nl});
  assign input_mem_banks_bank_a_nand_26_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_28_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_26_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_204_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_28_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_205_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_26_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_26_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_26_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_26_nl
      , while_and_204_nl , while_and_205_nl});
  assign input_mem_banks_bank_a_nand_27_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_29_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_27_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_208_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_29_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_209_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_27_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_27_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_27_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_27_nl
      , while_and_208_nl , while_and_209_nl});
  assign input_mem_banks_bank_a_nand_28_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_30_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_28_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_212_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_30_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_213_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_28_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_28_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_28_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_28_nl
      , while_and_212_nl , while_and_213_nl});
  assign input_mem_banks_bank_a_nand_29_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_31_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_29_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_216_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_31_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_217_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_29_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_29_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_29_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_29_nl
      , while_and_216_nl , while_and_217_nl});
  assign input_mem_banks_bank_a_nand_30_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_32_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_30_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_220_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_32_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_221_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_30_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_30_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_30_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_30_nl
      , while_and_220_nl , while_and_221_nl});
  assign input_mem_banks_bank_a_nand_31_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_33_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_31_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_224_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_33_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_225_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_31_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_31_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_31_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_31_nl
      , while_and_224_nl , while_and_225_nl});
  assign input_mem_banks_bank_a_nand_32_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_34_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_32_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_228_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_34_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_229_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_32_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_32_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_32_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_32_nl
      , while_and_228_nl , while_and_229_nl});
  assign input_mem_banks_bank_a_nand_33_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_35_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_33_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_232_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_35_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_233_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_33_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_33_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_33_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_33_nl
      , while_and_232_nl , while_and_233_nl});
  assign input_mem_banks_bank_a_nand_34_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_36_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_34_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_236_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_36_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_237_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_34_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_34_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_34_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_34_nl
      , while_and_236_nl , while_and_237_nl});
  assign input_mem_banks_bank_a_nand_35_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_37_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_35_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_240_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_37_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_241_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_35_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_35_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_35_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_35_nl
      , while_and_240_nl , while_and_241_nl});
  assign input_mem_banks_bank_a_nand_36_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_38_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_36_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_244_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_38_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_245_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_36_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_36_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_36_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_36_nl
      , while_and_244_nl , while_and_245_nl});
  assign input_mem_banks_bank_a_nand_37_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_39_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_37_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_248_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_39_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_249_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_37_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_37_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_37_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_37_nl
      , while_and_248_nl , while_and_249_nl});
  assign input_mem_banks_bank_a_nand_38_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_40_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_38_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_252_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_40_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_253_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_38_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_38_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_38_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_38_nl
      , while_and_252_nl , while_and_253_nl});
  assign input_mem_banks_bank_a_nand_39_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_41_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_39_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_256_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_41_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_257_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_39_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_39_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_39_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_39_nl
      , while_and_256_nl , while_and_257_nl});
  assign input_mem_banks_bank_a_nand_40_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_42_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_40_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_260_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_42_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_261_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_40_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_40_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_40_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_40_nl
      , while_and_260_nl , while_and_261_nl});
  assign input_mem_banks_bank_a_nand_41_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_43_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_41_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_264_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_43_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_265_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_41_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_41_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_41_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_41_nl
      , while_and_264_nl , while_and_265_nl});
  assign input_mem_banks_bank_a_nand_42_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_44_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_42_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_268_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_44_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_269_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_42_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_42_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_42_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_42_nl
      , while_and_268_nl , while_and_269_nl});
  assign input_mem_banks_bank_a_nand_43_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_45_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_43_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_272_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_45_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_273_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_43_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_43_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_43_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_43_nl
      , while_and_272_nl , while_and_273_nl});
  assign input_mem_banks_bank_a_nand_44_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_46_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_44_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_276_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_46_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_277_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_44_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_44_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_44_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_44_nl
      , while_and_276_nl , while_and_277_nl});
  assign input_mem_banks_bank_a_nand_45_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_47_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_45_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_280_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_47_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_281_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_45_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_45_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_45_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_45_nl
      , while_and_280_nl , while_and_281_nl});
  assign input_mem_banks_bank_a_nand_46_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_48_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_46_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_284_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_48_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_285_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_46_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_46_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_46_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_46_nl
      , while_and_284_nl , while_and_285_nl});
  assign input_mem_banks_bank_a_nand_47_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_49_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_47_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_288_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_49_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_289_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_47_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_47_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_47_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_47_nl
      , while_and_288_nl , while_and_289_nl});
  assign input_mem_banks_bank_a_nand_48_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_50_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_48_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_292_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_50_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_293_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_48_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_48_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_48_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_48_nl
      , while_and_292_nl , while_and_293_nl});
  assign input_mem_banks_bank_a_nand_49_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_51_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_49_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_296_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_51_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_297_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_49_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_49_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_49_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_49_nl
      , while_and_296_nl , while_and_297_nl});
  assign input_mem_banks_bank_a_nand_50_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_52_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_50_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_300_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_52_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_301_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_50_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_50_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_50_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_50_nl
      , while_and_300_nl , while_and_301_nl});
  assign input_mem_banks_bank_a_nand_51_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_53_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_51_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_304_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_53_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_305_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_51_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_51_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_51_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_51_nl
      , while_and_304_nl , while_and_305_nl});
  assign input_mem_banks_bank_a_nand_52_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_54_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_52_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_308_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_54_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_309_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_52_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_52_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_52_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_52_nl
      , while_and_308_nl , while_and_309_nl});
  assign input_mem_banks_bank_a_nand_53_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_55_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_53_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_312_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_55_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_313_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_53_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_53_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_53_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_53_nl
      , while_and_312_nl , while_and_313_nl});
  assign input_mem_banks_bank_a_nand_54_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_56_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_54_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_316_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_56_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_317_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_54_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_54_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_54_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_54_nl
      , while_and_316_nl , while_and_317_nl});
  assign input_mem_banks_bank_a_nand_55_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_57_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_55_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_320_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_57_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_321_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_55_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_55_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_55_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_55_nl
      , while_and_320_nl , while_and_321_nl});
  assign input_mem_banks_bank_a_nand_56_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_58_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_56_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_324_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_58_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_325_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_56_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_56_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_56_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_56_nl
      , while_and_324_nl , while_and_325_nl});
  assign input_mem_banks_bank_a_nand_57_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_59_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_57_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_328_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_59_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_329_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_57_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_57_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_57_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_57_nl
      , while_and_328_nl , while_and_329_nl});
  assign input_mem_banks_bank_a_nand_58_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_60_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_58_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_332_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_60_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_333_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_58_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_58_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_58_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_58_nl
      , while_and_332_nl , while_and_333_nl});
  assign input_mem_banks_bank_a_nand_59_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_61_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_59_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_336_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_61_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_337_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_59_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_59_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_59_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_59_nl
      , while_and_336_nl , while_and_337_nl});
  assign input_mem_banks_bank_a_nand_60_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_62_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_60_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_340_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_62_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_341_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_60_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_60_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_60_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_60_nl
      , while_and_340_nl , while_and_341_nl});
  assign input_mem_banks_bank_a_nand_61_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_63_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_61_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_344_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_63_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_345_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_61_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_61_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_61_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_61_nl
      , while_and_344_nl , while_and_345_nl});
  assign input_mem_banks_bank_a_nand_62_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_64_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_62_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_348_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_64_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_349_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_62_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_62_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_62_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_62_nl
      , while_and_348_nl , while_and_349_nl});
  assign input_mem_banks_bank_a_nand_63_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_65_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_63_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_352_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_65_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_353_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_63_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_63_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_63_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_63_nl
      , while_and_352_nl , while_and_353_nl});
  assign input_mem_banks_bank_a_nand_64_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_66_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_64_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_356_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_66_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_357_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_64_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_64_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_64_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_64_nl
      , while_and_356_nl , while_and_357_nl});
  assign input_mem_banks_bank_a_nand_65_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_67_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_65_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_360_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_67_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_361_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_65_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_65_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_65_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_65_nl
      , while_and_360_nl , while_and_361_nl});
  assign input_mem_banks_bank_a_nand_66_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_68_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_66_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_364_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_68_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_365_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_66_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_66_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_66_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_66_nl
      , while_and_364_nl , while_and_365_nl});
  assign input_mem_banks_bank_a_nand_67_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_69_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_67_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_368_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_69_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_369_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_67_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_67_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_67_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_67_nl
      , while_and_368_nl , while_and_369_nl});
  assign input_mem_banks_bank_a_nand_68_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_70_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_68_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_372_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_70_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_373_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_68_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_68_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_68_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_68_nl
      , while_and_372_nl , while_and_373_nl});
  assign input_mem_banks_bank_a_nand_69_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_71_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_69_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_376_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_71_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_377_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_69_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_69_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_69_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_69_nl
      , while_and_376_nl , while_and_377_nl});
  assign input_mem_banks_bank_a_nand_70_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_72_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_70_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_380_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_72_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_381_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_70_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_70_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_70_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_70_nl
      , while_and_380_nl , while_and_381_nl});
  assign input_mem_banks_bank_a_nand_71_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_73_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_71_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_384_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_73_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_385_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_71_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_71_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_71_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_71_nl
      , while_and_384_nl , while_and_385_nl});
  assign input_mem_banks_bank_a_nand_72_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_74_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_72_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_388_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_74_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_389_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_72_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_72_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_72_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_72_nl
      , while_and_388_nl , while_and_389_nl});
  assign input_mem_banks_bank_a_nand_73_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_75_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_73_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_392_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_75_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_393_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_73_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_73_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_73_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_73_nl
      , while_and_392_nl , while_and_393_nl});
  assign input_mem_banks_bank_a_nand_74_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_76_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_74_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_396_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_76_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_397_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_74_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_74_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_74_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_74_nl
      , while_and_396_nl , while_and_397_nl});
  assign input_mem_banks_bank_a_nand_75_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_77_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_75_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_400_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_77_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_401_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_75_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_75_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_75_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_75_nl
      , while_and_400_nl , while_and_401_nl});
  assign input_mem_banks_bank_a_nand_76_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_78_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_76_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_404_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_78_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_405_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_76_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_76_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_76_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_76_nl
      , while_and_404_nl , while_and_405_nl});
  assign input_mem_banks_bank_a_nand_77_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_79_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_77_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_408_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_79_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_409_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_77_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_77_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_77_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_77_nl
      , while_and_408_nl , while_and_409_nl});
  assign input_mem_banks_bank_a_nand_78_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_80_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_78_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_412_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_80_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_413_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_78_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_78_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_78_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_78_nl
      , while_and_412_nl , while_and_413_nl});
  assign input_mem_banks_bank_a_nand_79_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_81_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_79_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_416_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_81_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_417_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_79_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_79_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_79_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_79_nl
      , while_and_416_nl , while_and_417_nl});
  assign input_mem_banks_bank_a_nand_80_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_82_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_80_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_420_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_82_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_421_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_80_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_80_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_80_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_80_nl
      , while_and_420_nl , while_and_421_nl});
  assign input_mem_banks_bank_a_nand_81_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_83_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_81_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_424_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_83_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_425_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_81_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_81_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_81_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_81_nl
      , while_and_424_nl , while_and_425_nl});
  assign input_mem_banks_bank_a_nand_82_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_84_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_82_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_428_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_84_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_429_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_82_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_82_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_82_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_82_nl
      , while_and_428_nl , while_and_429_nl});
  assign input_mem_banks_bank_a_nand_83_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_85_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_83_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_432_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_85_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_433_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_83_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_83_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_83_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_83_nl
      , while_and_432_nl , while_and_433_nl});
  assign input_mem_banks_bank_a_nand_84_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_86_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_84_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_436_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_86_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_437_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_84_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_84_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_84_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_84_nl
      , while_and_436_nl , while_and_437_nl});
  assign input_mem_banks_bank_a_nand_85_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_87_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_85_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_440_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_87_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_441_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_85_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_85_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_85_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_85_nl
      , while_and_440_nl , while_and_441_nl});
  assign input_mem_banks_bank_a_nand_86_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_88_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_86_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_444_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_88_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_445_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_86_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_86_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_86_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_86_nl
      , while_and_444_nl , while_and_445_nl});
  assign input_mem_banks_bank_a_nand_87_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_89_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_87_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_448_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_89_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_449_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_87_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_87_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_87_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_87_nl
      , while_and_448_nl , while_and_449_nl});
  assign input_mem_banks_bank_a_nand_88_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_90_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_88_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_452_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_90_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_453_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_88_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_88_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_88_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_88_nl
      , while_and_452_nl , while_and_453_nl});
  assign input_mem_banks_bank_a_nand_89_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_91_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_89_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_456_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_91_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_457_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_89_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_89_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_89_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_89_nl
      , while_and_456_nl , while_and_457_nl});
  assign input_mem_banks_bank_a_nand_90_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_92_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_90_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_460_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_92_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_461_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_90_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_90_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_90_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_90_nl
      , while_and_460_nl , while_and_461_nl});
  assign input_mem_banks_bank_a_nand_91_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_93_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_91_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_464_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_93_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_465_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_91_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_91_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_91_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_91_nl
      , while_and_464_nl , while_and_465_nl});
  assign input_mem_banks_bank_a_nand_92_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_94_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_92_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_468_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_94_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_469_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_92_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_92_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_92_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_92_nl
      , while_and_468_nl , while_and_469_nl});
  assign input_mem_banks_bank_a_nand_93_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_95_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_93_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_472_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_95_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_473_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_93_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_93_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_93_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_93_nl
      , while_and_472_nl , while_and_473_nl});
  assign input_mem_banks_bank_a_nand_94_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_96_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_94_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_476_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_96_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_477_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_94_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_94_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_94_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_94_nl
      , while_and_476_nl , while_and_477_nl});
  assign input_mem_banks_bank_a_nand_95_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_97_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_95_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_480_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_97_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_481_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_95_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_95_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_95_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_95_nl
      , while_and_480_nl , while_and_481_nl});
  assign input_mem_banks_bank_a_nand_96_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_98_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_96_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_484_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_98_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_485_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_96_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_96_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_96_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_96_nl
      , while_and_484_nl , while_and_485_nl});
  assign input_mem_banks_bank_a_nand_97_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_99_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_97_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_488_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_99_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_489_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_97_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_97_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_97_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_97_nl
      , while_and_488_nl , while_and_489_nl});
  assign input_mem_banks_bank_a_nand_98_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_100_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_98_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_492_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_100_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_493_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_98_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_98_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_98_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_98_nl
      , while_and_492_nl , while_and_493_nl});
  assign input_mem_banks_bank_a_nand_99_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_101_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_99_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_496_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_101_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_497_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_99_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_99_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_99_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_99_nl
      , while_and_496_nl , while_and_497_nl});
  assign input_mem_banks_bank_a_nand_100_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_102_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_100_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_500_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_102_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_501_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_100_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_100_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_100_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_100_nl
      , while_and_500_nl , while_and_501_nl});
  assign input_mem_banks_bank_a_nand_101_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_103_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_101_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_504_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_103_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_505_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_101_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_101_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_101_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_101_nl
      , while_and_504_nl , while_and_505_nl});
  assign input_mem_banks_bank_a_nand_102_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_104_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_102_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_508_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_104_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_509_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_102_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_102_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_102_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_102_nl
      , while_and_508_nl , while_and_509_nl});
  assign input_mem_banks_bank_a_nand_103_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_105_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_103_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_512_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_105_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_513_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_103_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_103_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_103_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_103_nl
      , while_and_512_nl , while_and_513_nl});
  assign input_mem_banks_bank_a_nand_104_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_106_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_104_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_516_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_106_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_517_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_104_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_104_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_104_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_104_nl
      , while_and_516_nl , while_and_517_nl});
  assign input_mem_banks_bank_a_nand_105_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_107_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_105_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_520_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_107_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_521_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_105_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_105_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_105_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_105_nl
      , while_and_520_nl , while_and_521_nl});
  assign input_mem_banks_bank_a_nand_106_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_108_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_106_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_524_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_108_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_525_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_106_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_106_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_106_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_106_nl
      , while_and_524_nl , while_and_525_nl});
  assign input_mem_banks_bank_a_nand_107_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_109_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_107_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_528_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_109_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_529_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_107_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_107_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_107_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_107_nl
      , while_and_528_nl , while_and_529_nl});
  assign input_mem_banks_bank_a_nand_108_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_110_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_108_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_532_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_110_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_533_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_108_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_108_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_108_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_108_nl
      , while_and_532_nl , while_and_533_nl});
  assign input_mem_banks_bank_a_nand_109_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_111_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_109_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_536_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_111_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_537_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_109_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_109_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_109_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_109_nl
      , while_and_536_nl , while_and_537_nl});
  assign input_mem_banks_bank_a_nand_110_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_112_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_110_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_540_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_112_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_541_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_110_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_110_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_110_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_110_nl
      , while_and_540_nl , while_and_541_nl});
  assign input_mem_banks_bank_a_nand_111_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_113_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_111_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_544_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_113_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_545_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_111_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_111_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_111_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_111_nl
      , while_and_544_nl , while_and_545_nl});
  assign input_mem_banks_bank_a_nand_112_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_114_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_112_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_548_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_114_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_549_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_112_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_112_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_112_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_112_nl
      , while_and_548_nl , while_and_549_nl});
  assign input_mem_banks_bank_a_nand_113_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_115_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_113_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_552_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_115_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_553_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_113_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_113_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_113_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_113_nl
      , while_and_552_nl , while_and_553_nl});
  assign input_mem_banks_bank_a_nand_114_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_116_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_114_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_556_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_116_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_557_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_114_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_114_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_114_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_114_nl
      , while_and_556_nl , while_and_557_nl});
  assign input_mem_banks_bank_a_nand_115_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_117_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_115_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_560_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_117_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_561_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_115_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_115_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_115_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_115_nl
      , while_and_560_nl , while_and_561_nl});
  assign input_mem_banks_bank_a_nand_116_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_118_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_116_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_564_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_118_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_565_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_116_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_116_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_116_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_116_nl
      , while_and_564_nl , while_and_565_nl});
  assign input_mem_banks_bank_a_nand_117_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_119_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_117_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_568_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_119_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_569_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_117_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_117_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_117_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_117_nl
      , while_and_568_nl , while_and_569_nl});
  assign input_mem_banks_bank_a_nand_118_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_120_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_118_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_572_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_120_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_573_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_118_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_118_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_118_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_118_nl
      , while_and_572_nl , while_and_573_nl});
  assign input_mem_banks_bank_a_nand_119_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_121_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_119_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_576_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_121_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_577_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_119_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_119_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_119_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_119_nl
      , while_and_576_nl , while_and_577_nl});
  assign input_mem_banks_bank_a_nand_120_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_122_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_120_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_580_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_122_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_581_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_120_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_120_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_120_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_120_nl
      , while_and_580_nl , while_and_581_nl});
  assign input_mem_banks_bank_a_nand_121_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_123_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_121_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_584_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_123_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_585_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_121_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_121_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_121_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_121_nl
      , while_and_584_nl , while_and_585_nl});
  assign input_mem_banks_bank_a_nand_122_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_124_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_122_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_588_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_124_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_589_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_122_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_122_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_122_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_122_nl
      , while_and_588_nl , while_and_589_nl});
  assign input_mem_banks_bank_a_nand_123_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_125_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_123_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_592_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_125_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_593_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_123_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_123_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_123_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_123_nl
      , while_and_592_nl , while_and_593_nl});
  assign input_mem_banks_bank_a_nand_124_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_126_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_124_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_596_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_126_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_597_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_124_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_124_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_124_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_124_nl
      , while_and_596_nl , while_and_597_nl});
  assign input_mem_banks_bank_a_nand_125_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_127_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_125_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_600_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_127_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_601_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_125_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_125_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_125_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_125_nl
      , while_and_600_nl , while_and_601_nl});
  assign input_mem_banks_bank_a_nand_126_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_128_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_126_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_604_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_128_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_605_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_126_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_126_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_126_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_126_nl
      , while_and_604_nl , while_and_605_nl});
  assign input_mem_banks_bank_a_nand_127_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_129_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_127_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_608_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_129_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_609_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_127_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_127_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_127_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_127_nl
      , while_and_608_nl , while_and_609_nl});
  assign input_mem_banks_bank_a_nand_128_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_130_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_128_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_612_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_130_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_613_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_128_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_128_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_128_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_128_nl
      , while_and_612_nl , while_and_613_nl});
  assign input_mem_banks_bank_a_nand_129_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_131_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_129_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_616_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_131_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_617_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_129_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_129_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_129_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_129_nl
      , while_and_616_nl , while_and_617_nl});
  assign input_mem_banks_bank_a_nand_130_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_132_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_130_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_620_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_132_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_621_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_130_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_130_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_130_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_130_nl
      , while_and_620_nl , while_and_621_nl});
  assign input_mem_banks_bank_a_nand_131_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_133_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_131_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_624_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_133_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_625_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_131_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_131_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_131_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_131_nl
      , while_and_624_nl , while_and_625_nl});
  assign input_mem_banks_bank_a_nand_132_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_134_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_132_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_628_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_134_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_629_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_132_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_132_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_132_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_132_nl
      , while_and_628_nl , while_and_629_nl});
  assign input_mem_banks_bank_a_nand_133_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_135_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_133_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_632_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_135_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_633_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_133_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_133_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_133_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_133_nl
      , while_and_632_nl , while_and_633_nl});
  assign input_mem_banks_bank_a_nand_134_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_136_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_134_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_636_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_136_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_637_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_134_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_134_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_134_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_134_nl
      , while_and_636_nl , while_and_637_nl});
  assign input_mem_banks_bank_a_nand_135_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_137_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_135_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_640_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_137_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_641_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_135_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_135_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_135_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_135_nl
      , while_and_640_nl , while_and_641_nl});
  assign input_mem_banks_bank_a_nand_136_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_138_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_136_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_644_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_138_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_645_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_136_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_136_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_136_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_136_nl
      , while_and_644_nl , while_and_645_nl});
  assign input_mem_banks_bank_a_nand_137_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_139_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_137_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_648_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_139_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_649_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_137_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_137_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_137_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_137_nl
      , while_and_648_nl , while_and_649_nl});
  assign input_mem_banks_bank_a_nand_138_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_140_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_138_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_652_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_140_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_653_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_138_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_138_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_138_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_138_nl
      , while_and_652_nl , while_and_653_nl});
  assign input_mem_banks_bank_a_nand_139_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_141_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_139_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_656_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_141_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_657_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_139_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_139_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_139_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_139_nl
      , while_and_656_nl , while_and_657_nl});
  assign input_mem_banks_bank_a_nand_140_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_142_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_140_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_660_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_142_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_661_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_140_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_140_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_140_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_140_nl
      , while_and_660_nl , while_and_661_nl});
  assign input_mem_banks_bank_a_nand_141_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_143_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_141_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_664_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_143_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_665_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_141_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_141_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_141_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_141_nl
      , while_and_664_nl , while_and_665_nl});
  assign input_mem_banks_bank_a_nand_142_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_144_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_142_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_668_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_144_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_669_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_142_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_142_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_142_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_142_nl
      , while_and_668_nl , while_and_669_nl});
  assign input_mem_banks_bank_a_nand_143_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_145_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_143_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_672_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_145_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_673_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_143_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_143_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_143_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_143_nl
      , while_and_672_nl , while_and_673_nl});
  assign input_mem_banks_bank_a_nand_144_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_146_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_144_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_676_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_146_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_677_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_144_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_144_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_144_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_144_nl
      , while_and_676_nl , while_and_677_nl});
  assign input_mem_banks_bank_a_nand_145_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_147_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_145_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_680_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_147_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_681_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_145_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_145_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_145_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_145_nl
      , while_and_680_nl , while_and_681_nl});
  assign input_mem_banks_bank_a_nand_146_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_148_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_146_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_684_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_148_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_685_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_146_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_146_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_146_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_146_nl
      , while_and_684_nl , while_and_685_nl});
  assign input_mem_banks_bank_a_nand_147_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_149_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_147_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_688_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_149_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_689_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_147_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_147_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_147_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_147_nl
      , while_and_688_nl , while_and_689_nl});
  assign input_mem_banks_bank_a_nand_148_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_150_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_148_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_692_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_150_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_693_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_148_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_148_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_148_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_148_nl
      , while_and_692_nl , while_and_693_nl});
  assign input_mem_banks_bank_a_nand_149_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_151_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_149_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_696_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_151_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_697_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_149_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_149_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_149_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_149_nl
      , while_and_696_nl , while_and_697_nl});
  assign input_mem_banks_bank_a_nand_150_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_152_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_150_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_700_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_152_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_701_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_150_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_150_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_150_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_150_nl
      , while_and_700_nl , while_and_701_nl});
  assign input_mem_banks_bank_a_nand_151_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_153_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_151_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_704_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_153_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_705_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_151_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_151_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_151_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_151_nl
      , while_and_704_nl , while_and_705_nl});
  assign input_mem_banks_bank_a_nand_152_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_154_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_152_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_708_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_154_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_709_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_152_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_152_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_152_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_152_nl
      , while_and_708_nl , while_and_709_nl});
  assign input_mem_banks_bank_a_nand_153_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_155_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_153_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_712_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_155_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_713_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_153_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_153_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_153_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_153_nl
      , while_and_712_nl , while_and_713_nl});
  assign input_mem_banks_bank_a_nand_154_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_156_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_154_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_716_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_156_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_717_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_154_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_154_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_154_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_154_nl
      , while_and_716_nl , while_and_717_nl});
  assign input_mem_banks_bank_a_nand_155_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_157_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_155_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_720_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_157_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_721_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_155_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_155_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_155_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_155_nl
      , while_and_720_nl , while_and_721_nl});
  assign input_mem_banks_bank_a_nand_156_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_158_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_156_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_724_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_158_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_725_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_156_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_156_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_156_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_156_nl
      , while_and_724_nl , while_and_725_nl});
  assign input_mem_banks_bank_a_nand_157_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_159_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_157_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_728_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_159_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_729_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_157_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_157_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_157_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_157_nl
      , while_and_728_nl , while_and_729_nl});
  assign input_mem_banks_bank_a_nand_158_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_160_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_158_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_732_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_160_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_733_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_158_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_158_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_158_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_158_nl
      , while_and_732_nl , while_and_733_nl});
  assign input_mem_banks_bank_a_nand_159_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_161_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_159_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_736_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_161_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_737_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_159_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_159_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_159_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_159_nl
      , while_and_736_nl , while_and_737_nl});
  assign input_mem_banks_bank_a_nand_160_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_162_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_160_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_740_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_162_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_741_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_160_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_160_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_160_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_160_nl
      , while_and_740_nl , while_and_741_nl});
  assign input_mem_banks_bank_a_nand_161_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_163_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_161_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_744_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_163_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_745_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_161_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_161_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_161_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_161_nl
      , while_and_744_nl , while_and_745_nl});
  assign input_mem_banks_bank_a_nand_162_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_164_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_162_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_748_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_164_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_749_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_162_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_162_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_162_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_162_nl
      , while_and_748_nl , while_and_749_nl});
  assign input_mem_banks_bank_a_nand_163_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_165_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_163_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_752_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_165_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_753_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_163_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_163_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_163_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_163_nl
      , while_and_752_nl , while_and_753_nl});
  assign input_mem_banks_bank_a_nand_164_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_166_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_164_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_756_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_166_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_757_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_164_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_164_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_164_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_164_nl
      , while_and_756_nl , while_and_757_nl});
  assign input_mem_banks_bank_a_nand_165_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_167_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_165_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_760_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_167_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_761_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_165_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_165_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_165_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_165_nl
      , while_and_760_nl , while_and_761_nl});
  assign input_mem_banks_bank_a_nand_166_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_168_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_166_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_764_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_168_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_765_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_166_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_166_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_166_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_166_nl
      , while_and_764_nl , while_and_765_nl});
  assign input_mem_banks_bank_a_nand_167_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_169_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_167_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_768_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_169_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_769_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_167_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_167_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_167_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_167_nl
      , while_and_768_nl , while_and_769_nl});
  assign input_mem_banks_bank_a_nand_168_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_170_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_168_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_772_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_170_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_773_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_168_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_168_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_168_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_168_nl
      , while_and_772_nl , while_and_773_nl});
  assign input_mem_banks_bank_a_nand_169_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_171_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_169_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_776_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_171_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_777_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_169_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_169_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_169_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_169_nl
      , while_and_776_nl , while_and_777_nl});
  assign input_mem_banks_bank_a_nand_170_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_172_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_170_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_780_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_172_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_781_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_170_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_170_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_170_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_170_nl
      , while_and_780_nl , while_and_781_nl});
  assign input_mem_banks_bank_a_nand_171_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_173_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_171_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_784_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_173_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_785_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_171_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_171_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_171_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_171_nl
      , while_and_784_nl , while_and_785_nl});
  assign input_mem_banks_bank_a_nand_172_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_174_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_172_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_788_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_174_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_789_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_172_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_172_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_172_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_172_nl
      , while_and_788_nl , while_and_789_nl});
  assign input_mem_banks_bank_a_nand_173_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_175_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_173_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_792_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_175_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_793_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_173_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_173_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_173_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_173_nl
      , while_and_792_nl , while_and_793_nl});
  assign input_mem_banks_bank_a_nand_174_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_176_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_174_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_796_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_176_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_797_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_174_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_174_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_174_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_174_nl
      , while_and_796_nl , while_and_797_nl});
  assign input_mem_banks_bank_a_nand_175_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_177_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_175_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_800_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_177_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_801_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_175_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_175_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_175_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_175_nl
      , while_and_800_nl , while_and_801_nl});
  assign input_mem_banks_bank_a_nand_176_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_178_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_176_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_804_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_178_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_805_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_176_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_176_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_176_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_176_nl
      , while_and_804_nl , while_and_805_nl});
  assign input_mem_banks_bank_a_nand_177_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_179_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_177_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_808_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_179_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_809_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_177_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_177_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_177_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_177_nl
      , while_and_808_nl , while_and_809_nl});
  assign input_mem_banks_bank_a_nand_178_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_180_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_178_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_812_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_180_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_813_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_178_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_178_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_178_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_178_nl
      , while_and_812_nl , while_and_813_nl});
  assign input_mem_banks_bank_a_nand_179_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_181_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_179_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_816_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_181_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_817_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_179_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_179_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_179_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_179_nl
      , while_and_816_nl , while_and_817_nl});
  assign input_mem_banks_bank_a_nand_180_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_182_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_180_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_820_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_182_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_821_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_180_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_180_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_180_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_180_nl
      , while_and_820_nl , while_and_821_nl});
  assign input_mem_banks_bank_a_nand_181_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_183_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_181_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_824_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_183_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_825_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_181_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_181_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_181_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_181_nl
      , while_and_824_nl , while_and_825_nl});
  assign input_mem_banks_bank_a_nand_182_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_184_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_182_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_828_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_184_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_829_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_182_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_182_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_182_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_182_nl
      , while_and_828_nl , while_and_829_nl});
  assign input_mem_banks_bank_a_nand_183_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_185_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_183_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_832_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_185_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_833_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_183_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_183_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_183_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_183_nl
      , while_and_832_nl , while_and_833_nl});
  assign input_mem_banks_bank_a_nand_184_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_186_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_184_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_836_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_186_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_837_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_184_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_184_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_184_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_184_nl
      , while_and_836_nl , while_and_837_nl});
  assign input_mem_banks_bank_a_nand_185_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_187_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_185_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_840_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_187_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_841_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_185_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_185_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_185_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_185_nl
      , while_and_840_nl , while_and_841_nl});
  assign input_mem_banks_bank_a_nand_186_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_188_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_186_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_844_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_188_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_845_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_186_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_186_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_186_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_186_nl
      , while_and_844_nl , while_and_845_nl});
  assign input_mem_banks_bank_a_nand_187_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_189_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_187_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_848_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_189_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_849_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_187_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_187_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_187_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_187_nl
      , while_and_848_nl , while_and_849_nl});
  assign input_mem_banks_bank_a_nand_188_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_190_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_188_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_852_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_190_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_853_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_188_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_188_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_188_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_188_nl
      , while_and_852_nl , while_and_853_nl});
  assign input_mem_banks_bank_a_nand_189_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_191_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_189_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_856_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_191_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_857_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_189_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_189_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_189_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_189_nl
      , while_and_856_nl , while_and_857_nl});
  assign input_mem_banks_bank_a_nand_190_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_192_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_190_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_860_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_192_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_861_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_190_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_190_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_190_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_190_nl
      , while_and_860_nl , while_and_861_nl});
  assign input_mem_banks_bank_a_nand_191_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_193_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_191_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_864_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_193_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_865_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_191_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_191_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_191_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_191_nl
      , while_and_864_nl , while_and_865_nl});
  assign input_mem_banks_bank_a_nand_192_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_194_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_192_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_868_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_194_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_869_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_192_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_192_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_192_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_192_nl
      , while_and_868_nl , while_and_869_nl});
  assign input_mem_banks_bank_a_nand_193_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_195_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_193_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_872_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_195_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_873_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_193_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_193_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_193_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_193_nl
      , while_and_872_nl , while_and_873_nl});
  assign input_mem_banks_bank_a_nand_194_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_196_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_194_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_876_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_196_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_877_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_194_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_194_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_194_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_194_nl
      , while_and_876_nl , while_and_877_nl});
  assign input_mem_banks_bank_a_nand_195_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_197_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_195_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_880_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_197_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_881_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_195_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_195_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_195_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_195_nl
      , while_and_880_nl , while_and_881_nl});
  assign input_mem_banks_bank_a_nand_196_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_198_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_196_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_884_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_198_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_885_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_196_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_196_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_196_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_196_nl
      , while_and_884_nl , while_and_885_nl});
  assign input_mem_banks_bank_a_nand_197_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_199_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_197_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_888_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_199_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_889_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_197_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_197_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_197_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_197_nl
      , while_and_888_nl , while_and_889_nl});
  assign input_mem_banks_bank_a_nand_198_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_200_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_198_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_892_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_200_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_893_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_198_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_198_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_198_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_198_nl
      , while_and_892_nl , while_and_893_nl});
  assign input_mem_banks_bank_a_nand_199_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_201_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_199_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_896_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_201_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_897_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_199_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_199_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_199_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_199_nl
      , while_and_896_nl , while_and_897_nl});
  assign input_mem_banks_bank_a_nand_200_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_202_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_200_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_900_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_202_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_901_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_200_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_200_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_200_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_200_nl
      , while_and_900_nl , while_and_901_nl});
  assign input_mem_banks_bank_a_nand_201_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_203_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_201_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_904_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_203_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_905_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_201_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_201_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_201_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_201_nl
      , while_and_904_nl , while_and_905_nl});
  assign input_mem_banks_bank_a_nand_202_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_204_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_202_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_908_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_204_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_909_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_202_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_202_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_202_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_202_nl
      , while_and_908_nl , while_and_909_nl});
  assign input_mem_banks_bank_a_nand_203_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_205_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_203_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_912_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_205_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_913_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_203_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_203_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_203_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_203_nl
      , while_and_912_nl , while_and_913_nl});
  assign input_mem_banks_bank_a_nand_204_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_206_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_204_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_916_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_206_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_917_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_204_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_204_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_204_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_204_nl
      , while_and_916_nl , while_and_917_nl});
  assign input_mem_banks_bank_a_nand_205_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_207_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_205_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_920_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_207_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_921_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_205_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_205_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_205_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_205_nl
      , while_and_920_nl , while_and_921_nl});
  assign input_mem_banks_bank_a_nand_206_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_208_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_206_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_924_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_208_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_925_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_206_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_206_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_206_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_206_nl
      , while_and_924_nl , while_and_925_nl});
  assign input_mem_banks_bank_a_nand_207_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_209_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_207_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_928_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_209_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_929_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_207_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_207_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_207_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_207_nl
      , while_and_928_nl , while_and_929_nl});
  assign input_mem_banks_bank_a_nand_208_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_210_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_208_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_932_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_210_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_933_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_208_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_208_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_208_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_208_nl
      , while_and_932_nl , while_and_933_nl});
  assign input_mem_banks_bank_a_nand_209_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_211_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_209_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_936_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_211_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_937_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_209_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_209_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_209_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_209_nl
      , while_and_936_nl , while_and_937_nl});
  assign input_mem_banks_bank_a_nand_210_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_212_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_210_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_940_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_212_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_941_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_210_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_210_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_210_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_210_nl
      , while_and_940_nl , while_and_941_nl});
  assign input_mem_banks_bank_a_nand_211_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_213_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_211_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_944_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_213_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_945_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_211_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_211_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_211_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_211_nl
      , while_and_944_nl , while_and_945_nl});
  assign input_mem_banks_bank_a_nand_212_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_214_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_212_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_948_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_214_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_949_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_212_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_212_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_212_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_212_nl
      , while_and_948_nl , while_and_949_nl});
  assign input_mem_banks_bank_a_nand_213_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_215_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_213_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_952_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_215_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_953_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_213_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_213_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_213_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_213_nl
      , while_and_952_nl , while_and_953_nl});
  assign input_mem_banks_bank_a_nand_214_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_216_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_214_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_956_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_216_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_957_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_214_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_214_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_214_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_214_nl
      , while_and_956_nl , while_and_957_nl});
  assign input_mem_banks_bank_a_nand_215_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_217_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_215_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_960_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_217_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_961_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_215_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_215_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_215_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_215_nl
      , while_and_960_nl , while_and_961_nl});
  assign input_mem_banks_bank_a_nand_216_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_218_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_216_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_964_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_218_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_965_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_216_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_216_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_216_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_216_nl
      , while_and_964_nl , while_and_965_nl});
  assign input_mem_banks_bank_a_nand_217_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_219_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_217_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_968_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_219_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_969_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_217_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_217_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_217_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_217_nl
      , while_and_968_nl , while_and_969_nl});
  assign input_mem_banks_bank_a_nand_218_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_220_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_218_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_972_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_220_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_973_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_218_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_218_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_218_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_218_nl
      , while_and_972_nl , while_and_973_nl});
  assign input_mem_banks_bank_a_nand_219_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_221_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_219_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_976_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_221_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_977_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_219_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_219_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_219_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_219_nl
      , while_and_976_nl , while_and_977_nl});
  assign input_mem_banks_bank_a_nand_220_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_222_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_220_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_980_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_222_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_981_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_220_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_220_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_220_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_220_nl
      , while_and_980_nl , while_and_981_nl});
  assign input_mem_banks_bank_a_nand_221_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_223_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_221_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_984_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_223_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_985_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_221_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_221_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_221_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_221_nl
      , while_and_984_nl , while_and_985_nl});
  assign input_mem_banks_bank_a_nand_222_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_224_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_222_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_988_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_224_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_989_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_222_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_222_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_222_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_222_nl
      , while_and_988_nl , while_and_989_nl});
  assign input_mem_banks_bank_a_nand_223_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_225_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_223_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_992_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_225_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_993_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_223_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_223_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_223_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_223_nl
      , while_and_992_nl , while_and_993_nl});
  assign input_mem_banks_bank_a_nand_224_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_226_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_224_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_996_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_226_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_997_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_224_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_224_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_224_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_224_nl
      , while_and_996_nl , while_and_997_nl});
  assign input_mem_banks_bank_a_nand_225_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_227_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_225_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_1000_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_227_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_1001_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_225_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_225_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_225_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_225_nl
      , while_and_1000_nl , while_and_1001_nl});
  assign input_mem_banks_bank_a_nand_226_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_228_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_226_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_1004_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_228_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_1005_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_226_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_226_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_226_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_226_nl
      , while_and_1004_nl , while_and_1005_nl});
  assign input_mem_banks_bank_a_nand_227_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_229_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_227_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_1008_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_229_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_1009_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_227_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_227_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_227_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_227_nl
      , while_and_1008_nl , while_and_1009_nl});
  assign input_mem_banks_bank_a_nand_228_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_230_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_228_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_1012_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_230_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_1013_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_228_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_228_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_228_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_228_nl
      , while_and_1012_nl , while_and_1013_nl});
  assign input_mem_banks_bank_a_nand_229_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_231_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_229_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_1016_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_231_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_1017_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_229_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_229_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_229_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_229_nl
      , while_and_1016_nl , while_and_1017_nl});
  assign input_mem_banks_bank_a_nand_230_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_232_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_230_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_1020_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_232_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_1021_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_230_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_230_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_230_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_230_nl
      , while_and_1020_nl , while_and_1021_nl});
  assign input_mem_banks_bank_a_nand_231_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_233_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_231_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_1024_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_233_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_1025_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_231_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_231_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_231_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_231_nl
      , while_and_1024_nl , while_and_1025_nl});
  assign input_mem_banks_bank_a_nand_232_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_234_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_232_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_1028_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_234_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_1029_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_232_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_232_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_232_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_232_nl
      , while_and_1028_nl , while_and_1029_nl});
  assign input_mem_banks_bank_a_nand_233_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_235_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_233_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_1032_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_235_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_1033_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_233_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_233_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_233_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_233_nl
      , while_and_1032_nl , while_and_1033_nl});
  assign input_mem_banks_bank_a_nand_234_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_236_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_234_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_1036_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_236_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_1037_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_234_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_234_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_234_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_234_nl
      , while_and_1036_nl , while_and_1037_nl});
  assign input_mem_banks_bank_a_nand_235_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_237_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_235_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_1040_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_237_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_1041_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_235_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_235_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_235_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_235_nl
      , while_and_1040_nl , while_and_1041_nl});
  assign input_mem_banks_bank_a_nand_236_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_238_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_236_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_1044_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_238_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_1045_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_236_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_236_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_236_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_236_nl
      , while_and_1044_nl , while_and_1045_nl});
  assign input_mem_banks_bank_a_nand_237_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_239_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_237_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_1048_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_239_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_1049_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_237_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_237_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_237_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_237_nl
      , while_and_1048_nl , while_and_1049_nl});
  assign input_mem_banks_bank_a_nand_238_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_240_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_238_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_1052_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_240_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_1053_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_238_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_238_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_238_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_238_nl
      , while_and_1052_nl , while_and_1053_nl});
  assign input_mem_banks_bank_a_nand_239_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_241_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_239_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_1056_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_241_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_1057_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_239_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_239_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_239_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_239_nl
      , while_and_1056_nl , while_and_1057_nl});
  assign input_mem_banks_bank_a_nand_240_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_242_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_240_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_1060_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_242_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_1061_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_240_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_240_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_240_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_240_nl
      , while_and_1060_nl , while_and_1061_nl});
  assign input_mem_banks_bank_a_nand_241_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_243_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_241_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_1064_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_243_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_1065_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_241_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_241_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_241_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_241_nl
      , while_and_1064_nl , while_and_1065_nl});
  assign input_mem_banks_bank_a_nand_242_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_244_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_242_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_1068_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_244_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_1069_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_242_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_242_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_242_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_242_nl
      , while_and_1068_nl , while_and_1069_nl});
  assign input_mem_banks_bank_a_nand_243_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_245_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_243_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_1072_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_245_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_1073_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_243_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_243_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_243_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_243_nl
      , while_and_1072_nl , while_and_1073_nl});
  assign input_mem_banks_bank_a_nand_244_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_246_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_244_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_1076_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_246_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_1077_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_244_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_244_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_244_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_244_nl
      , while_and_1076_nl , while_and_1077_nl});
  assign input_mem_banks_bank_a_nand_245_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_247_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_245_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_1080_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_247_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_1081_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_245_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_245_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_245_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_245_nl
      , while_and_1080_nl , while_and_1081_nl});
  assign input_mem_banks_bank_a_nand_246_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_248_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_246_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_1084_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_248_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_1085_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_246_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_246_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_246_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_246_nl
      , while_and_1084_nl , while_and_1085_nl});
  assign input_mem_banks_bank_a_nand_247_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_249_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_247_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_1088_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_249_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_1089_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_247_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_247_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_247_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_247_nl
      , while_and_1088_nl , while_and_1089_nl});
  assign input_mem_banks_bank_a_nand_248_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_250_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_248_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_1092_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_250_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_1093_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_248_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_248_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_248_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_248_nl
      , while_and_1092_nl , while_and_1093_nl});
  assign input_mem_banks_bank_a_nand_249_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_251_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_249_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_1096_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_251_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_1097_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_249_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_249_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_249_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_249_nl
      , while_and_1096_nl , while_and_1097_nl});
  assign input_mem_banks_bank_a_nand_250_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_252_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_250_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_1100_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_252_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_1101_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_250_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_250_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_250_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_250_nl
      , while_and_1100_nl , while_and_1101_nl});
  assign input_mem_banks_bank_a_nand_251_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_253_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_251_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_1104_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_253_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_1105_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_251_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_251_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_251_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_251_nl
      , while_and_1104_nl , while_and_1105_nl});
  assign input_mem_banks_bank_a_nand_252_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_254_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_252_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_1108_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_254_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_1109_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_252_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_252_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_252_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_252_nl
      , while_and_1108_nl , while_and_1109_nl});
  assign input_mem_banks_bank_a_nand_253_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_255_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_253_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_1112_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_255_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_1113_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_253_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_253_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_253_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_253_nl
      , while_and_1112_nl , while_and_1113_nl});
  assign input_mem_banks_bank_a_nand_254_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_256_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_254_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_1116_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_256_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_1117_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_254_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_254_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_254_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_254_nl
      , while_and_1116_nl , while_and_1117_nl});
  assign input_mem_banks_bank_a_nand_255_nl = ~(while_stage_0_3 & (~((~(input_mem_write_arbxbar_xbar_1_for_3_if_1_and_257_tmp_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      | ((~ input_mem_write_arbxbar_xbar_for_3_if_1_and_255_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))));
  assign while_and_1120_nl = input_mem_write_arbxbar_xbar_1_for_3_if_1_and_257_tmp_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign while_and_1121_nl = input_mem_write_arbxbar_xbar_for_3_if_1_and_255_tmp_1
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign input_mem_banks_bank_a_255_sva_dfm_2_mx1 = MUX1HOT_v_64_3_2(input_mem_banks_bank_a_255_sva_dfm_2,
      input_port_PopNB_mioi_data_data_data_rsc_z_mxwt, rva_in_reg_data_sva_1, {input_mem_banks_bank_a_nand_255_nl
      , while_and_1120_nl , while_and_1121_nl});
  assign accum_vector_data_3_sva_1_load_mx0w0 = PECore_UpdateFSM_switch_lp_equal_tmp_2_1
      | accum_vector_data_3_sva_1_load;
  assign accum_vector_data_2_sva_1_load_mx0w0 = PECore_UpdateFSM_switch_lp_equal_tmp_2_1
      | accum_vector_data_2_sva_1_load;
  assign accum_vector_data_1_sva_1_load_mx0w0 = PECore_UpdateFSM_switch_lp_equal_tmp_2_1
      | accum_vector_data_1_sva_1_load;
  assign accum_vector_data_0_sva_1_load_mx0w0 = PECore_UpdateFSM_switch_lp_equal_tmp_2_1
      | accum_vector_data_0_sva_1_load;
  assign pe_manager_base_input_sva_mx1_7_0 = MUX_v_8_2_2((pe_manager_base_input_sva[7:0]),
      (pe_manager_base_input_sva_dfm_3_1[7:0]), while_stage_0_3);
  assign pe_manager_base_input_sva_mx2 = MUX_v_15_2_2(pe_manager_base_input_sva,
      pe_manager_base_input_sva_dfm_3_1, while_stage_0_3);
  assign accum_vector_data_7_sva_1_load_mx0w1 = PECore_UpdateFSM_switch_lp_equal_tmp_2_1
      | accum_vector_data_7_sva_1_load;
  assign accum_vector_data_5_sva_1_load_mx0w1 = PECore_UpdateFSM_switch_lp_equal_tmp_2_1
      | accum_vector_data_5_sva_1_load;
  assign accum_vector_data_4_sva_1_load_mx0w1 = PECore_UpdateFSM_switch_lp_equal_tmp_2_1
      | accum_vector_data_4_sva_1_load;
  assign PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_mx0w0 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])
      & PECore_DecodeAxiRead_case_4_switch_lp_nor_8_tmp;
  assign PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_mx0w0 = ~(PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_mx0w0
      | and_321_cse);
  assign PECore_RunScale_PECore_RunScale_if_and_1_svs_1 = (state_mux_1_cse[0]) &
      state_0_sva_mx1 & (~ (state_mux_1_cse[1]));
  assign PECore_DecodeAxiRead_switch_lp_nor_tmp_mx0w0 = ~(PECore_DecodeAxiRead_switch_lp_equal_tmp_4
      | PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_and_5 | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0);
  assign PECore_DecodeAxiRead_switch_lp_nor_9_cse_1 = ~(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_9
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_9 | PECore_DecodeAxiRead_switch_lp_nor_tmp_9);
  assign PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_m1c_1 = ~(input_read_req_valid_lpi_1_dfm_1_9
      | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000000
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:8]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:8]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[7:0]),
      {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_12_itm_2});
  assign weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0 = MUX_v_64_2_2(weight_mem_banks_read_1_read_data_7_lpi_1_dfm_1,
      weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d, weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2);
  assign weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0 = MUX_v_56_2_2(weight_mem_banks_read_1_read_data_lpi_1_dfm_1_63_8,
      (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[63:8]), weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_2_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:8]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:8]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[7:0]),
      {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_1_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_1_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[7:0]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[7:0]), BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9,
      {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_1_itm_2});
  assign weight_mem_banks_load_store_1_for_else_else_and_nl = (~(weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2))
      & weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_1_m1c_1
      & weight_mem_banks_load_store_1_for_else_else_and_10_m1c_1;
  assign weight_mem_banks_load_store_1_for_else_else_or_nl = (weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & (~ weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2)
      & weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_1_m1c_1
      & weight_mem_banks_load_store_1_for_else_else_and_10_m1c_1) | (weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_1_m1c_1
      & weight_mem_banks_load_store_1_for_else_else_and_10_m1c_1) | (weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & weight_mem_banks_load_store_1_for_else_else_and_10_m1c_1) | (weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_3_m1c_1);
  assign weight_mem_banks_load_store_1_for_else_else_and_4_nl = weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & (~ weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2)
      & weight_mem_banks_load_store_1_for_else_else_and_10_m1c_1;
  assign weight_mem_banks_load_store_1_for_else_else_and_6_nl = weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & (~ weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2)
      & weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_3_m1c_1;
  assign weight_mem_banks_load_store_1_for_else_else_and_8_nl = weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      & (~ weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2);
  assign BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9 = MUX1HOT_v_8_6_2(BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_8,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_21_itm_1,
      weight_mem_banks_load_store_1_for_3_result_val_Marshall_64U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1,
      weight_mem_banks_load_store_1_for_5_result_val_Marshall_64U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1,
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[7:0]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[7:0]),
      {weight_mem_banks_load_store_1_for_else_else_and_nl , weight_mem_banks_load_store_1_for_else_else_or_nl
      , weight_mem_banks_load_store_1_for_else_else_and_4_nl , weight_mem_banks_load_store_1_for_else_else_and_6_nl
      , weight_mem_banks_load_store_1_for_else_else_and_8_nl , weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_2_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:8]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:8]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[7:0]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_2_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_1_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[7:0]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[7:0]), BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9,
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_2_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_81_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_10_itm_1
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000000
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:8]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:8]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[7:0]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_81_nl , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_118
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_120 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_84_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_122 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_86_itm_2
      , PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4 , PECore_DecodeAxiRead_switch_lp_equal_tmp_2_5});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_89_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_11_itm_1
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000001
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[7:0]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[7:0]), BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9,
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_89_nl , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_118
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_120 , PECore_DecodeAxiRead_switch_lp_equal_tmp_3_5
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_122 , PECore_DecodeAxiRead_switch_lp_nor_tmp_5
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_95_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_124});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000000
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[15:8]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15:8]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15:8]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15:8]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[7:0]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_100 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_60_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_62_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000001
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[7:0]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[7:0]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[7:0]), BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9,
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_98 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_60_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_62_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_cse = ~((reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[2:1]!=2'b00));
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1 = (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[0])
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_cse & weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 = (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1])
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_1_cse & weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 = (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[2])
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_2_cse & weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1 = (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse==3'b111)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  assign weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_1_m1c_1
      = ~(weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2);
  assign weight_mem_banks_load_store_1_for_else_else_and_10_m1c_1 = (~(weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2))
      & weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_3_m1c_1;
  assign weight_mem_banks_load_store_1_for_else_else_weight_mem_banks_load_store_1_for_else_else_nor_3_m1c_1
      = ~(weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_8_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_13_sva_1 & (~ Arbiter_8U_Roundrobin_pick_1_priority_14_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_nl
      = (~ operator_2_false_3_operator_2_false_3_or_mdf_sva_1) & not_tmp_469;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_1_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_sva_1 & not_tmp_469;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_nl
      = ~(operator_2_false_4_operator_2_false_4_or_mdf_sva_1 | mux_306_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_3_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_sva_1 & (~ mux_306_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_4_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_sva_1) & and_dcpl_625;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_5_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_sva_1 & and_dcpl_625;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_8_nl,
      Arbiter_8U_Roundrobin_pick_1_priority_9_sva_1, Arbiter_8U_Roundrobin_pick_1_priority_11_sva_1,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[7]),
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]),
      {mux_tmp_280 , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_1_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_3_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_4_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_5_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_1_priority_14_sva_1, operator_2_false_3_operator_2_false_3_or_mdf_sva_1,
      operator_2_false_4_operator_2_false_4_or_mdf_sva_1, operator_2_false_5_operator_2_false_5_or_mdf_sva_1,
      {mux_tmp_280 , not_tmp_469 , (~ mux_306_itm) , and_dcpl_625});
  assign weight_mem_read_arbxbar_xbar_1_for_3_8_operator_4_false_2_operator_4_false_2_or_nl
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_8_operator_3_false_1_operator_3_false_1_or_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_14_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_13_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_12_sva_1;
  assign mux_316_nl = MUX_s_1_2_2(mux_tmp_295, mux_tmp_294, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]);
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_8_operator_4_false_2_operator_4_false_2_or_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_8_operator_3_false_1_operator_3_false_1_or_nl,
      mux_316_nl);
  assign Arbiter_8U_Roundrobin_pick_1_priority_9_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_2_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_11_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_4_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]);
  assign operator_2_false_3_operator_2_false_3_or_mdf_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_11_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_10_sva_1;
  assign Arbiter_8U_Roundrobin_pick_1_priority_10_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_3_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_13_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_6_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_14_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_7_sva_mx0
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_12_sva_1 = weight_mem_read_arbxbar_arbiters_next_7_5_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_9_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_13_7_sva_1 & (~ Arbiter_8U_Roundrobin_pick_1_priority_14_7_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_1_nl
      = ~(operator_2_false_3_operator_2_false_3_or_mdf_7_sva_1 | mux_330_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_7_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_7_sva_1 & (~ mux_330_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_2_nl
      = ~(operator_2_false_4_operator_2_false_4_or_mdf_7_sva_1 | mux_343_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_9_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_7_sva_1 & (~ mux_343_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_10_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_7_sva_1) & and_dcpl_626;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_11_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_7_sva_1 & and_dcpl_626;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_7_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_9_nl,
      Arbiter_8U_Roundrobin_pick_1_priority_9_7_sva_1, Arbiter_8U_Roundrobin_pick_1_priority_11_7_sva_1,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[6]),
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]),
      {mux_tmp_319 , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_1_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_7_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_2_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_9_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_10_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_11_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_7_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_1_priority_14_7_sva_1, operator_2_false_3_operator_2_false_3_or_mdf_7_sva_1,
      operator_2_false_4_operator_2_false_4_or_mdf_7_sva_1, operator_2_false_5_operator_2_false_5_or_mdf_7_sva_1,
      {mux_tmp_319 , (~ mux_330_itm) , (~ mux_343_itm) , and_dcpl_626});
  assign weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_2_operator_4_false_2_or_nl
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_7_operator_3_false_1_operator_3_false_1_or_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_14_7_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_13_7_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_12_7_sva_1;
  assign mux_353_nl = MUX_s_1_2_2(mux_tmp_332, mux_tmp_330, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]);
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_2_operator_4_false_2_or_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_7_operator_3_false_1_operator_3_false_1_or_nl,
      mux_353_nl);
  assign Arbiter_8U_Roundrobin_pick_1_priority_9_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_2_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_11_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_4_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]);
  assign operator_2_false_3_operator_2_false_3_or_mdf_7_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_11_7_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_10_7_sva_1;
  assign Arbiter_8U_Roundrobin_pick_1_priority_10_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_3_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_13_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_6_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_14_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_7_sva_mx0
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_12_7_sva_1 = weight_mem_read_arbxbar_arbiters_next_6_5_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_7_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_7_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_10_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_13_6_sva_1 & (~ weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_12_nl
      = (~ operator_2_false_3_operator_2_false_3_or_mdf_6_sva_1) & and_dcpl_629;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_13_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_6_sva_1 & and_dcpl_629;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_14_nl
      = (~ operator_2_false_4_operator_2_false_4_or_mdf_6_sva_1) & and_dcpl_632;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_15_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_6_sva_1 & and_dcpl_632;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_16_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_6_sva_1) & and_dcpl_639;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_17_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_6_sva_1 & and_dcpl_639;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_6_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_10_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_3_tmp,
      Arbiter_8U_Roundrobin_pick_1_priority_11_6_sva_1, (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]),
      (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[5]), (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[5]),
      (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5]), {or_dcpl_677 , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_12_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_13_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_14_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_15_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_16_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_17_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_6_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp,
      operator_2_false_3_operator_2_false_3_or_mdf_6_sva_1, operator_2_false_4_operator_2_false_4_or_mdf_6_sva_1,
      operator_2_false_5_operator_2_false_5_or_mdf_6_sva_1, {or_dcpl_677 , and_dcpl_629
      , and_dcpl_632 , and_dcpl_639});
  assign weight_mem_read_arbxbar_xbar_1_for_3_6_operator_3_false_1_operator_3_false_1_or_nl
      = weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp
      | Arbiter_8U_Roundrobin_pick_1_priority_13_6_sva_1 | weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp;
  assign weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_2_operator_4_false_2_or_nl
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5]);
  assign and_667_nl = (~ mux_tmp_362) & and_dcpl_631;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_6_operator_3_false_1_operator_3_false_1_or_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_2_operator_4_false_2_or_nl,
      and_667_nl);
  assign weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_3_tmp
      = weight_mem_read_arbxbar_arbiters_next_5_2_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[5]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_11_6_sva_1 = weight_mem_read_arbxbar_arbiters_next_5_4_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5]);
  assign operator_2_false_3_operator_2_false_3_or_mdf_6_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_11_6_sva_1
      | (weight_mem_read_arbxbar_arbiters_next_5_3_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5]));
  assign Arbiter_8U_Roundrobin_pick_1_priority_13_6_sva_1 = weight_mem_read_arbxbar_arbiters_next_5_6_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp
      = weight_mem_read_arbxbar_arbiters_next_5_7_sva_mx0 & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp
      = weight_mem_read_arbxbar_arbiters_next_5_5_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_6_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_6_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5]);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_11_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_13_5_sva_1 & (~ Arbiter_8U_Roundrobin_pick_1_priority_14_5_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_3_nl
      = ~(operator_2_false_3_operator_2_false_3_or_mdf_5_sva_1 | mux_373_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_19_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_5_sva_1 & (~ mux_373_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_4_nl
      = ~(operator_2_false_4_operator_2_false_4_or_mdf_5_sva_1 | mux_380_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_21_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_5_sva_1 & (~ mux_380_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_22_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_5_sva_1) & and_dcpl_641;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_23_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_5_sva_1 & and_dcpl_641;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_5_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_11_nl,
      Arbiter_8U_Roundrobin_pick_1_priority_9_5_sva_1, Arbiter_8U_Roundrobin_pick_1_priority_11_5_sva_1,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[4]),
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[4]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4]),
      {mux_tmp_366 , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_3_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_19_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_4_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_21_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_22_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_23_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_5_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_1_priority_14_5_sva_1, operator_2_false_3_operator_2_false_3_or_mdf_5_sva_1,
      operator_2_false_4_operator_2_false_4_or_mdf_5_sva_1, operator_2_false_5_operator_2_false_5_or_mdf_5_sva_1,
      {mux_tmp_366 , (~ mux_373_itm) , (~ mux_380_itm) , and_dcpl_641});
  assign weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_2_operator_4_false_2_or_nl
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_5_operator_3_false_1_operator_3_false_1_or_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_14_5_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_13_5_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_12_5_sva_1;
  assign mux_388_nl = MUX_s_1_2_2(mux_tmp_371, mux_tmp_370, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4]);
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_2_operator_4_false_2_or_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_5_operator_3_false_1_operator_3_false_1_or_nl,
      mux_388_nl);
  assign Arbiter_8U_Roundrobin_pick_1_priority_9_5_sva_1 = weight_mem_read_arbxbar_arbiters_next_4_2_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[4]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_11_5_sva_1 = weight_mem_read_arbxbar_arbiters_next_4_4_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4]);
  assign operator_2_false_3_operator_2_false_3_or_mdf_5_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_11_5_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_10_5_sva_1;
  assign Arbiter_8U_Roundrobin_pick_1_priority_10_5_sva_1 = weight_mem_read_arbxbar_arbiters_next_4_3_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_13_5_sva_1 = weight_mem_read_arbxbar_arbiters_next_4_6_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_14_5_sva_1 = weight_mem_read_arbxbar_arbiters_next_4_7_sva_mx0
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_12_5_sva_1 = weight_mem_read_arbxbar_arbiters_next_4_5_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_5_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_5_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4]);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_12_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_13_4_sva_1 & (~ Arbiter_8U_Roundrobin_pick_1_priority_14_4_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_5_nl
      = ~(operator_2_false_3_operator_2_false_3_or_mdf_4_sva_1 | mux_394_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_25_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_4_sva_1 & (~ mux_394_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_6_nl
      = ~(operator_2_false_4_operator_2_false_4_or_mdf_4_sva_1 | mux_401_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_27_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_4_sva_1 & (~ mux_401_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_28_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_4_sva_1) & and_dcpl_642;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_29_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_4_sva_1 & and_dcpl_642;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_4_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_12_nl,
      Arbiter_8U_Roundrobin_pick_1_priority_9_4_sva_1, Arbiter_8U_Roundrobin_pick_1_priority_11_4_sva_1,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[3]),
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[3]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[3]),
      {mux_tmp_387 , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_5_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_25_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_6_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_27_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_28_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_29_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_4_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_1_priority_14_4_sva_1, operator_2_false_3_operator_2_false_3_or_mdf_4_sva_1,
      operator_2_false_4_operator_2_false_4_or_mdf_4_sva_1, operator_2_false_5_operator_2_false_5_or_mdf_4_sva_1,
      {mux_tmp_387 , (~ mux_394_itm) , (~ mux_401_itm) , and_dcpl_642});
  assign weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_2_operator_4_false_2_or_nl
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_4_operator_3_false_1_operator_3_false_1_or_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_14_4_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_13_4_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_12_4_sva_1;
  assign mux_409_nl = MUX_s_1_2_2(mux_tmp_392, mux_tmp_391, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3]);
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_2_operator_4_false_2_or_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_4_operator_3_false_1_operator_3_false_1_or_nl,
      mux_409_nl);
  assign Arbiter_8U_Roundrobin_pick_1_priority_9_4_sva_1 = weight_mem_read_arbxbar_arbiters_next_3_2_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[3]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_11_4_sva_1 = weight_mem_read_arbxbar_arbiters_next_3_4_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[3]);
  assign operator_2_false_3_operator_2_false_3_or_mdf_4_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_11_4_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_10_4_sva_1;
  assign Arbiter_8U_Roundrobin_pick_1_priority_10_4_sva_1 = weight_mem_read_arbxbar_arbiters_next_3_3_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_13_4_sva_1 = weight_mem_read_arbxbar_arbiters_next_3_6_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_14_4_sva_1 = weight_mem_read_arbxbar_arbiters_next_3_7_sva_mx0
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_12_4_sva_1 = weight_mem_read_arbxbar_arbiters_next_3_5_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_4_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_4_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[3])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3]);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_13_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_13_3_sva_1 & (~ Arbiter_8U_Roundrobin_pick_1_priority_14_3_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_7_nl
      = ~(operator_2_false_3_operator_2_false_3_or_mdf_3_sva_1 | mux_415_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_31_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_3_sva_1 & (~ mux_415_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_8_nl
      = ~(operator_2_false_4_operator_2_false_4_or_mdf_3_sva_1 | mux_422_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_33_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_3_sva_1 & (~ mux_422_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_34_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_3_sva_1) & and_dcpl_643;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_35_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_3_sva_1 & and_dcpl_643;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_3_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_13_nl,
      Arbiter_8U_Roundrobin_pick_1_priority_9_3_sva_1, Arbiter_8U_Roundrobin_pick_1_priority_11_3_sva_1,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[2]),
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2]),
      {mux_tmp_408 , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_7_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_31_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_8_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_33_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_34_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_35_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_3_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_1_priority_14_3_sva_1, operator_2_false_3_operator_2_false_3_or_mdf_3_sva_1,
      operator_2_false_4_operator_2_false_4_or_mdf_3_sva_1, operator_2_false_5_operator_2_false_5_or_mdf_3_sva_1,
      {mux_tmp_408 , (~ mux_415_itm) , (~ mux_422_itm) , and_dcpl_643});
  assign weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_2_operator_4_false_2_or_nl
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_3_operator_3_false_1_operator_3_false_1_or_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_14_3_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_13_3_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_12_3_sva_1;
  assign mux_430_nl = MUX_s_1_2_2(mux_tmp_413, mux_tmp_412, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2]);
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_2_operator_4_false_2_or_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_3_operator_3_false_1_operator_3_false_1_or_nl,
      mux_430_nl);
  assign Arbiter_8U_Roundrobin_pick_1_priority_9_3_sva_1 = weight_mem_read_arbxbar_arbiters_next_2_2_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_11_3_sva_1 = weight_mem_read_arbxbar_arbiters_next_2_4_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2]);
  assign operator_2_false_3_operator_2_false_3_or_mdf_3_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_11_3_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_10_3_sva_1;
  assign Arbiter_8U_Roundrobin_pick_1_priority_10_3_sva_1 = weight_mem_read_arbxbar_arbiters_next_2_3_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_13_3_sva_1 = weight_mem_read_arbxbar_arbiters_next_2_6_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_14_3_sva_1 = weight_mem_read_arbxbar_arbiters_next_2_7_sva_mx0
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_12_3_sva_1 = weight_mem_read_arbxbar_arbiters_next_2_5_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_3_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_3_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2]);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_14_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_13_2_sva_1 & (~ Arbiter_8U_Roundrobin_pick_1_priority_14_2_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_9_nl
      = ~(operator_2_false_3_operator_2_false_3_or_mdf_2_sva_1 | mux_438_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_37_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_2_sva_1 & (~ mux_438_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_10_nl
      = ~(operator_2_false_4_operator_2_false_4_or_mdf_2_sva_1 | mux_445_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_39_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_2_sva_1 & (~ mux_445_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_40_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_2_sva_1) & and_dcpl_644;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_41_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_2_sva_1 & and_dcpl_644;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_2_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_14_nl,
      Arbiter_8U_Roundrobin_pick_1_priority_9_2_sva_1, Arbiter_8U_Roundrobin_pick_1_priority_11_2_sva_1,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[1]),
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]),
      {mux_tmp_429 , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_9_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_37_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_10_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_39_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_40_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_41_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_2_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_1_priority_14_2_sva_1, operator_2_false_3_operator_2_false_3_or_mdf_2_sva_1,
      operator_2_false_4_operator_2_false_4_or_mdf_2_sva_1, operator_2_false_5_operator_2_false_5_or_mdf_2_sva_1,
      {mux_tmp_429 , (~ mux_438_itm) , (~ mux_445_itm) , and_dcpl_644});
  assign weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_2_operator_4_false_2_or_nl
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1]);
  assign weight_mem_read_arbxbar_xbar_1_for_3_2_operator_3_false_1_operator_3_false_1_or_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_14_2_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_13_2_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_12_2_sva_1;
  assign mux_455_nl = MUX_s_1_2_2(mux_tmp_436, mux_tmp_435, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1]);
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_2_operator_4_false_2_or_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_2_operator_3_false_1_operator_3_false_1_or_nl,
      mux_455_nl);
  assign Arbiter_8U_Roundrobin_pick_1_priority_9_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_2_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_11_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_4_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]);
  assign operator_2_false_3_operator_2_false_3_or_mdf_2_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_11_2_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_10_2_sva_1;
  assign Arbiter_8U_Roundrobin_pick_1_priority_10_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_3_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_13_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_6_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_14_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_7_sva_mx0
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_12_2_sva_1 = weight_mem_read_arbxbar_arbiters_next_1_5_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_2_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_2_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1]);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_15_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_13_1_sva_1 & (~ Arbiter_8U_Roundrobin_pick_1_priority_14_1_sva_1);
  assign weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_3_nl
      = weight_mem_read_arbxbar_arbiters_next_0_2_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0]);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_11_nl
      = ~(operator_2_false_3_operator_2_false_3_or_mdf_1_sva_1 | mux_461_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_43_nl
      = operator_2_false_3_operator_2_false_3_or_mdf_1_sva_1 & (~ mux_461_itm);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_44_nl
      = (~ operator_2_false_4_operator_2_false_4_or_mdf_1_sva_1) & and_dcpl_646;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_45_nl
      = operator_2_false_4_operator_2_false_4_or_mdf_1_sva_1 & and_dcpl_646;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_46_nl
      = (~ operator_2_false_5_operator_2_false_5_or_mdf_1_sva_1) & and_dcpl_651;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_47_nl
      = operator_2_false_5_operator_2_false_5_or_mdf_1_sva_1 & and_dcpl_651;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_1_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2(nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_15_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_3_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp,
      (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]), (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0]),
      (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0]), (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0]),
      {mux_tmp_454 , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_nor_11_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_43_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_44_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_45_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_46_nl
      , nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_1_and_47_nl});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_1_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_1_priority_14_1_sva_1, operator_2_false_3_operator_2_false_3_or_mdf_1_sva_1,
      operator_2_false_4_operator_2_false_4_or_mdf_1_sva_1, operator_2_false_5_operator_2_false_5_or_mdf_1_sva_1,
      {mux_tmp_454 , (~ mux_461_itm) , and_dcpl_646 , and_dcpl_651});
  assign weight_mem_read_arbxbar_xbar_1_for_3_1_operator_3_false_1_operator_3_false_1_or_nl
      = Arbiter_8U_Roundrobin_pick_1_priority_14_1_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_13_1_sva_1
      | (weight_mem_read_arbxbar_arbiters_next_0_5_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0]));
  assign weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_2_operator_4_false_2_or_nl
      = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0]);
  assign mux_470_nl = MUX_s_1_2_2(mux_tmp_459, mux_tmp_458, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]);
  assign and_679_nl = (~ mux_470_nl) & and_dcpl_645;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0
      = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_1_operator_3_false_1_operator_3_false_1_or_nl,
      weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_2_operator_4_false_2_or_nl,
      and_679_nl);
  assign weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp
      = weight_mem_read_arbxbar_arbiters_next_0_4_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0]);
  assign operator_2_false_3_operator_2_false_3_or_mdf_1_sva_1 = weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_1_tmp;
  assign weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_1_tmp
      = weight_mem_read_arbxbar_arbiters_next_0_3_sva_mx1 & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[0]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_13_1_sva_1 = weight_mem_read_arbxbar_arbiters_next_0_6_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]);
  assign Arbiter_8U_Roundrobin_pick_1_priority_14_1_sva_1 = weight_mem_read_arbxbar_arbiters_next_0_7_sva_mx0
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0]);
  assign operator_2_false_4_operator_2_false_4_or_mdf_1_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0]);
  assign operator_2_false_5_operator_2_false_5_or_mdf_1_sva_1 = (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[0]);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_3_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_3,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_3,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_4_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_4,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_5_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_5,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_5_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_6_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_6,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_0_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_0,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_2_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_2,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_2,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_1_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_1,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_3_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_3_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_3,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_4_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_4_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_4_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_5_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_5_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_5_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_6_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_6_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_6_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_0_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_0_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_2_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_2_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_2,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_1_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_1_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_3_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_3_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_3,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_4_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_4_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_5_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_5_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_5_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_6_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_6_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_0_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_0_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_2_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_2_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_2,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_1_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_1_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_1,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_3_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_3_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_3,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_4_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_4_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_5_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_5_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_5_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_6_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_6_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_0_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_0_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_2_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_2_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_2,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_1_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_1_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_3_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_3_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_3_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_4_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_4_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_5_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_5_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_5_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_6_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_6_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_0_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_0_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_2_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_2_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_2_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_1_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_1_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_1_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_53_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_5_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_65_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_5_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_77_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_5_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_89_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_5_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_101_tmp =
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_5_cse & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_113_tmp =
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_5_cse & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_2_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_3
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_6_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_3
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_10_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_3
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_14_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_3
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_18_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_3
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_22_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_3_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_26_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_3
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_30_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_3
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_52_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_1
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_64_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_1
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_76_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_1
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_88_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_1
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_100_tmp =
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_1_cse & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_112_tmp =
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_1 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_124_tmp =
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_1 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_122_tmp =
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_2 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_126_tmp =
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_0 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_110_tmp =
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_2 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_114_tmp =
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_0 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_98_tmp = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_2_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_102_tmp =
      Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_0 & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_86_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_2
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_90_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_0
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_74_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_2
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_78_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_0
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_6_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_6_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_4_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_4_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_62_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_2
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_66_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_0
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_1 = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_cse
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_50_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_2
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_54_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_0
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_6_1 = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_6
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  assign Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_4_1 = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_4
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_38_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_2
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  assign Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_42_tmp = Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_0
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1;
  assign nl_PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1 = (pe_manager_base_weight_sva_mx2[14:4])
      + PEManager_15U_GetWeightAddr_else_acc_3_1;
  assign PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1 = nl_PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1[10:0];
  assign weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_1_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_1_lpi_1_dfm_mx0);
  assign weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_2_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_2_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_2_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_2_sva_1));
  assign operator_7_false_1_operator_7_false_1_or_mdf_2_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_14_2_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_13_2_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_12_2_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_11_2_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_10_2_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_9_2_sva_1 | (weight_mem_read_arbxbar_arbiters_next_1_1_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1]));
  assign weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_3_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_3_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_3_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_3_sva_1));
  assign operator_7_false_1_operator_7_false_1_or_mdf_3_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_14_3_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_13_3_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_12_3_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_11_3_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_10_3_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_9_3_sva_1 | (weight_mem_read_arbxbar_arbiters_next_2_1_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[2]));
  assign weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_4_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_4_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_4_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_4_sva_1));
  assign operator_7_false_1_operator_7_false_1_or_mdf_4_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_14_4_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_13_4_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_12_4_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_11_4_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_10_4_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_9_4_sva_1 | (weight_mem_read_arbxbar_arbiters_next_3_1_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[3]));
  assign weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_5_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_5_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_5_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_5_sva_1));
  assign operator_7_false_1_operator_7_false_1_or_mdf_5_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_14_5_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_13_5_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_12_5_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_11_5_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_10_5_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_9_5_sva_1 | (weight_mem_read_arbxbar_arbiters_next_4_1_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[4]));
  assign weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_6_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_6_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_6_lpi_1_dfm_mx0);
  assign weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_7_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_7_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_7_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_7_sva_1));
  assign operator_7_false_1_operator_7_false_1_or_mdf_7_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_14_7_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_13_7_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_12_7_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_11_7_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_10_7_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_9_7_sva_1 | (weight_mem_read_arbxbar_arbiters_next_6_1_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6]));
  assign operator_7_false_1_operator_7_false_1_or_mdf_sva_1 = Arbiter_8U_Roundrobin_pick_1_priority_14_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_13_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_12_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_11_sva_1 | Arbiter_8U_Roundrobin_pick_1_priority_10_sva_1
      | Arbiter_8U_Roundrobin_pick_1_priority_9_sva_1 | (weight_mem_read_arbxbar_arbiters_next_7_1_sva_mx1
      & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7]));
  assign weight_read_addrs_0_3_0_lpi_1_dfm_4 = MUX_v_4_2_2(4'b0000, pe_manager_base_weight_sva_mx1_3_0,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign nl_operator_4_false_acc_sdt_sva_1 = conv_u2s_4_5(pe_config_num_manager_sva)
      + 5'b11111;
  assign operator_4_false_acc_sdt_sva_1 = nl_operator_4_false_acc_sdt_sva_1[4:0];
  assign while_and_1129_cse_1 = (~ while_if_and_tmp_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign while_if_and_tmp_1 = PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_nor_1_cse_1
      & reg_rva_in_reg_rw_sva_st_1_1_cse;
  assign PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_nor_1_cse_1
      = ~(PECore_DecodeAxiWrite_switch_lp_equal_tmp_1 | PECore_DecodeAxiWrite_switch_lp_equal_tmp_2
      | PECore_DecodeAxiWrite_switch_lp_nor_tmp_1);
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_8_nl = start_PopNB_mioi_data_rsc_z_mxwt
      & pe_config_is_valid_sva & start_PopNB_mioi_return_rsc_z_mxwt;
  assign PECore_UpdateFSM_case_1_if_PECore_UpdateFSM_case_1_if_and_nl = pe_config_is_zero_first_sva
      & pe_manager_zero_active_sva;
  assign PECore_UpdateFSM_switch_lp_pe_config_UpdateManagerCounter_nand_nl = ~(pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_if_nor_mdf_sva_1
      & pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1);
  assign PECore_UpdateFSM_switch_lp_mux1h_14_nl = MUX1HOT_s_1_4_2(PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_and_8_nl,
      PECore_UpdateFSM_case_1_if_PECore_UpdateFSM_case_1_if_and_nl, pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_nor_mdf_sva_st_1,
      PECore_UpdateFSM_switch_lp_pe_config_UpdateManagerCounter_nand_nl, {PECore_UpdateFSM_switch_lp_and_7_itm_1
      , PECore_UpdateFSM_switch_lp_equal_tmp_2_1 , PECore_UpdateFSM_switch_lp_equal_tmp_3_1
      , PECore_UpdateFSM_switch_lp_equal_tmp_5_1});
  assign PECore_UpdateFSM_next_state_0_lpi_1_dfm_4 = PECore_UpdateFSM_switch_lp_mux1h_14_nl
      & PECore_UpdateFSM_switch_lp_nor_7_itm_1;
  assign pe_config_UpdateManagerCounter_if_if_unequal_tmp = pe_config_output_counter_sva
      != (operator_8_false_acc_sdt_sva_1[7:0]);
  assign pe_config_UpdateManagerCounter_if_pe_config_UpdateManagerCounter_if_if_nor_mdf_sva_1
      = ~(pe_config_UpdateManagerCounter_if_if_unequal_tmp | (operator_8_false_acc_sdt_sva_1[8]));
  assign input_write_req_valid_lpi_1_dfm_5 = PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva_mx1
      & PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_cse_1;
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_cse_1 = ~(PECore_RunFSM_switch_lp_equal_tmp_1_mx0w1
      | PECore_RunFSM_switch_lp_nor_tmp_1);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_pmx_sva_1
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:56]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:56]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[55:48]),
      {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_12_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000002
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[55:48]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[55:48]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[47:40]),
      {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_12_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000003
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:40]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:40]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[39:32]),
      {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_12_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000004
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[39:32]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[39:32]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[31:24]),
      {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_12_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000005
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[23:16]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[23:16]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[15:8]),
      {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_12_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000006
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:24]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31:24]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[23:16]),
      {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_12_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:56]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:56]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[55:48]),
      {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_1_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[55:48]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[55:48]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[47:40]),
      {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_1_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_6_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:40]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:40]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[39:32]),
      {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_1_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_5_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[39:32]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[39:32]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[31:24]),
      {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_1_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:24]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31:24]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[23:16]),
      {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_1_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_3_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[23:16]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[23:16]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[15:8]),
      {weight_read_addrs_4_14_2_lpi_1_dfm_3_0 , pe_manager_base_weight_slc_pe_manager_base_weight_1_0_1_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:56]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:56]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[55:48]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_2_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[55:48]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[55:48]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[47:40]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_2_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_6_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:40]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:40]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[39:32]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_2_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_5_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[39:32]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[39:32]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[31:24]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_2_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:24]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31:24]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[23:16]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_2_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_3_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2
      = MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[23:16]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[23:16]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[15:8]),
      {weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 , reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_2_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_65_cse = reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_2_cse
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000002
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:24]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31:24]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[23:16]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_65_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_118
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_120 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_122 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_71_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_72_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000003
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[23:16]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[23:16]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[15:8]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_65_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_118
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_120 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_76_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_122 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_78_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_79_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_80_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000002
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:24]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31:24]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[23:16]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_100 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_44_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_62_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_48_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000003
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[23:16]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[23:16]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[15:8]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_100 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_44_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_46_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_47_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_48_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000004
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:40]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:40]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[39:32]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_100 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_60_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_62_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_48_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000005
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[39:32]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[39:32]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[31:24]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_98 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_60_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_62_itm_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_48_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_mux1h_34_nl = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[63:56]),
      (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63:56]),
      (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63:56]), (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63:56]),
      (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[55:48]), {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_100
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_44_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_62_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_8_cse_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_pmx_000000
      = MUX_v_8_2_2(8'b00000000, crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_mux1h_34_nl,
      weight_mem_run_3_for_land_2_lpi_1_dfm_2);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000006
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[55:48]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[55:48]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[47:40]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_100 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_2_cse_1
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_3_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_44_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_5_cse_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_46_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_47_itm_1 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_48_itm_1});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000000
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[55:48]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[55:48]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[55:48]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[55:48]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[47:40]),
      {weight_mem_run_3_for_5_and_161_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_14_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_15_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_17_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_3
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_19_itm_2 , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_20_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_21_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_2_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000001
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[47:40]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[47:40]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[47:40]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[47:40]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[39:32]),
      {crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_21_nl , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_54_itm_2
      , reg_weight_mem_run_3_for_5_and_163_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_itm_2
      , reg_weight_mem_run_3_for_5_and_165_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_2
      , reg_weight_mem_run_3_for_5_and_167_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_44_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000002
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[39:32]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[39:32]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[39:32]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[39:32]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[31:24]),
      {weight_mem_run_3_for_5_and_161_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_54_itm_2
      , reg_weight_mem_run_3_for_5_and_163_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_56_itm_2
      , reg_weight_mem_run_3_for_5_and_165_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_34_itm_2
      , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_35_itm_2 , reg_weight_mem_run_3_for_5_and_168_itm_2_cse});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000003
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:24]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[31:24]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[31:24]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[31:24]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[23:16]),
      {weight_mem_run_3_for_5_and_161_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_54_itm_2
      , reg_weight_mem_run_3_for_5_and_163_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_56_itm_2
      , reg_weight_mem_run_3_for_5_and_165_itm_2_cse , reg_weight_mem_run_3_for_5_and_166_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_167_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_44_itm_2});
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000004
      = MUX1HOT_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[23:16]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[23:16]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[23:16]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[23:16]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[15:8]),
      {weight_mem_run_3_for_5_and_161_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_54_itm_2
      , reg_weight_mem_run_3_for_5_and_163_itm_2_cse , crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_56_itm_2
      , reg_weight_mem_run_3_for_5_and_165_itm_2_cse , reg_weight_mem_run_3_for_5_and_166_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_167_itm_2_cse , reg_weight_mem_run_3_for_5_and_168_itm_2_cse});
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_5_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
      = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_8 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_8 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_8 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_8 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_8 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0;
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_3_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_3,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_3_mx0,
      or_dcpl_678);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_4_mx0
      = MUX_s_1_2_2(reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4_cse,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_4_mx0,
      or_dcpl_678);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_5_mx0
      = MUX_s_1_2_2(reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_5_cse,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_5_mx0,
      or_dcpl_678);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_6_mx0
      = MUX_s_1_2_2(reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6_cse,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_6_mx0,
      or_dcpl_678);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_0_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_0_mx0,
      or_dcpl_678);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_2_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_2,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_2_mx0,
      or_dcpl_678);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_1_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1_1,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_1_mx0,
      or_dcpl_678);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_3_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_3_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_4_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_4_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_5_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_5_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_5_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_6_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_6_mx0,
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_0_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_0_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_0,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_2_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_2_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_2,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_1_mx0
      = MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_1_mx0,
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1,
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_8 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0);
  assign nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_0_1
      = Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_8 & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_1_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_8 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_1_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_1_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_8 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_1_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_1_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_8 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_1_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_1_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_8 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_1_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_1_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_9 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_2_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_2_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_9 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_2_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_2_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_9 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_2_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_2_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_9 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_2_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_2_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_10 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_3_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_3_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_10 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_3_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_3_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_10 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_3_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_3_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_10 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_3_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_3_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_11 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_4_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_4_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_11 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_4_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_4_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_11 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_4_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_4_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_11 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_4_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_4_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_12 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_5_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_5_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_12 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_5_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_5_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_12 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_5_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_5_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_12 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_5_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_5_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_13 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_6_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_6_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_13 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_6_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_6_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_13 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_6_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_6_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_13 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_6_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_6_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_14 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_7_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_7_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_14 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_7_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_7_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_14 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_7_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_7_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_14 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_7_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_7_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_2_15 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_0_15 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_1_15 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_and_stg_1_3_15 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_lpi_1_dfm_mx0;
  assign PECore_DecodeAxiWrite_case_4_switch_lp_or_cse_1 = and_321_cse | PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_mx0w0;
  assign nl_operator_16_false_acc_sdt_sva_1 = conv_u2s_8_9(pe_manager_num_input_sva)
      + 9'b111111111;
  assign operator_16_false_acc_sdt_sva_1 = nl_operator_16_false_acc_sdt_sva_1[8:0];
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_1_cse_1 = ~((state_mux_1_cse!=2'b00)
      | state_0_sva_mx1);
  assign PECore_UpdateFSM_switch_lp_nor_tmp_1 = ~(PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_1_cse_1
      | PECore_UpdateFSM_switch_lp_equal_tmp_6 | PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_1_cse_1
      | PECore_RunScale_PECore_RunScale_if_and_1_svs_1 | PECore_PushOutput_PECore_PushOutput_if_and_svs_1);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_136_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_1_itm_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_54_nl
      = MUX_v_4_2_2(4'b0000, (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[55:52]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_136_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_137_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_1_itm_2[1]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_62_nl
      = MUX_v_4_2_2(4'b0000, (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[55:52]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_137_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_8_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_64_63_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_2_0_8_7_0_sdt_47_40_sva_1_7_4
      = MUX_v_4_8_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_6_itm_1[7:4]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1_7_4,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_22_itm_1[7:4]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_30_itm_1[7:4]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_38_itm_1[7:4]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_46_itm_1[7:4]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_54_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_62_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_89_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_1_itm_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_64_nl
      = MUX_v_4_2_2(4'b0000, (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[51:48]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_89_nl);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_82_nl = ~ (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_1_itm_2[1]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_65_nl
      = MUX_v_4_2_2(4'b0000, (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[51:48]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_82_nl);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_8_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_64_63_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_2_0_8_7_0_sdt_47_40_sva_1_3_0
      = MUX_v_4_8_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_6_itm_1[3:0]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1_3_0,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_22_itm_1[3:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_30_itm_1[3:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_38_itm_1[3:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_46_itm_1[3:0]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_64_nl,
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_65_nl,
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse);
  assign mux1h_7_nl = MUX1HOT_s_1_8_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_7_itm_1[7]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1_7,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_23_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_31_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_47_itm_1[7]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[63]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[63]),
      weight_port_read_out_data_0_7_sva_dfm_2_7, {and_931_cse , and_932_cse , and_933_cse
      , and_934_cse , and_935_cse , and_936_cse , and_937_cse , nor_524_cse});
  assign weight_port_read_out_data_0_7_sva_dfm_3_7 = mux1h_7_nl & (~ or_dcpl_684);
  assign mux1h_16_nl = MUX1HOT_v_7_8_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_7_itm_1[6:0]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1_6_0,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_23_itm_1[6:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_31_itm_1[6:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_47_itm_1[6:0]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[62:56]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[62:56]),
      weight_port_read_out_data_0_7_sva_dfm_2_6_0, {and_931_cse , and_932_cse , and_933_cse
      , and_934_cse , and_935_cse , and_936_cse , and_937_cse , nor_524_cse});
  assign not_2551_nl = ~ or_dcpl_684;
  assign weight_port_read_out_data_0_7_sva_dfm_3_6_0 = MUX_v_7_2_2(7'b0000000, mux1h_16_nl,
      not_2551_nl);
  assign or_1407_tmp = ((pe_manager_base_weight_slc_pe_manager_base_weight_1_0_1_itm_2[1])
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_44_itm_2) | and_dcpl_665;
  assign and_967_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_for_and_52 & (~ or_1407_tmp);
  assign and_968_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_for_asn_56 & (~ or_1407_tmp);
  assign and_969_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_for_or_cse & (~ or_1407_tmp);
  assign and_970_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_71_itm_1
      & (~ or_1407_tmp);
  assign and_971_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_60_itm_1
      & (~ or_1407_tmp);
  assign and_972_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_47_itm_1
      & (~ or_1407_tmp);
  assign and_973_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_44_itm_2
      & (~ or_1407_tmp);
  assign nor_528_ssc = ~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3
      | or_1407_tmp);
  assign mux1h_8_nl = MUX1HOT_v_4_8_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_5_itm_1[7:4]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1_7_4,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_21_itm_1[7:4]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_29_itm_1[7:4]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_45_itm_1[7:4]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[47:44]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[47:44]),
      weight_port_read_out_data_0_5_sva_dfm_2_7_4, {and_967_ssc , and_968_ssc , and_969_ssc
      , and_970_ssc , and_971_ssc , and_972_ssc , and_973_ssc , nor_528_ssc});
  assign not_2552_nl = ~ or_1407_tmp;
  assign weight_port_read_out_data_0_5_sva_dfm_3_7_4 = MUX_v_4_2_2(4'b0000, mux1h_8_nl,
      not_2552_nl);
  assign mux1h_17_nl = MUX1HOT_v_4_8_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_5_itm_1[3:0]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1_3_0,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_21_itm_1[3:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_29_itm_1[3:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_45_itm_1[3:0]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[43:40]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[43:40]),
      weight_port_read_out_data_0_5_sva_dfm_2_3_0, {and_967_ssc , and_968_ssc , and_969_ssc
      , and_970_ssc , and_971_ssc , and_972_ssc , and_973_ssc , nor_528_ssc});
  assign not_2463_nl = ~ or_1407_tmp;
  assign weight_port_read_out_data_0_5_sva_dfm_3_3_0 = MUX_v_4_2_2(4'b0000, mux1h_17_nl,
      not_2463_nl);
  assign and_976_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_for_and_54 & (~ or_dcpl_684);
  assign and_979_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_71_itm_1
      & (~ or_dcpl_684);
  assign and_980_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_72_itm_1
      & (~ or_dcpl_684);
  assign mux1h_9_nl = MUX1HOT_s_1_8_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_4_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_itm_1_7_6[1]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1_7,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_28_itm_1[7]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_44_itm_1[7]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[39]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[39]),
      weight_port_read_out_data_0_4_sva_dfm_2_7, {and_976_ssc , and_932_cse , and_933_cse
      , and_979_ssc , and_980_ssc , and_936_cse , and_937_cse , nor_524_cse});
  assign weight_port_read_out_data_0_4_sva_dfm_3_7 = mux1h_9_nl & (~ or_dcpl_684);
  assign mux1h_18_nl = MUX1HOT_s_1_8_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_4_itm_1[6]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_itm_1_7_6[0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1_6_0[6]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_28_itm_1[6]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_44_itm_1[6]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[38]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[38]),
      weight_port_read_out_data_0_4_sva_dfm_2_6, {and_976_ssc , and_932_cse , and_933_cse
      , and_979_ssc , and_980_ssc , and_936_cse , and_937_cse , nor_524_cse});
  assign weight_port_read_out_data_0_4_sva_dfm_3_6 = mux1h_18_nl & (~ or_dcpl_684);
  assign mux1h_19_nl = MUX1HOT_v_6_8_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_4_itm_1[5:0]),
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_itm_1_5_0,
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1_6_0[5:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_28_itm_1[5:0]),
      (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_44_itm_1[5:0]),
      (weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d[37:32]), (weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[37:32]),
      weight_port_read_out_data_0_4_sva_dfm_2_5_0, {and_976_ssc , and_932_cse , and_933_cse
      , and_979_ssc , and_980_ssc , and_936_cse , and_937_cse , nor_524_cse});
  assign not_2553_nl = ~ or_dcpl_684;
  assign weight_port_read_out_data_0_4_sva_dfm_3_5_0 = MUX_v_6_2_2(6'b000000, mux1h_19_nl,
      not_2553_nl);
  assign weight_mem_run_1_if_for_weight_mem_run_1_if_for_weight_mem_run_1_if_for_nor_tmp
      = ~((~ PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2) | reg_rva_in_reg_rw_sva_2_cse
      | (~((weight_mem_read_arbxbar_xbar_for_1_lshift_tmp!=8'b00000000))) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[0])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[0])) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[1])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[1])) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[2])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[2])) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[3])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[3])) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[4])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[4])) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[5])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[5])) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[6])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[6])) | ((weight_mem_write_arbxbar_xbar_for_lshift_tmp[7])
      & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[7])));
  assign PECore_DecodeAxiWrite_switch_lp_or_5_cse_1 = PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0 | PECore_DecodeAxiWrite_switch_lp_nor_tmp_1_1;
  assign rva_out_reg_data_63_sva_dfm_7 = PECore_PushAxiRsp_mux_13_itm_1 & rva_in_reg_rw_sva_5;
  assign PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1 = ~(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_11_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign input_mem_banks_write_if_for_if_and_stg_6_0_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_0_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_1_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_1_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_2_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_2_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_3_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_3_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_4_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_4_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_5_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_5_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_6_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_6_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_7_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_7_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_8_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_8_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_9_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_9_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_10_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_10_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_11_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_11_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_12_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_12_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_13_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_13_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_14_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_14_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_15_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_15_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_16_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_16_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_17_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_17_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_18_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_18_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_19_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_19_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_20_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_20_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_21_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_21_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_22_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_22_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_23_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_23_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_24_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_24_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_25_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_25_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_26_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_26_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_27_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_27_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_28_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_28_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_29_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_29_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_30_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_30_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_31_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_31_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_32_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_32_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_33_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_33_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_34_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_34_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_35_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_35_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_36_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_36_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_37_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_37_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_38_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_38_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_39_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_39_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_40_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_40_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_41_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_41_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_42_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_42_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_43_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_43_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_44_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_44_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_45_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_45_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_46_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_46_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_47_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_47_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_48_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_48_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_49_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_49_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_50_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_50_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_51_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_51_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_52_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_52_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_53_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_53_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_54_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_54_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_55_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_55_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_56_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_56_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_57_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_57_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_58_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_58_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_59_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_59_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_60_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_60_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_61_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_61_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_62_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_62_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_63_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_63_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]));
  assign input_mem_banks_write_if_for_if_and_stg_6_64_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_0_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_65_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_1_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_66_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_2_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_67_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_3_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_68_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_4_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_69_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_5_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_70_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_6_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_71_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_7_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_72_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_8_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_73_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_9_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_74_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_10_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_75_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_11_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_76_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_12_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_77_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_13_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_78_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_14_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_79_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_15_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_80_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_16_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_81_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_17_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_82_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_18_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_83_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_19_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_84_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_20_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_85_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_21_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_86_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_22_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_87_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_23_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_88_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_24_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_89_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_25_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_90_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_26_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_91_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_27_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_92_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_28_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_93_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_29_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_94_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_30_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_95_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_31_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_96_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_32_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_97_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_33_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_98_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_34_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_99_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_35_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_100_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_36_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_101_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_37_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_102_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_38_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_103_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_39_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_104_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_40_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_105_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_41_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_106_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_42_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_107_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_43_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_108_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_44_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_109_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_45_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_110_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_46_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_111_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_47_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_112_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_48_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_113_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_49_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_114_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_50_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_115_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_51_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_116_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_52_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_117_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_53_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_118_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_54_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_119_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_55_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_120_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_56_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_121_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_57_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_122_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_58_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_123_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_59_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_124_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_60_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_125_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_61_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_126_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_62_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_6_127_sva_1 = input_mem_banks_write_if_for_if_and_stg_5_63_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[6]);
  assign input_mem_banks_write_if_for_if_and_stg_5_0_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_0_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_1_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_1_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_2_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_2_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_3_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_3_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_4_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_4_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_5_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_5_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_6_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_6_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_7_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_7_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_8_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_8_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_9_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_9_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_10_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_10_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_11_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_11_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_12_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_12_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_13_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_13_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_14_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_14_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_15_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_15_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_16_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_16_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_17_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_17_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_18_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_18_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_19_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_19_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_20_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_20_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_21_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_21_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_22_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_22_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_23_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_23_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_24_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_24_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_25_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_25_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_26_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_26_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_27_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_27_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_28_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_28_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_29_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_29_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_30_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_30_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_31_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_31_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]));
  assign input_mem_banks_write_if_for_if_and_stg_5_32_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_0_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_33_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_1_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_34_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_2_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_35_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_3_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_36_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_4_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_37_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_5_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_38_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_6_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_39_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_7_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_40_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_8_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_41_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_9_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_42_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_10_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_43_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_11_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_44_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_12_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_45_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_13_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_46_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_14_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_47_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_15_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_48_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_16_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_49_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_17_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_50_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_18_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_51_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_19_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_52_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_20_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_53_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_21_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_54_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_22_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_55_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_23_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_56_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_24_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_57_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_25_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_58_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_26_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_59_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_27_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_60_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_28_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_61_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_29_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_62_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_30_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_5_63_sva_1 = input_mem_banks_write_if_for_if_and_stg_4_31_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[5]);
  assign input_mem_banks_write_if_for_if_and_stg_4_0_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_0_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_1_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_1_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_2_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_2_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_3_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_3_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_4_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_4_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_5_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_5_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_6_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_6_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_7_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_7_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_8_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_8_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_9_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_9_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_10_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_10_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_11_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_11_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_12_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_12_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_13_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_13_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_14_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_14_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_15_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_15_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]));
  assign input_mem_banks_write_if_for_if_and_stg_4_16_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_0_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_17_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_1_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_18_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_2_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_19_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_3_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_20_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_4_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_21_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_5_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_22_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_6_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_23_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_7_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_24_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_8_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_25_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_9_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_26_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_10_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_27_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_11_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_28_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_12_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_29_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_13_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_30_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_14_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_4_31_sva_1 = input_mem_banks_write_if_for_if_and_stg_3_15_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[4]);
  assign input_mem_banks_write_if_for_if_and_stg_3_0_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_0_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_1_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_1_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_2_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_2_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_3_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_3_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_4_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_4_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_5_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_5_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_6_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_6_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_7_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_7_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]));
  assign input_mem_banks_write_if_for_if_and_stg_3_8_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_0_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_3_9_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_1_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_3_10_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_2_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_3_11_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_3_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_3_12_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_4_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_3_13_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_5_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_3_14_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_6_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_3_15_sva_1 = input_mem_banks_write_if_for_if_and_stg_2_7_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[3]);
  assign input_mem_banks_write_if_for_if_and_stg_2_0_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_0_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]));
  assign input_mem_banks_write_if_for_if_and_stg_2_1_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_1_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]));
  assign input_mem_banks_write_if_for_if_and_stg_2_2_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_2_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]));
  assign input_mem_banks_write_if_for_if_and_stg_2_3_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_3_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]));
  assign input_mem_banks_write_if_for_if_and_stg_2_4_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_0_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]);
  assign input_mem_banks_write_if_for_if_and_stg_2_5_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_1_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]);
  assign input_mem_banks_write_if_for_if_and_stg_2_6_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_2_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]);
  assign input_mem_banks_write_if_for_if_and_stg_2_7_sva_1 = input_mem_banks_write_if_for_if_and_stg_1_3_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[2]);
  assign input_mem_banks_write_if_for_if_and_stg_1_0_sva_1 = ~((while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[1:0]!=2'b00));
  assign input_mem_banks_write_if_for_if_and_stg_1_1_sva_1 = (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[1:0]==2'b01);
  assign input_mem_banks_write_if_for_if_and_stg_1_2_sva_1 = (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[1:0]==2'b10);
  assign input_mem_banks_write_if_for_if_and_stg_1_3_sva_1 = (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[1:0]==2'b11);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_0_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_0_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_1_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_1_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_2_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_2_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_3_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_3_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_4_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_4_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_5_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_5_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_6_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_6_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_7_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_7_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_8_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_8_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_9_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_9_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_10_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_10_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_11_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_11_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_12_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_12_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_13_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_13_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_14_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_14_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_15_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_15_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_16_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_16_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_17_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_17_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_18_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_18_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_19_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_19_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_20_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_20_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_21_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_21_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_22_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_22_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_23_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_23_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_24_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_24_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_25_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_25_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_26_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_26_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_27_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_27_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_28_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_28_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_29_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_29_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_30_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_30_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_31_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_31_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_32_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_32_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_33_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_33_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_34_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_34_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_35_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_35_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_36_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_36_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_37_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_37_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_38_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_38_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_39_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_39_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_40_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_40_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_41_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_41_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_42_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_42_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_43_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_43_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_44_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_44_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_45_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_45_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_46_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_46_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_47_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_47_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_48_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_48_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_49_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_49_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_50_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_50_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_51_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_51_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_52_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_52_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_53_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_53_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_54_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_54_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_55_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_55_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_56_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_56_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_57_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_57_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_58_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_58_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_59_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_59_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_60_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_60_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_61_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_61_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_62_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_62_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_63_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_63_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[6]));
  assign input_mem_banks_write_1_if_for_if_and_stg_6_64_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_0_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_65_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_1_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_66_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_2_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_67_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_3_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_68_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_4_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_69_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_5_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_70_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_6_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_71_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_7_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_72_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_8_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_73_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_9_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_74_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_10_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_75_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_11_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_76_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_12_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_77_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_13_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_78_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_14_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_79_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_15_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_80_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_16_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_81_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_17_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_82_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_18_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_83_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_19_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_84_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_20_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_85_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_21_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_86_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_22_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_87_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_23_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_88_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_24_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_89_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_25_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_90_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_26_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_91_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_27_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_92_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_28_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_93_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_29_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_94_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_30_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_95_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_31_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_96_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_32_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_97_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_33_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_98_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_34_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_99_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_35_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_100_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_36_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_101_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_37_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_102_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_38_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_103_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_39_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_104_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_40_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_105_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_41_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_106_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_42_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_107_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_43_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_108_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_44_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_109_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_45_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_110_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_46_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_111_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_47_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_112_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_48_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_113_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_49_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_114_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_50_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_115_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_51_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_116_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_52_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_117_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_53_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_118_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_54_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_119_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_55_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_120_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_56_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_121_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_57_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_122_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_58_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_123_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_59_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_124_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_60_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_125_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_61_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_126_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_62_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign input_mem_banks_write_1_if_for_if_and_stg_6_127_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_5_63_sva_1
      & (input_write_addrs_lpi_1_dfm_2[6]);
  assign nl_PEManager_15U_GetInputAddr_acc_tmp = input_port_PopNB_mioi_data_logical_addr_rsc_z_mxwt
      + (pe_manager_base_input_sva[7:0]);
  assign PEManager_15U_GetInputAddr_acc_tmp = nl_PEManager_15U_GetInputAddr_acc_tmp[7:0];
  assign input_write_addrs_lpi_1_dfm_2 = PEManager_15U_GetInputAddr_acc_tmp & ({{7{PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva_mx1}},
      PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva_mx1})
      & ({{7{PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_cse_1}}, PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_cse_1});
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_257_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_127_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_255_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_127_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_256_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_126_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_254_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_126_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_255_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_125_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_253_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_125_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_254_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_124_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_252_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_124_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_253_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_123_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_251_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_123_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_252_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_122_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_250_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_122_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_251_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_121_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_249_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_121_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_250_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_120_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_248_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_120_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_249_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_119_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_247_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_119_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_248_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_118_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_246_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_118_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_247_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_117_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_245_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_117_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_246_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_116_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_244_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_116_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_245_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_115_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_243_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_115_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_244_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_114_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_242_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_114_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_243_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_113_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_241_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_113_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_242_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_112_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_240_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_112_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_241_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_111_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_239_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_111_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_240_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_110_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_238_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_110_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_239_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_109_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_237_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_109_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_238_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_108_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_236_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_108_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_237_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_107_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_235_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_107_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_236_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_106_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_234_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_106_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_235_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_105_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_233_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_105_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_234_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_104_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_232_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_104_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_233_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_103_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_231_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_103_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_232_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_102_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_230_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_102_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_231_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_101_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_229_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_101_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_230_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_100_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_228_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_100_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_229_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_99_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_227_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_99_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_228_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_98_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_226_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_98_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_227_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_97_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_225_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_97_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_226_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_96_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_224_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_96_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_225_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_95_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_223_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_95_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_224_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_94_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_222_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_94_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_223_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_93_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_221_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_93_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_222_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_92_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_220_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_92_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_221_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_91_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_219_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_91_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_220_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_90_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_218_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_90_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_219_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_89_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_217_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_89_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_218_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_88_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_216_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_88_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_217_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_87_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_215_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_87_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_216_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_86_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_214_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_86_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_215_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_85_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_213_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_85_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_214_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_84_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_212_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_84_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_213_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_83_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_211_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_83_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_212_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_82_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_210_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_82_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_211_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_81_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_209_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_81_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_210_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_80_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_208_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_80_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_209_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_79_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_207_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_79_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_208_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_78_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_206_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_78_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_207_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_77_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_205_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_77_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_206_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_76_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_204_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_76_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_205_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_75_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_203_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_75_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_204_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_74_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_202_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_74_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_203_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_73_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_201_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_73_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_202_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_72_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_200_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_72_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_201_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_71_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_199_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_71_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_200_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_70_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_198_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_70_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_199_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_69_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_197_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_69_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_198_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_68_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_196_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_68_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_197_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_67_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_195_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_67_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_196_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_66_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_194_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_66_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_195_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_65_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_193_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_65_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_194_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_64_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_192_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_64_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_193_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_63_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_191_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_63_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_192_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_62_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_190_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_62_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_191_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_61_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_189_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_61_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_190_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_60_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_188_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_60_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_189_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_59_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_187_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_59_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_188_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_58_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_186_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_58_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_187_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_57_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_185_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_57_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_186_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_56_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_184_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_56_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_185_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_55_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_183_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_55_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_184_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_54_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_182_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_54_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_183_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_53_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_181_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_53_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_182_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_52_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_180_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_52_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_181_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_51_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_179_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_51_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_180_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_50_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_178_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_50_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_179_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_49_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_177_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_49_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_178_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_48_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_176_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_48_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_177_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_47_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_175_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_47_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_176_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_46_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_174_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_46_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_175_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_45_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_173_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_45_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_174_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_44_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_172_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_44_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_173_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_43_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_171_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_43_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_172_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_42_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_170_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_42_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_171_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_41_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_169_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_41_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_170_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_40_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_168_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_40_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_169_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_39_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_167_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_39_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_168_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_38_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_166_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_38_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_167_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_37_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_165_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_37_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_166_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_36_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_164_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_36_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_165_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_35_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_163_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_35_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_164_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_34_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_162_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_34_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_163_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_33_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_161_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_33_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_162_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_32_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_160_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_32_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_161_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_31_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_159_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_31_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_160_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_30_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_158_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_30_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_159_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_29_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_157_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_29_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_158_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_28_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_156_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_28_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_157_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_27_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_155_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_27_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_156_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_26_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_154_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_26_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_155_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_25_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_153_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_25_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_154_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_24_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_152_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_24_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_153_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_23_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_151_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_23_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_152_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_22_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_150_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_22_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_151_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_21_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_149_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_21_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_150_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_20_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_148_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_20_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_149_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_19_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_147_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_19_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_148_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_18_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_146_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_18_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_147_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_17_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_145_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_17_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_146_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_16_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_144_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_16_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_145_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_15_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_143_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_15_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_144_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_14_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_142_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_14_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_143_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_13_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_141_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_13_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_142_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_12_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_140_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_12_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_141_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_11_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_139_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_11_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_140_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_10_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_138_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_10_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_139_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_9_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_137_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_9_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_138_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_8_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_136_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_8_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_137_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_7_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_135_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_7_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_136_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_6_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_134_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_6_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_135_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_5_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_133_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_5_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_134_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_4_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_132_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_4_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_133_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_3_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_131_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_3_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_132_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_2_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_130_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_2_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_131_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_1_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_129_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_1_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_130_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_0_sva_1
      & (input_write_addrs_lpi_1_dfm_2[7]) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_128_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_0_sva_1
      & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7])
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_129_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_127_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_127_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_127_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_128_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_126_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_126_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_126_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_127_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_125_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_125_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_125_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_126_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_124_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_124_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_124_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_125_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_123_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_123_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_123_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_124_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_122_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_122_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_122_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_123_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_121_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_121_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_121_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_122_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_120_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_120_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_120_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_121_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_119_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_119_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_119_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_120_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_118_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_118_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_118_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_119_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_117_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_117_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_117_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_118_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_116_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_116_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_116_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_117_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_115_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_115_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_115_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_116_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_114_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_114_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_114_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_115_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_113_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_113_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_113_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_114_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_112_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_112_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_112_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_113_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_111_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_111_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_111_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_112_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_110_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_110_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_110_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_111_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_109_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_109_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_109_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_110_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_108_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_108_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_108_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_109_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_107_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_107_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_107_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_108_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_106_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_106_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_106_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_107_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_105_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_105_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_105_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_106_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_104_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_104_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_104_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_105_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_103_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_103_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_103_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_104_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_102_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_102_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_102_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_103_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_101_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_101_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_101_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_102_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_100_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_100_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_100_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_101_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_99_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_99_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_99_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_100_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_98_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_98_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_98_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_99_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_97_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_97_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_97_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_98_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_96_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_96_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_96_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_97_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_95_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_95_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_95_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_96_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_94_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_94_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_94_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_95_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_93_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_93_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_93_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_94_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_92_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_92_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_92_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_93_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_91_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_91_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_91_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_92_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_90_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_90_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_90_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_91_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_89_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_89_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_89_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_90_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_88_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_88_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_88_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_89_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_87_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_87_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_87_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_88_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_86_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_86_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_86_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_87_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_85_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_85_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_85_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_86_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_84_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_84_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_84_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_85_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_83_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_83_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_83_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_84_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_82_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_82_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_82_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_83_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_81_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_81_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_81_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_82_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_80_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_80_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_80_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_81_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_79_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_79_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_79_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_80_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_78_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_78_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_78_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_79_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_77_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_77_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_77_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_78_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_76_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_76_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_76_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_77_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_75_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_75_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_75_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_76_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_74_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_74_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_74_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_75_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_73_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_73_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_73_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_74_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_72_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_72_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_72_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_73_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_71_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_71_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_71_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_72_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_70_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_70_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_70_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_71_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_69_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_69_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_69_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_70_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_68_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_68_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_68_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_69_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_67_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_67_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_67_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_68_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_66_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_66_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_66_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_67_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_65_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_65_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_65_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_66_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_64_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_64_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_64_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_65_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_63_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_63_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_63_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_64_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_62_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_62_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_62_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_63_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_61_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_61_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_61_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_62_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_60_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_60_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_60_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_61_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_59_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_59_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_59_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_60_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_58_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_58_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_58_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_59_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_57_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_57_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_57_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_58_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_56_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_56_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_56_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_57_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_55_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_55_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_55_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_56_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_54_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_54_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_54_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_55_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_53_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_53_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_53_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_54_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_52_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_52_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_52_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_53_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_51_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_51_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_51_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_52_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_50_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_50_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_50_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_51_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_49_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_49_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_49_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_50_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_48_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_48_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_48_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_49_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_47_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_47_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_47_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_48_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_46_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_46_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_46_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_47_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_45_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_45_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_45_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_46_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_44_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_44_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_44_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_45_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_43_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_43_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_43_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_44_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_42_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_42_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_42_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_43_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_41_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_41_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_41_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_42_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_40_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_40_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_40_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_41_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_39_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_39_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_39_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_40_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_38_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_38_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_38_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_39_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_37_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_37_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_37_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_38_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_36_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_36_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_36_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_37_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_35_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_35_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_35_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_36_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_34_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_34_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_34_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_35_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_33_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_33_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_33_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_34_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_32_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_32_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_32_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_33_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_31_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_31_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_31_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_32_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_30_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_30_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_30_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_31_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_29_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_29_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_29_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_30_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_28_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_28_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_28_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_29_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_27_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_27_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_27_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_28_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_26_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_26_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_26_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_27_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_25_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_25_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_25_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_26_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_24_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_24_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_24_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_25_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_23_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_23_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_23_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_24_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_22_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_22_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_22_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_23_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_21_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_21_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_21_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_22_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_20_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_20_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_20_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_21_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_19_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_19_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_19_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_20_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_18_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_18_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_18_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_19_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_17_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_17_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_17_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_18_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_16_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_16_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_16_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_17_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_15_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_15_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_15_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_16_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_14_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_14_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_14_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_15_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_13_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_13_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_13_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_14_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_12_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_12_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_12_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_13_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_11_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_11_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_11_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_12_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_10_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_10_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_10_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_11_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_9_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_9_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_9_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_10_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_8_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_8_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_8_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_9_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_7_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_7_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_7_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_8_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_6_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_6_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_6_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_7_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_5_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_5_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_5_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_6_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_4_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_4_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_4_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_5_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_3_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_3_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_3_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_4_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_2_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_2_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_2_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_3_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_1_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_1_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_1_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_write_arbxbar_xbar_1_for_3_if_1_and_2_tmp_1 = input_mem_banks_write_1_if_for_if_and_stg_6_0_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[7])) & input_write_req_valid_lpi_1_dfm_5;
  assign input_mem_write_arbxbar_xbar_for_3_if_1_and_tmp_1 = input_mem_banks_write_if_for_if_and_stg_6_0_sva_1
      & (~ (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7]))
      & input_write_req_valid_lpi_1_dfm_1_1;
  assign input_mem_banks_write_1_if_for_if_and_stg_5_0_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_0_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_1_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_1_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_2_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_2_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_3_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_3_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_4_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_4_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_5_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_5_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_6_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_6_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_7_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_7_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_8_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_8_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_9_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_9_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_10_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_10_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_11_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_11_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_12_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_12_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_13_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_13_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_14_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_14_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_15_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_15_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_16_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_16_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_17_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_17_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_18_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_18_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_19_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_19_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_20_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_20_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_21_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_21_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_22_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_22_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_23_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_23_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_24_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_24_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_25_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_25_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_26_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_26_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_27_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_27_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_28_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_28_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_29_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_29_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_30_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_30_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_31_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_31_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[5]));
  assign input_mem_banks_write_1_if_for_if_and_stg_5_32_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_0_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_33_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_1_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_34_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_2_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_35_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_3_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_36_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_4_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_37_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_5_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_38_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_6_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_39_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_7_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_40_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_8_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_41_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_9_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_42_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_10_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_43_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_11_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_44_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_12_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_45_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_13_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_46_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_14_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_47_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_15_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_48_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_16_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_49_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_17_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_50_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_18_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_51_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_19_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_52_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_20_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_53_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_21_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_54_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_22_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_55_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_23_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_56_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_24_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_57_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_25_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_58_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_26_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_59_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_27_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_60_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_28_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_61_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_29_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_62_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_30_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_5_63_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_4_31_sva_1
      & (input_write_addrs_lpi_1_dfm_2[5]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_0_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_0_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_1_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_1_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_2_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_2_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_3_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_3_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_4_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_4_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_5_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_5_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_6_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_6_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_7_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_7_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_8_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_8_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_9_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_9_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_10_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_10_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_11_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_11_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_12_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_12_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_13_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_13_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_14_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_14_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_15_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_15_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[4]));
  assign input_mem_banks_write_1_if_for_if_and_stg_4_16_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_0_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_17_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_1_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_18_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_2_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_19_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_3_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_20_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_4_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_21_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_5_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_22_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_6_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_23_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_7_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_24_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_8_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_25_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_9_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_26_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_10_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_27_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_11_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_28_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_12_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_29_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_13_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_30_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_14_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_4_31_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_3_15_sva_1
      & (input_write_addrs_lpi_1_dfm_2[4]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_0_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_0_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_1_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_1_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_2_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_2_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_3_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_3_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_4_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_4_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_5_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_5_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_6_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_6_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_7_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_7_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[3]));
  assign input_mem_banks_write_1_if_for_if_and_stg_3_8_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_0_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_9_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_1_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_10_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_2_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_11_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_3_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_12_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_4_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_13_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_5_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_14_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_6_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_3_15_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_2_7_sva_1
      & (input_write_addrs_lpi_1_dfm_2[3]);
  assign input_mem_banks_write_1_if_for_if_and_stg_2_0_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_0_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[2]));
  assign input_mem_banks_write_1_if_for_if_and_stg_2_1_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_1_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[2]));
  assign input_mem_banks_write_1_if_for_if_and_stg_2_2_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_2_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[2]));
  assign input_mem_banks_write_1_if_for_if_and_stg_2_3_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_3_sva_1
      & (~ (input_write_addrs_lpi_1_dfm_2[2]));
  assign input_mem_banks_write_1_if_for_if_and_stg_2_4_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_0_sva_1
      & (input_write_addrs_lpi_1_dfm_2[2]);
  assign input_mem_banks_write_1_if_for_if_and_stg_2_5_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_1_sva_1
      & (input_write_addrs_lpi_1_dfm_2[2]);
  assign input_mem_banks_write_1_if_for_if_and_stg_2_6_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_2_sva_1
      & (input_write_addrs_lpi_1_dfm_2[2]);
  assign input_mem_banks_write_1_if_for_if_and_stg_2_7_sva_1 = input_mem_banks_write_1_if_for_if_and_stg_1_3_sva_1
      & (input_write_addrs_lpi_1_dfm_2[2]);
  assign input_mem_banks_write_1_if_for_if_and_stg_1_0_sva_1 = ~((input_write_addrs_lpi_1_dfm_2[1:0]!=2'b00));
  assign input_mem_banks_write_1_if_for_if_and_stg_1_1_sva_1 = (input_write_addrs_lpi_1_dfm_2[1:0]==2'b01);
  assign input_mem_banks_write_1_if_for_if_and_stg_1_2_sva_1 = (input_write_addrs_lpi_1_dfm_2[1:0]==2'b10);
  assign input_mem_banks_write_1_if_for_if_and_stg_1_3_sva_1 = (input_write_addrs_lpi_1_dfm_2[1:0]==2'b11);
  assign PECore_DecodeAxiRead_case_4_switch_lp_nor_5_cse_1 = ~(PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_2
      | PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_2);
  assign PECore_DecodeAxiRead_switch_lp_equal_tmp_4 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:16]==4'b0011);
  assign PECore_DecodeAxiRead_switch_lp_nor_13_cse_1 = ~(PECore_DecodeAxiRead_switch_lp_equal_tmp_4
      | PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0 | PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0
      | PECore_DecodeAxiRead_switch_lp_nor_tmp_mx0w0);
  assign Arbiter_8U_Roundrobin_pick_1_if_1_not_185 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_2_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_1_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_1_idx_0_lpi_1_dfm_mx0
      & (~ operator_7_false_1_operator_7_false_1_or_mdf_sva_1);
  assign PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_and_5 =
      (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:16]==4'b0100);
  assign PECore_DecodeAxiRead_case_4_switch_lp_nor_6_tmp = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[15])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[14]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[13])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[12]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[10]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[9])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[8]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]));
  assign PECore_DecodeAxiRead_case_4_switch_lp_nor_8_tmp = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[15:1]!=15'b000000000000000));
  assign PECore_PushAxiRsp_if_asn_55 = (~ rva_in_reg_rw_sva_9) & PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_m1c_1;
  assign PECore_PushAxiRsp_if_asn_57 = rva_in_reg_rw_sva_9 & PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_m1c_1;
  assign PECore_PushAxiRsp_if_asn_59 = input_read_req_valid_lpi_1_dfm_1_9 & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7);
  assign weight_mem_run_3_for_5_asn_309 = (weight_read_addrs_7_lpi_1_dfm_3_2_0==3'b001)
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_asn_311 = (weight_read_addrs_7_lpi_1_dfm_3_2_0==3'b010)
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_asn_313 = (weight_read_addrs_7_lpi_1_dfm_3_2_0[2])
      & nor_894_cse & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_asn_315 = (weight_read_addrs_5_lpi_1_dfm_3_2_0==3'b001)
      & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_asn_317 = (weight_read_addrs_5_lpi_1_dfm_3_2_0==3'b010)
      & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_asn_319 = (weight_read_addrs_5_lpi_1_dfm_3_2_0[2])
      & nor_896_cse & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_118 = (weight_read_addrs_3_lpi_1_dfm_3_2_0==3'b001)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_120 = (weight_read_addrs_3_lpi_1_dfm_3_2_0==3'b010)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_122 = (weight_read_addrs_3_lpi_1_dfm_3_2_0==3'b100)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_asn_124 = (weight_read_addrs_3_lpi_1_dfm_3_2_0==3'b111)
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_3
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_4
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_5
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_6;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_1
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_2
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_5
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_6;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_2
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_4
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_6;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_3_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_1_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_0_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_3_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_3_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_1_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_0_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_5_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_3_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_1_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_0_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_7_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_3_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_1_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_0_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_9_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_3_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_1_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_0_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_11_6_mx0;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_asn_56 = (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[0])
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_cse & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_asn_321 = (weight_read_addrs_7_lpi_1_dfm_3_2_0==3'b111)
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_asn_323 = (weight_read_addrs_5_lpi_1_dfm_3_2_0==3'b111)
      & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_3_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_1_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_0_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_13_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_2 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_3_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_1 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_1_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_5_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_6_mx0;
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_0 = nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_0_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_2_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_4_mx0
      | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_15_6_mx0;
  assign PECore_PushAxiRsp_if_asn_61 = (~ rva_in_reg_rw_sva_5) & PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1;
  assign PECore_PushAxiRsp_if_asn_63 = rva_in_reg_rw_sva_5 & PECore_PushAxiRsp_if_PECore_PushAxiRsp_if_nor_2_m1c_1;
  assign PECore_PushAxiRsp_if_asn_65 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_11_itm_1
      & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign weight_mem_run_3_for_5_and_166 = weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_3_itm_1
      & weight_mem_run_3_for_land_4_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_98 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_7_itm_1
      & weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_and_168 = weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_12_itm_1
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_100 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_6_itm_2
      & weight_mem_run_3_for_land_2_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_and_172 = weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_5_itm_2
      & weight_mem_run_3_for_land_6_lpi_1_dfm_2;
  assign weight_mem_run_3_for_5_and_174 = weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_13_itm_2
      & weight_mem_run_3_for_land_lpi_1_dfm_2;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_and_52 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_80_itm_1
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_and_54 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_10_itm_1
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3;
  assign while_mux_1298_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_576_itm_1,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_600_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_5_6_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_391_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign while_mux_1285_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_600_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_36_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_601_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_4_1_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_323_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign while_mux_1283_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_601_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_34_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_602_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_4_2_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_322_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign while_mux_1282_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_602_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_33_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_603_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_4_3_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_321_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign while_mux_1281_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_603_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_32_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_604_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_4_4_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_320_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign while_mux_1280_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_604_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_31_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_605_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_4_5_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_319_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign while_mux_1279_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_605_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_30_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_606_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_4_6_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_318_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign while_mux_1278_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_606_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_29_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign while_mux_1277_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_350_itm_1,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_607_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_3_1_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_250_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign while_mux_1276_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_607_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_27_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_608_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_3_2_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_249_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign while_mux_1275_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_608_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_26_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_609_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_3_3_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_248_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign while_mux_1274_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_609_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_25_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_610_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_3_4_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_247_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign while_mux_1273_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_610_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_24_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_611_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_3_5_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_246_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign while_mux_1272_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_611_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_23_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_612_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_3_6_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_245_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1);
  assign while_mux_1271_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_612_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_22_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign while_mux_1270_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_277_itm_1,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_613_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_2_1_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_177_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign while_mux_1269_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_613_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_20_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_614_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_2_2_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_176_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign while_mux_1268_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_614_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_19_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_615_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_2_3_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_175_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign while_mux_1267_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_615_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_18_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_616_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_2_4_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_174_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign while_mux_1266_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_616_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_17_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_617_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_2_5_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_173_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign while_mux_1265_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_617_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_16_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_618_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_2_6_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_172_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1);
  assign while_mux_1264_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_618_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_15_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign while_mux_1263_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_204_itm_1,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_619_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_1_1_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_104_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign while_mux_1262_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_619_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_13_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_620_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_1_2_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_103_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign while_mux_1261_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_620_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_12_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_621_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_1_3_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_102_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign while_mux_1260_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_621_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_11_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_622_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_1_4_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_101_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign while_mux_1259_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_622_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_10_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_623_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_1_5_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_100_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign while_mux_1258_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_623_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_9_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_624_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_1_6_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_99_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1);
  assign while_mux_1257_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_624_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_8_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign while_mux_1256_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_131_itm_1,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_629_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_0_5_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_27_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1);
  assign while_mux_1251_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_629_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_2_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign Arbiter_8U_Roundrobin_pick_1_mux_630_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_0_6_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_26_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1);
  assign while_mux_1250_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_630_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_1_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign while_mux_1249_tmp = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_57_itm_1,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_dcpl_4 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8
      & while_stage_0_10;
  assign and_dcpl_5 = and_dcpl_4 & (~ rva_in_reg_rw_sva_st_1_8);
  assign and_dcpl_6 = and_dcpl_5 & (~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6
      | rva_in_reg_rw_sva_8 | input_read_req_valid_lpi_1_dfm_1_8));
  assign and_dcpl_27 = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7)
      & while_stage_0_9;
  assign and_dcpl_31 = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
      & PECore_RunMac_PECore_RunMac_if_and_svs_st_5 & while_stage_0_7;
  assign and_dcpl_32 = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
      & while_stage_0_7;
  assign or_tmp_2 = (~ PECore_RunMac_PECore_RunMac_if_and_svs_st_5) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
  assign or_tmp_3 = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
      | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3;
  assign and_dcpl_40 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & while_stage_0_6;
  assign and_dcpl_41 = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      & while_stage_0_6;
  assign or_tmp_4 = rva_in_reg_rw_sva_st_1_4 | rva_in_reg_rw_sva_4 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_17_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2;
  assign and_tmp = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & or_tmp_4;
  assign or_tmp_5 = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      | rva_in_reg_rw_sva_st_1_4 | rva_in_reg_rw_sva_4 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_17_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2;
  assign nor_tmp_1 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_95_itm_1
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2;
  assign and_dcpl_69 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      & while_stage_0_5;
  assign and_dcpl_78 = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign and_dcpl_79 = and_dcpl_78 & weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp;
  assign and_dcpl_80 = and_dcpl_78 & weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp;
  assign and_dcpl_82 = weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign and_dcpl_84 = weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign and_dcpl_86 = weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign and_dcpl_88 = weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign and_dcpl_90 = weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign and_dcpl_92 = weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign or_dcpl_13 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      | (~ while_stage_0_4);
  assign nor_227_cse = ~((weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]));
  assign and_100_cse = (~((weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]) |
      (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]))) & (~((weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]))) & (~((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]))) & nor_227_cse;
  assign nor_230_cse = ~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]));
  assign nor_231_cse = ~((weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]));
  assign nor_228_cse = ~((weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]));
  assign nor_229_cse = ~((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]));
  assign and_114_cse = (~((weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[5]) |
      (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5]))) & (~((weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[5]))) & (~((weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[5]))) & (~((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5])));
  assign or_dcpl_16 = and_114_cse | or_dcpl_13;
  assign nor_238_cse = ~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]));
  assign nor_239_cse = ~((weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4]));
  assign nor_236_cse = ~((weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4]));
  assign nor_237_cse = ~((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[4]) | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[4]));
  assign nor_242_cse = ~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]));
  assign nor_243_cse = ~((weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3]));
  assign nor_240_cse = ~((weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[3]));
  assign nor_241_cse = ~((weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[3]) | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[3]));
  assign nor_246_cse = ~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]));
  assign nor_247_cse = ~((weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2]));
  assign nor_244_cse = ~((weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]));
  assign nor_245_cse = ~((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[2]) | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2]));
  assign nor_250_cse = ~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]));
  assign nor_251_cse = ~((weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1]));
  assign nor_248_cse = ~((weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1]));
  assign nor_249_cse = ~((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1]) | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]));
  assign and_149_cse = (~((weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[0]) |
      (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[0]))) & (~((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0]))) & (~((weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0]))) & (~((weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0])));
  assign or_dcpl_21 = and_149_cse | or_dcpl_13;
  assign and_dcpl_149 = (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5])) & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[5]);
  assign and_dcpl_150 = (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4])) & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[4]);
  assign and_dcpl_151 = (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[0])) & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[0]);
  assign and_dcpl_152 = (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3])) & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[3]);
  assign and_dcpl_153 = (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[2])) & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[2]);
  assign and_dcpl_154 = (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1])) & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[1]);
  assign and_dcpl_155 = (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7])) & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[7]);
  assign and_dcpl_156 = (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6])) & (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[6]);
  assign and_dcpl_162 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4;
  assign and_dcpl_168 = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2)
      & while_stage_0_4;
  assign and_dcpl_178 = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4;
  assign and_dcpl_179 = and_dcpl_151 & and_dcpl_162;
  assign and_dcpl_181 = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1]) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4;
  assign and_dcpl_182 = and_dcpl_154 & and_dcpl_162;
  assign and_dcpl_184 = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[2]) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4;
  assign and_dcpl_185 = and_dcpl_153 & and_dcpl_162;
  assign and_dcpl_187 = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3]) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4;
  assign and_dcpl_188 = and_dcpl_152 & and_dcpl_162;
  assign and_dcpl_190 = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4]) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4;
  assign and_dcpl_191 = and_dcpl_150 & and_dcpl_162;
  assign and_dcpl_193 = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5]) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4;
  assign and_dcpl_194 = and_dcpl_149 & and_dcpl_162;
  assign and_dcpl_196 = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6]) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4;
  assign and_dcpl_197 = and_dcpl_156 & and_dcpl_162;
  assign and_dcpl_199 = (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7]) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      & while_stage_0_4;
  assign and_dcpl_200 = and_dcpl_155 & and_dcpl_162;
  assign and_dcpl_203 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      & while_stage_0_3;
  assign and_dcpl_204 = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      & while_stage_0_3;
  assign and_dcpl_207 = nor_340_cse & (state_2_1_sva[0]) & and_dcpl_204;
  assign or_120_nl = nor_340_cse | PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva;
  assign and_691_nl = or_2088_cse & PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva;
  assign or_117_nl = (~ input_port_PopNB_mioi_return_rsc_z_mxwt) | (state_2_1_sva[0]);
  assign mux_19_nl = MUX_s_1_2_2(or_120_nl, and_691_nl, or_117_nl);
  assign and_dcpl_209 = mux_19_nl & and_dcpl_204 & (~ PECore_RunFSM_switch_lp_nor_tmp_1);
  assign or_dcpl_87 = ~(rva_in_PopNB_mioi_return_rsc_z_mxwt & reg_rva_in_PopNB_mioi_iswt0_cse);
  assign and_dcpl_210 = (~ rva_in_PopNB_mioi_return_rsc_z_mxwt) & reg_rva_in_PopNB_mioi_iswt0_cse;
  assign or_dcpl_91 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:18]!=2'b01);
  assign and_dcpl_211 = reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  assign and_dcpl_215 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_return_rsc_z_mxwt;
  assign and_dcpl_216 = and_dcpl_215 & and_dcpl_211 & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]);
  assign and_dcpl_217 = reg_rva_in_PopNB_mioi_iswt0_cse & (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt);
  assign and_dcpl_219 = and_dcpl_215 & and_dcpl_217 & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]);
  assign and_dcpl_221 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7
      & (~ rva_in_reg_rw_sva_st_1_7);
  assign or_tmp_33 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
      | PECore_RunMac_PECore_RunMac_if_and_svs_st_2;
  assign and_692_cse = rva_in_PopNB_mioi_return_rsc_z_mxwt & reg_rva_in_PopNB_mioi_iswt0_cse;
  assign and_dcpl_228 = crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4;
  assign and_dcpl_241 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      & while_stage_0_7;
  assign and_dcpl_242 = and_692_cse & (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt);
  assign and_dcpl_246 = PECore_RunMac_PECore_RunMac_if_and_svs_st_3 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign and_dcpl_248 = PECore_RunFSM_switch_lp_equal_tmp_1_2 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3)
      & while_stage_0_5;
  assign and_dcpl_266 = and_dcpl_221 & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5);
  assign and_696_nl = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1 & Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_3
      & PECore_RunFSM_switch_lp_equal_tmp_1_2;
  assign mux_28_nl = MUX_s_1_2_2(and_696_nl, PECore_RunFSM_switch_lp_equal_tmp_1_2,
      Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_2_tmp);
  assign or_187_nl = Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_22_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_26_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_14_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_10_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_6_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_18_tmp;
  assign mux_tmp_25 = MUX_s_1_2_2(mux_28_nl, PECore_RunFSM_switch_lp_equal_tmp_1_2,
      or_187_nl);
  assign or_tmp_43 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~ mux_tmp_25);
  assign and_dcpl_281 = and_dcpl_221 & while_stage_0_9;
  assign and_dcpl_282 = ~(rva_in_reg_rw_sva_7 | input_read_req_valid_lpi_1_dfm_1_7);
  assign and_dcpl_293 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6
      & (~ rva_in_reg_rw_sva_st_1_6);
  assign and_dcpl_294 = and_dcpl_293 & (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_4);
  assign or_tmp_206 = (~(rva_in_reg_rw_sva_st_1_4 | rva_in_reg_rw_sva_4 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_17_itm_1))
      | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2;
  assign nor_288_nl = ~((~ weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1)
      | weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
  assign nor_289_nl = ~((~(weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | (~ weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1)))
      | weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
  assign or_365_nl = (~(weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1))
      | weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
  assign not_tmp_203 = MUX_s_1_2_2(nor_288_nl, nor_289_nl, or_365_nl);
  assign or_tmp_215 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | not_tmp_203;
  assign nor_290_nl = ~(weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | not_tmp_203);
  assign mux_tmp_108 = MUX_s_1_2_2(nor_290_nl, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign and_dcpl_312 = nor_536_cse & and_692_cse;
  assign not_tmp_217 = ~(crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1_1
      | reg_rva_in_reg_rw_sva_2_cse);
  assign and_dcpl_329 = ~(input_read_req_valid_lpi_1_dfm_1_6 | rva_in_reg_rw_sva_6);
  assign and_dcpl_355 = while_and_23_cse & while_stage_0_7;
  assign nand_27_cse = ~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      & while_stage_0_7);
  assign and_dcpl_376 = ~(pe_manager_base_weight_slc_pe_manager_base_weight_2_0_178_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1);
  assign or_tmp_334 = rva_in_reg_rw_sva_3 | input_read_req_valid_lpi_1_dfm_1_3 |
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1 | pe_manager_base_weight_slc_pe_manager_base_weight_2_0_178_itm_1;
  assign and_dcpl_389 = and_dcpl_376 & (~ input_read_req_valid_lpi_1_dfm_1_3);
  assign and_dcpl_398 = (~ reg_rva_in_reg_rw_sva_2_cse) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2;
  assign nor_320_cse = ~(reg_rva_in_reg_rw_sva_2_cse | accum_vector_operator_1_for_asn_7_itm_1);
  assign and_dcpl_401 = ((~ weight_mem_run_1_if_for_weight_mem_run_1_if_for_weight_mem_run_1_if_for_nor_tmp)
      | crossbar_spec_PE_Weight_WordType_8U_8U_for_mux_1_tmp) & nor_320_cse;
  assign and_dcpl_419 = ~(reg_rva_in_reg_rw_sva_st_1_1_cse | ProductSum_for_asn_64_itm_1);
  assign and_dcpl_420 = and_dcpl_419 & and_dcpl_203;
  assign mux_tmp_182 = ~(reg_rva_in_reg_rw_sva_st_1_1_cse | (while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1!=4'b0100));
  assign and_dcpl_431 = ~(reg_rva_in_reg_rw_sva_st_1_1_cse | ProductSum_for_asn_64_itm_1
      | (while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1[0]));
  assign nand_36_cse = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]) & PECore_DecodeAxiRead_case_4_switch_lp_nor_6_tmp);
  assign and_dcpl_459 = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6)
      & PECore_RunMac_PECore_RunMac_if_and_svs_st_6 & while_stage_0_8;
  assign and_dcpl_467 = and_dcpl_69 & ProductSum_for_asn_73_itm_3;
  assign or_tmp_341 = weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_2
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_54_itm_1;
  assign or_tmp_342 = (~ weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2)
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
  assign nor_360_nl = ~(weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign mux_187_nl = MUX_s_1_2_2(or_tmp_342, nor_360_nl, weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_3);
  assign mux_188_itm = MUX_s_1_2_2(mux_187_nl, or_tmp_342, weight_mem_run_3_for_5_and_108_itm_1);
  assign and_dcpl_469 = and_dcpl_69 & ProductSum_for_asn_64_itm_3;
  assign or_tmp_347 = weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_2
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_44_itm_1;
  assign nor_361_nl = ~(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_7_itm_1
      | (~ weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_3));
  assign not_tmp_312 = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2,
      nor_361_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign or_tmp_352 = (~ weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_2)
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_35_itm_1;
  assign not_tmp_314 = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1,
      (~ or_tmp_352), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign or_tmp_358 = (~ weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_2)
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_34_itm_1;
  assign not_tmp_316 = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1,
      (~ or_tmp_358), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign or_tmp_364 = PECore_RunScale_PECore_RunScale_if_and_1_svs_st_3 | ProductSum_for_asn_25_itm_3;
  assign or_tmp_365 = (~ reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_3_1_itm_2_cse)
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_1;
  assign not_tmp_319 = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1,
      (~ or_tmp_365), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign not_tmp_322 = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1,
      nor_17_cse, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign not_tmp_325 = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1,
      nor_18_cse, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign or_tmp_382 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | (~ weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
  assign mux_229_nl = MUX_s_1_2_2(or_tmp_382, nor_469_cse, reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_0_1_itm_2_cse);
  assign mux_230_itm = MUX_s_1_2_2(mux_229_nl, or_tmp_382, crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_19_itm_1);
  assign and_704_cse = PECore_UpdateFSM_switch_lp_and_7_itm_1 & pe_config_is_valid_sva;
  assign or_dcpl_603 = reg_PECore_RunMac_PECore_RunMac_if_and_svs_st_8_cse | (~ PECore_RunScale_PECore_RunScale_if_and_1_svs_8);
  assign and_dcpl_504 = weight_mem_run_3_for_land_2_lpi_1_dfm_2 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign and_dcpl_505 = ~(weight_mem_run_3_for_land_2_lpi_1_dfm_2 | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign or_dcpl_606 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      | (~ while_stage_0_7);
  assign and_dcpl_525 = and_dcpl_78 & (~ while_stage_0_4);
  assign or_dcpl_615 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~ while_stage_0_5);
  assign and_dcpl_529 = nor_230_cse & nor_231_cse;
  assign and_dcpl_532 = nor_228_cse & nor_229_cse;
  assign and_dcpl_533 = and_dcpl_532 & and_dcpl_529;
  assign and_dcpl_543 = nor_238_cse & nor_239_cse;
  assign and_dcpl_547 = nor_236_cse & nor_237_cse & and_dcpl_543;
  assign and_dcpl_550 = nor_242_cse & nor_243_cse;
  assign and_dcpl_554 = nor_240_cse & nor_241_cse & and_dcpl_550;
  assign and_dcpl_557 = nor_246_cse & nor_247_cse;
  assign and_dcpl_561 = nor_244_cse & nor_245_cse & and_dcpl_557;
  assign and_dcpl_564 = nor_250_cse & nor_251_cse;
  assign and_dcpl_568 = nor_248_cse & nor_249_cse & and_dcpl_564;
  assign or_dcpl_616 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
      | (~ while_stage_0_3);
  assign or_dcpl_627 = or_dcpl_87 | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt);
  assign or_dcpl_628 = or_dcpl_91 | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]);
  assign or_dcpl_632 = or_2088_cse | (state_2_1_sva[0]);
  assign or_dcpl_635 = (~ while_stage_0_11) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_9;
  assign or_dcpl_658 = (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])
      | nand_36_cse;
  assign and_dcpl_580 = crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2
      & (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0]);
  assign and_dcpl_582 = crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2
      & (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1:0]==2'b10);
  assign and_dcpl_584 = crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2
      & (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1:0]==2'b00);
  assign and_dcpl_588 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & (~ (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1]));
  assign and_dcpl_592 = ~(weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
  assign or_dcpl_665 = (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6)
      | rva_in_reg_rw_sva_6 | (~ while_stage_0_8);
  assign and_dcpl_611 = (~(rva_in_PopNB_mioi_return_rsc_z_mxwt | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
      & while_stage_0_3;
  assign and_dcpl_612 = or_dcpl_616 & (~ rva_in_PopNB_mioi_return_rsc_z_mxwt);
  assign or_1079_nl = while_stage_0_3 | (state_2_1_sva!=2'b01) | state_0_sva;
  assign or_1078_nl = (state_2_1_sva!=2'b01) | state_0_sva;
  assign mux_269_nl = MUX_s_1_2_2(or_1078_nl, mux_246_cse, while_stage_0_3);
  assign nor_27_nl = ~((state_2_1_sva_dfm_1!=2'b01));
  assign mux_270_nl = MUX_s_1_2_2(or_1079_nl, mux_269_nl, nor_27_nl);
  assign and_dcpl_616 = (~ mux_270_nl) & and_dcpl_210;
  assign nor_tmp_39 = weight_mem_read_arbxbar_arbiters_next_7_6_sva & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]);
  assign and_714_cse = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]) & weight_mem_read_arbxbar_arbiters_next_7_5_sva;
  assign or_tmp_415 = and_714_cse | nor_tmp_39;
  assign nor_tmp_41 = Arbiter_8U_Roundrobin_pick_1_mux_537_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]);
  assign and_716_cse = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]) & Arbiter_8U_Roundrobin_pick_1_mux_538_itm_1;
  assign or_1099_cse = and_716_cse | nor_tmp_41;
  assign mux_280_nl = MUX_s_1_2_2(or_tmp_415, or_1099_cse, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1);
  assign or_1097_nl = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]);
  assign mux_279_nl = MUX_s_1_2_2(or_tmp_415, or_1097_nl, weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign mux_tmp_277 = MUX_s_1_2_2(mux_280_nl, mux_279_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_283_nl = MUX_s_1_2_2(or_tmp_415, mux_tmp_277, while_stage_0_5);
  assign or_1101_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1
      | or_tmp_415;
  assign or_1100_nl = while_mux_1298_tmp | mux_tmp_277;
  assign mux_282_nl = MUX_s_1_2_2(or_1101_nl, or_1100_nl, while_stage_0_5);
  assign mux_tmp_280 = MUX_s_1_2_2(mux_283_nl, mux_282_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]);
  assign and_720_cse = weight_mem_read_arbxbar_arbiters_next_7_3_sva & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]);
  assign and_721_cse = weight_mem_read_arbxbar_arbiters_next_7_2_sva & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]);
  assign and_722_cse = weight_mem_read_arbxbar_arbiters_next_7_1_sva & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7]);
  assign nand_1_nl = ~(weight_mem_read_arbxbar_arbiters_next_7_4_sva & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7])
      & (~ or_tmp_415));
  assign mux_285_nl = MUX_s_1_2_2(nand_1_nl, or_tmp_415, and_720_cse);
  assign mux_286_nl = MUX_s_1_2_2(mux_285_nl, or_tmp_415, and_721_cse);
  assign mux_tmp_283 = MUX_s_1_2_2(mux_286_nl, or_tmp_415, and_722_cse);
  assign and_728_cse = Arbiter_8U_Roundrobin_pick_1_mux_540_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]);
  assign and_729_cse = Arbiter_8U_Roundrobin_pick_1_mux_541_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]);
  assign and_730_cse = Arbiter_8U_Roundrobin_pick_1_mux_542_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7]);
  assign nor_404_nl = ~((Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7])) | mux_tmp_283);
  assign nand_2_nl = ~(Arbiter_8U_Roundrobin_pick_1_mux_539_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7])
      & (~ or_1099_cse));
  assign mux_289_nl = MUX_s_1_2_2(nand_2_nl, or_1099_cse, and_728_cse);
  assign mux_290_nl = MUX_s_1_2_2(mux_289_nl, or_1099_cse, and_729_cse);
  assign mux_291_nl = MUX_s_1_2_2(mux_290_nl, or_1099_cse, and_730_cse);
  assign mux_292_nl = MUX_s_1_2_2(mux_tmp_283, mux_291_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1);
  assign or_1103_nl = (~((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7])))
      | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]);
  assign mux_288_nl = MUX_s_1_2_2(mux_tmp_283, or_1103_nl, weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign mux_293_nl = MUX_s_1_2_2(mux_292_nl, mux_288_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign nor_405_nl = ~((while_mux_1298_tmp & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]))
      | mux_293_nl);
  assign not_tmp_469 = MUX_s_1_2_2(nor_404_nl, nor_405_nl, while_stage_0_5);
  assign and_732_cse = weight_mem_read_arbxbar_arbiters_next_7_4_sva & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]);
  assign or_tmp_427 = and_720_cse | and_732_cse | nor_tmp_39;
  assign or_tmp_430 = and_721_cse | and_722_cse | and_714_cse | or_tmp_427;
  assign and_737_cse = Arbiter_8U_Roundrobin_pick_1_mux_539_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]);
  assign or_tmp_432 = and_728_cse | and_737_cse | nor_tmp_41;
  assign or_1118_nl = and_729_cse | and_730_cse | and_716_cse | or_tmp_432;
  assign mux_296_nl = MUX_s_1_2_2(or_tmp_430, or_1118_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1);
  assign or_1108_nl = (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]) | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]);
  assign mux_295_nl = MUX_s_1_2_2(or_tmp_430, or_1108_nl, weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7]);
  assign mux_tmp_293 = MUX_s_1_2_2(mux_296_nl, mux_295_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign or_1120_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1
      | or_tmp_430;
  assign or_1119_nl = while_mux_1298_tmp | mux_tmp_293;
  assign mux_tmp_294 = MUX_s_1_2_2(or_1120_nl, or_1119_nl, while_stage_0_5);
  assign mux_tmp_295 = MUX_s_1_2_2(or_tmp_430, mux_tmp_293, while_stage_0_5);
  assign or_1124_nl = and_720_cse | and_732_cse | weight_mem_read_arbxbar_arbiters_next_7_6_sva
      | (~ (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]));
  assign or_1121_nl = weight_mem_read_arbxbar_arbiters_next_7_5_sva | or_tmp_427;
  assign mux_300_nl = MUX_s_1_2_2(or_1124_nl, or_1121_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]);
  assign or_tmp_443 = and_721_cse | and_722_cse | mux_300_nl;
  assign or_1131_nl = and_728_cse | and_737_cse | Arbiter_8U_Roundrobin_pick_1_mux_537_itm_1
      | (~ (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7]));
  assign or_1128_nl = Arbiter_8U_Roundrobin_pick_1_mux_538_itm_1 | or_tmp_432;
  assign mux_301_nl = MUX_s_1_2_2(or_1131_nl, or_1128_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]);
  assign or_1133_nl = and_729_cse | and_730_cse | mux_301_nl;
  assign mux_302_nl = MUX_s_1_2_2(or_tmp_443, or_1133_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1);
  assign or_1127_nl = (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7])
      | or_tmp_443;
  assign mux_303_nl = MUX_s_1_2_2(mux_302_nl, or_1127_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_304_nl = MUX_s_1_2_2(or_tmp_443, mux_303_nl, while_stage_0_5);
  assign mux_305_nl = MUX_s_1_2_2(mux_304_nl, mux_tmp_295, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[7]);
  assign mux_306_itm = MUX_s_1_2_2(mux_305_nl, mux_tmp_294, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[7]);
  assign or_tmp_451 = and_720_cse | and_732_cse;
  assign or_1139_nl = weight_mem_read_arbxbar_arbiters_next_7_4_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]));
  assign or_1138_nl = weight_mem_read_arbxbar_arbiters_next_7_3_sva | and_732_cse;
  assign mux_307_nl = MUX_s_1_2_2(or_1139_nl, or_1138_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]);
  assign or_1137_nl = weight_mem_read_arbxbar_arbiters_next_7_1_sva | or_tmp_451;
  assign mux_308_nl = MUX_s_1_2_2(mux_307_nl, or_1137_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7]);
  assign or_1136_nl = weight_mem_read_arbxbar_arbiters_next_7_2_sva | and_722_cse
      | or_tmp_451;
  assign mux_tmp_305 = MUX_s_1_2_2(mux_308_nl, or_1136_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]);
  assign or_tmp_458 = and_728_cse | and_737_cse;
  assign or_1146_nl = Arbiter_8U_Roundrobin_pick_1_mux_539_itm_1 | (~ (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[7]));
  assign or_1145_nl = Arbiter_8U_Roundrobin_pick_1_mux_540_itm_1 | and_737_cse;
  assign mux_310_nl = MUX_s_1_2_2(or_1146_nl, or_1145_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[7]);
  assign or_1144_nl = Arbiter_8U_Roundrobin_pick_1_mux_542_itm_1 | or_tmp_458;
  assign mux_311_nl = MUX_s_1_2_2(mux_310_nl, or_1144_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[7]);
  assign or_1143_nl = Arbiter_8U_Roundrobin_pick_1_mux_541_itm_1 | and_730_cse |
      or_tmp_458;
  assign mux_312_nl = MUX_s_1_2_2(mux_311_nl, or_1143_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[7]);
  assign mux_313_nl = MUX_s_1_2_2(mux_tmp_305, mux_312_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1);
  assign or_1140_nl = (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[7])
      | mux_tmp_305;
  assign mux_314_nl = MUX_s_1_2_2(mux_313_nl, or_1140_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_315_nl = MUX_s_1_2_2(mux_tmp_305, mux_314_nl, while_stage_0_5);
  assign and_dcpl_625 = (~ mux_315_nl) & (~((weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[7])
      | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[7]))) & nor_227_cse;
  assign and_755_cse = (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]) & weight_mem_read_arbxbar_arbiters_next_6_6_sva;
  assign and_756_cse = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6]) & weight_mem_read_arbxbar_arbiters_next_6_5_sva;
  assign or_tmp_465 = and_755_cse | and_756_cse;
  assign or_1147_nl = (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6]);
  assign mux_tmp_313 = MUX_s_1_2_2(or_tmp_465, or_1147_nl, weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[6]);
  assign and_757_cse = (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]) & Arbiter_8U_Roundrobin_pick_1_mux_464_itm_1;
  assign and_758_cse = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6]) & Arbiter_8U_Roundrobin_pick_1_mux_465_itm_1;
  assign or_1150_nl = and_757_cse | and_758_cse;
  assign mux_tmp_314 = MUX_s_1_2_2(or_tmp_465, or_1150_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign mux_321_nl = MUX_s_1_2_2(mux_tmp_314, mux_tmp_313, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_322_nl = MUX_s_1_2_2(or_tmp_465, mux_321_nl, while_stage_0_5);
  assign or_1152_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1
      | or_tmp_465;
  assign or_1151_nl = Arbiter_8U_Roundrobin_pick_1_mux_496_itm_1 | mux_tmp_314;
  assign or_1149_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1
      | mux_tmp_313;
  assign mux_319_nl = MUX_s_1_2_2(or_1151_nl, or_1149_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_320_nl = MUX_s_1_2_2(or_1152_nl, mux_319_nl, while_stage_0_5);
  assign mux_tmp_319 = MUX_s_1_2_2(mux_322_nl, mux_320_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]);
  assign nor_tmp_89 = weight_mem_read_arbxbar_arbiters_next_6_3_sva & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]);
  assign or_tmp_472 = ((weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]) & weight_mem_read_arbxbar_arbiters_next_6_4_sva)
      | nor_tmp_89;
  assign or_tmp_473 = ((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6]) & weight_mem_read_arbxbar_arbiters_next_6_1_sva)
      | or_tmp_472;
  assign or_tmp_474 = ((weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]) & weight_mem_read_arbxbar_arbiters_next_6_2_sva)
      | or_tmp_473;
  assign or_tmp_476 = and_755_cse | (~((~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6])
      & weight_mem_read_arbxbar_arbiters_next_6_5_sva)) & or_tmp_474));
  assign or_1154_nl = (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6])
      | and_dcpl_532;
  assign mux_tmp_320 = MUX_s_1_2_2(or_tmp_476, or_1154_nl, weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[6]);
  assign nor_tmp_95 = Arbiter_8U_Roundrobin_pick_1_mux_467_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]);
  assign or_tmp_478 = ((weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]) & Arbiter_8U_Roundrobin_pick_1_mux_466_itm_1)
      | nor_tmp_95;
  assign or_tmp_479 = ((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6]) & Arbiter_8U_Roundrobin_pick_1_mux_469_itm_1)
      | or_tmp_478;
  assign or_tmp_480 = ((weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]) & Arbiter_8U_Roundrobin_pick_1_mux_468_itm_1)
      | or_tmp_479;
  assign or_1165_nl = and_757_cse | (~((~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6])
      & Arbiter_8U_Roundrobin_pick_1_mux_465_itm_1)) & or_tmp_480));
  assign mux_tmp_321 = MUX_s_1_2_2(or_tmp_476, or_1165_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign mux_328_nl = MUX_s_1_2_2(mux_tmp_321, mux_tmp_320, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_329_nl = MUX_s_1_2_2(or_tmp_476, mux_328_nl, while_stage_0_5);
  assign or_1167_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1
      | or_tmp_476;
  assign or_1166_nl = Arbiter_8U_Roundrobin_pick_1_mux_496_itm_1 | mux_tmp_321;
  assign or_1160_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1
      | mux_tmp_320;
  assign mux_326_nl = MUX_s_1_2_2(or_1166_nl, or_1160_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_327_nl = MUX_s_1_2_2(or_1167_nl, mux_326_nl, while_stage_0_5);
  assign mux_330_itm = MUX_s_1_2_2(mux_329_nl, mux_327_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]);
  assign or_tmp_486 = and_756_cse | or_tmp_474;
  assign or_tmp_487 = and_755_cse | or_tmp_486;
  assign or_1168_nl = (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6])
      | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]) | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]);
  assign mux_tmp_327 = MUX_s_1_2_2(or_tmp_487, or_1168_nl, weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[6]);
  assign or_tmp_489 = and_758_cse | or_tmp_480;
  assign or_1173_nl = and_757_cse | or_tmp_489;
  assign mux_tmp_328 = MUX_s_1_2_2(or_tmp_487, or_1173_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign or_1175_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1
      | or_tmp_487;
  assign or_1174_nl = Arbiter_8U_Roundrobin_pick_1_mux_496_itm_1 | mux_tmp_328;
  assign or_1171_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1
      | mux_tmp_327;
  assign mux_333_nl = MUX_s_1_2_2(or_1174_nl, or_1171_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_tmp_330 = MUX_s_1_2_2(or_1175_nl, mux_333_nl, while_stage_0_5);
  assign mux_335_nl = MUX_s_1_2_2(mux_tmp_328, mux_tmp_327, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_tmp_332 = MUX_s_1_2_2(or_tmp_487, mux_335_nl, while_stage_0_5);
  assign or_1178_nl = (~ (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6])) |
      weight_mem_read_arbxbar_arbiters_next_6_5_sva | or_tmp_474;
  assign or_1176_nl = weight_mem_read_arbxbar_arbiters_next_6_6_sva | or_tmp_486;
  assign mux_tmp_333 = MUX_s_1_2_2(or_1178_nl, or_1176_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]);
  assign or_1182_nl = (~ (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[6])) |
      Arbiter_8U_Roundrobin_pick_1_mux_465_itm_1 | or_tmp_480;
  assign or_1180_nl = Arbiter_8U_Roundrobin_pick_1_mux_464_itm_1 | or_tmp_489;
  assign mux_338_nl = MUX_s_1_2_2(or_1182_nl, or_1180_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[6]);
  assign mux_339_nl = MUX_s_1_2_2(mux_tmp_333, mux_338_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign or_1179_nl = (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[6])
      | mux_tmp_333;
  assign mux_340_nl = MUX_s_1_2_2(mux_339_nl, or_1179_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_341_nl = MUX_s_1_2_2(mux_tmp_333, mux_340_nl, while_stage_0_5);
  assign mux_342_nl = MUX_s_1_2_2(mux_341_nl, mux_tmp_332, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[6]);
  assign mux_343_itm = MUX_s_1_2_2(mux_342_nl, mux_tmp_330, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[6]);
  assign or_1186_nl = weight_mem_read_arbxbar_arbiters_next_6_3_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]));
  assign or_1185_nl = weight_mem_read_arbxbar_arbiters_next_6_4_sva | nor_tmp_89;
  assign mux_344_nl = MUX_s_1_2_2(or_1186_nl, or_1185_nl, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]);
  assign or_1184_nl = weight_mem_read_arbxbar_arbiters_next_6_1_sva | or_tmp_472;
  assign mux_345_nl = MUX_s_1_2_2(mux_344_nl, or_1184_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6]);
  assign or_1183_nl = weight_mem_read_arbxbar_arbiters_next_6_2_sva | or_tmp_473;
  assign mux_tmp_342 = MUX_s_1_2_2(mux_345_nl, or_1183_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]);
  assign or_1191_nl = Arbiter_8U_Roundrobin_pick_1_mux_467_itm_1 | (~ (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[6]));
  assign or_1190_nl = Arbiter_8U_Roundrobin_pick_1_mux_466_itm_1 | nor_tmp_95;
  assign mux_347_nl = MUX_s_1_2_2(or_1191_nl, or_1190_nl, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[6]);
  assign or_1189_nl = Arbiter_8U_Roundrobin_pick_1_mux_469_itm_1 | or_tmp_478;
  assign mux_348_nl = MUX_s_1_2_2(mux_347_nl, or_1189_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[6]);
  assign or_1188_nl = Arbiter_8U_Roundrobin_pick_1_mux_468_itm_1 | or_tmp_479;
  assign mux_349_nl = MUX_s_1_2_2(mux_348_nl, or_1188_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[6]);
  assign mux_350_nl = MUX_s_1_2_2(mux_tmp_342, mux_349_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign or_1187_nl = (weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[6])
      | mux_tmp_342;
  assign mux_351_nl = MUX_s_1_2_2(mux_350_nl, or_1187_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign mux_352_nl = MUX_s_1_2_2(mux_tmp_342, mux_351_nl, while_stage_0_5);
  assign and_dcpl_626 = (~ mux_352_nl) & and_dcpl_529;
  assign mux_354_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_5_6_sva,
      while_mux_1285_tmp, while_stage_0_5);
  assign or_dcpl_677 = (mux_354_nl & (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]))
      | weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp;
  assign and_775_cse = (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5]) & weight_mem_read_arbxbar_arbiters_next_5_3_sva;
  assign and_776_cse = weight_mem_read_arbxbar_arbiters_next_5_4_sva & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5]);
  assign or_tmp_511 = and_775_cse | and_776_cse | weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_3_tmp;
  assign Arbiter_8U_Roundrobin_pick_1_mux_595_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_5_1_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_396_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign and_777_cse = (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[5]) & Arbiter_8U_Roundrobin_pick_1_mux_595_nl;
  assign and_778_cse = (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5]) & Arbiter_8U_Roundrobin_pick_1_mux_394_itm_1;
  assign and_779_cse = Arbiter_8U_Roundrobin_pick_1_mux_393_itm_1 & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5]);
  assign and_780_cse = (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[5]) & Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_41_mx1w0;
  assign or_1199_nl = and_778_cse | and_779_cse | weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_3_tmp;
  assign mux_356_nl = MUX_s_1_2_2(or_tmp_511, or_1199_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign or_1200_nl = and_777_cse | mux_356_nl;
  assign or_1194_nl = (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[5])
      | weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_3_tmp;
  assign mux_355_nl = MUX_s_1_2_2(or_tmp_511, or_1194_nl, weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[5]);
  assign or_1197_nl = and_780_cse | mux_355_nl;
  assign mux_tmp_353 = MUX_s_1_2_2(or_1200_nl, or_1197_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_781_cse = (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[5]) & weight_mem_read_arbxbar_arbiters_next_5_1_sva;
  assign or_tmp_517 = and_781_cse | or_tmp_511;
  assign mux_359_nl = MUX_s_1_2_2(or_tmp_517, mux_tmp_353, while_stage_0_5);
  assign nor_407_nl = ~(weight_mem_read_arbxbar_arbiters_next_5_6_sva | (~ or_tmp_517));
  assign nor_408_nl = ~(while_mux_1285_tmp | (~ mux_tmp_353));
  assign mux_358_nl = MUX_s_1_2_2(nor_407_nl, nor_408_nl, while_stage_0_5);
  assign mux_360_nl = MUX_s_1_2_2(mux_359_nl, mux_358_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]);
  assign and_dcpl_629 = mux_360_nl & (~(weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp));
  assign and_dcpl_631 = ~(weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_3_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_4_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_8_tmp);
  assign or_tmp_521 = and_775_cse | and_776_cse;
  assign or_1208_nl = and_778_cse | and_779_cse;
  assign mux_362_nl = MUX_s_1_2_2(or_tmp_521, or_1208_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign or_1209_nl = and_777_cse | mux_362_nl;
  assign mux_361_nl = MUX_s_1_2_2(or_tmp_521, operator_2_false_5_operator_2_false_5_or_mdf_6_sva_1,
      weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1[5]);
  assign or_1207_nl = and_780_cse | mux_361_nl;
  assign mux_tmp_359 = MUX_s_1_2_2(or_1209_nl, or_1207_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign or_tmp_526 = and_781_cse | or_tmp_521;
  assign or_1212_nl = weight_mem_read_arbxbar_arbiters_next_5_6_sva | or_tmp_526;
  assign or_1210_nl = while_mux_1285_tmp | mux_tmp_359;
  assign mux_tmp_360 = MUX_s_1_2_2(or_1212_nl, or_1210_nl, while_stage_0_5);
  assign mux_tmp_361 = MUX_s_1_2_2(or_tmp_526, mux_tmp_359, while_stage_0_5);
  assign mux_tmp_362 = MUX_s_1_2_2(mux_tmp_361, mux_tmp_360, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]);
  assign nand_3_nl = ~((weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]) & (~
      mux_tmp_360));
  assign or_1204_nl = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[5]);
  assign mux_367_nl = MUX_s_1_2_2(nand_3_nl, mux_tmp_362, or_1204_nl);
  assign and_dcpl_632 = (~ mux_367_nl) & and_dcpl_631;
  assign and_dcpl_639 = ~(mux_tmp_361 | weight_mem_read_arbxbar_xbar_1_for_3_6_Arbiter_8U_Roundrobin_pick_1_priority_and_3_tmp
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[5])
      | (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[5]) | (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[5]));
  assign and_789_cse = (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]) & while_mux_1278_tmp;
  assign and_790_cse = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4]) & while_mux_1279_tmp;
  assign or_tmp_528 = and_789_cse | and_790_cse;
  assign and_791_cse = (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]) & weight_mem_read_arbxbar_arbiters_next_4_6_sva;
  assign and_792_cse = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4]) & weight_mem_read_arbxbar_arbiters_next_4_5_sva;
  assign or_tmp_530 = and_791_cse | and_792_cse;
  assign mux_369_nl = MUX_s_1_2_2(or_tmp_530, or_tmp_528, while_stage_0_5);
  assign or_1216_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_itm_1
      | or_tmp_530;
  assign or_1214_nl = while_mux_1277_tmp | or_tmp_528;
  assign mux_368_nl = MUX_s_1_2_2(or_1216_nl, or_1214_nl, while_stage_0_5);
  assign mux_tmp_366 = MUX_s_1_2_2(mux_369_nl, mux_368_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4]);
  assign nor_tmp_123 = while_mux_1280_tmp & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4]);
  assign or_tmp_532 = ((weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4]) & while_mux_1281_tmp)
      | nor_tmp_123;
  assign or_tmp_533 = ((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[4]) & while_mux_1283_tmp)
      | or_tmp_532;
  assign or_tmp_534 = ((weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[4]) & while_mux_1282_tmp)
      | or_tmp_533;
  assign or_tmp_536 = and_789_cse | (~((~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4])
      & while_mux_1279_tmp)) & or_tmp_534));
  assign nor_tmp_129 = weight_mem_read_arbxbar_arbiters_next_4_4_sva & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4]);
  assign or_tmp_538 = ((weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4]) & weight_mem_read_arbxbar_arbiters_next_4_3_sva)
      | nor_tmp_129;
  assign or_tmp_539 = ((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[4]) & weight_mem_read_arbxbar_arbiters_next_4_1_sva)
      | or_tmp_538;
  assign or_tmp_540 = ((weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[4]) & weight_mem_read_arbxbar_arbiters_next_4_2_sva)
      | or_tmp_539;
  assign or_tmp_542 = and_791_cse | (~((~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4])
      & weight_mem_read_arbxbar_arbiters_next_4_5_sva)) & or_tmp_540));
  assign mux_372_nl = MUX_s_1_2_2(or_tmp_542, or_tmp_536, while_stage_0_5);
  assign or_1228_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_itm_1
      | or_tmp_542;
  assign or_1222_nl = while_mux_1277_tmp | or_tmp_536;
  assign mux_371_nl = MUX_s_1_2_2(or_1228_nl, or_1222_nl, while_stage_0_5);
  assign mux_373_itm = MUX_s_1_2_2(mux_372_nl, mux_371_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4]);
  assign or_tmp_544 = and_790_cse | or_tmp_534;
  assign or_tmp_545 = and_789_cse | or_tmp_544;
  assign or_tmp_547 = and_792_cse | or_tmp_540;
  assign or_tmp_548 = and_791_cse | or_tmp_547;
  assign or_1234_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_itm_1
      | or_tmp_548;
  assign or_1231_nl = while_mux_1277_tmp | or_tmp_545;
  assign mux_tmp_370 = MUX_s_1_2_2(or_1234_nl, or_1231_nl, while_stage_0_5);
  assign mux_tmp_371 = MUX_s_1_2_2(or_tmp_548, or_tmp_545, while_stage_0_5);
  assign or_1240_nl = (~ (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4])) |
      weight_mem_read_arbxbar_arbiters_next_4_5_sva | or_tmp_540;
  assign or_1238_nl = weight_mem_read_arbxbar_arbiters_next_4_6_sva | or_tmp_547;
  assign mux_377_nl = MUX_s_1_2_2(or_1240_nl, or_1238_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]);
  assign or_1237_nl = (~ (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[4])) |
      while_mux_1279_tmp | or_tmp_534;
  assign or_1235_nl = while_mux_1278_tmp | or_tmp_544;
  assign mux_376_nl = MUX_s_1_2_2(or_1237_nl, or_1235_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[4]);
  assign mux_378_nl = MUX_s_1_2_2(mux_377_nl, mux_376_nl, while_stage_0_5);
  assign mux_379_nl = MUX_s_1_2_2(mux_378_nl, mux_tmp_371, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[4]);
  assign mux_380_itm = MUX_s_1_2_2(mux_379_nl, mux_tmp_370, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[4]);
  assign nor_417_nl = ~(weight_mem_read_arbxbar_arbiters_next_4_4_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4])));
  assign nor_418_nl = ~(weight_mem_read_arbxbar_arbiters_next_4_3_sva | nor_tmp_129);
  assign mux_384_nl = MUX_s_1_2_2(nor_417_nl, nor_418_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4]);
  assign nor_419_nl = ~(weight_mem_read_arbxbar_arbiters_next_4_1_sva | or_tmp_538);
  assign mux_385_nl = MUX_s_1_2_2(mux_384_nl, nor_419_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[4]);
  assign nor_420_nl = ~(weight_mem_read_arbxbar_arbiters_next_4_2_sva | or_tmp_539);
  assign mux_386_nl = MUX_s_1_2_2(mux_385_nl, nor_420_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[4]);
  assign nor_421_nl = ~(while_mux_1280_tmp | (~ (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[4])));
  assign nor_422_nl = ~(while_mux_1281_tmp | nor_tmp_123);
  assign mux_381_nl = MUX_s_1_2_2(nor_421_nl, nor_422_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[4]);
  assign nor_423_nl = ~(while_mux_1283_tmp | or_tmp_532);
  assign mux_382_nl = MUX_s_1_2_2(mux_381_nl, nor_423_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[4]);
  assign nor_424_nl = ~(while_mux_1282_tmp | or_tmp_533);
  assign mux_383_nl = MUX_s_1_2_2(mux_382_nl, nor_424_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[4]);
  assign mux_387_nl = MUX_s_1_2_2(mux_386_nl, mux_383_nl, while_stage_0_5);
  assign and_dcpl_641 = mux_387_nl & and_dcpl_543;
  assign and_809_cse = (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]) & while_mux_1271_tmp;
  assign and_810_cse = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3]) & while_mux_1272_tmp;
  assign or_tmp_564 = and_809_cse | and_810_cse;
  assign and_811_cse = (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]) & weight_mem_read_arbxbar_arbiters_next_3_6_sva;
  assign and_812_cse = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3]) & weight_mem_read_arbxbar_arbiters_next_3_5_sva;
  assign or_tmp_566 = and_811_cse | and_812_cse;
  assign mux_390_nl = MUX_s_1_2_2(or_tmp_566, or_tmp_564, while_stage_0_5);
  assign or_1252_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_itm_1
      | or_tmp_566;
  assign or_1250_nl = while_mux_1270_tmp | or_tmp_564;
  assign mux_389_nl = MUX_s_1_2_2(or_1252_nl, or_1250_nl, while_stage_0_5);
  assign mux_tmp_387 = MUX_s_1_2_2(mux_390_nl, mux_389_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3]);
  assign nor_tmp_143 = while_mux_1274_tmp & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3]);
  assign or_tmp_568 = ((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[3]) & while_mux_1276_tmp)
      | nor_tmp_143;
  assign or_tmp_569 = ((weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[3]) & while_mux_1275_tmp)
      | or_tmp_568;
  assign or_tmp_570 = ((weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[3]) & while_mux_1273_tmp)
      | or_tmp_569;
  assign or_tmp_572 = and_809_cse | (~((~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3])
      & while_mux_1272_tmp)) & or_tmp_570));
  assign nor_tmp_149 = weight_mem_read_arbxbar_arbiters_next_3_3_sva & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3]);
  assign or_tmp_574 = ((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[3]) & weight_mem_read_arbxbar_arbiters_next_3_1_sva)
      | nor_tmp_149;
  assign or_tmp_575 = ((weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[3]) & weight_mem_read_arbxbar_arbiters_next_3_2_sva)
      | or_tmp_574;
  assign or_tmp_576 = ((weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[3]) & weight_mem_read_arbxbar_arbiters_next_3_4_sva)
      | or_tmp_575;
  assign or_tmp_578 = and_811_cse | (~((~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3])
      & weight_mem_read_arbxbar_arbiters_next_3_5_sva)) & or_tmp_576));
  assign mux_393_nl = MUX_s_1_2_2(or_tmp_578, or_tmp_572, while_stage_0_5);
  assign or_1264_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_itm_1
      | or_tmp_578;
  assign or_1258_nl = while_mux_1270_tmp | or_tmp_572;
  assign mux_392_nl = MUX_s_1_2_2(or_1264_nl, or_1258_nl, while_stage_0_5);
  assign mux_394_itm = MUX_s_1_2_2(mux_393_nl, mux_392_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3]);
  assign or_tmp_580 = and_810_cse | or_tmp_570;
  assign or_tmp_581 = and_809_cse | or_tmp_580;
  assign or_tmp_583 = and_812_cse | or_tmp_576;
  assign or_tmp_584 = and_811_cse | or_tmp_583;
  assign or_1270_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_itm_1
      | or_tmp_584;
  assign or_1267_nl = while_mux_1270_tmp | or_tmp_581;
  assign mux_tmp_391 = MUX_s_1_2_2(or_1270_nl, or_1267_nl, while_stage_0_5);
  assign mux_tmp_392 = MUX_s_1_2_2(or_tmp_584, or_tmp_581, while_stage_0_5);
  assign or_1276_nl = (~ (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3])) |
      weight_mem_read_arbxbar_arbiters_next_3_5_sva | or_tmp_576;
  assign or_1274_nl = weight_mem_read_arbxbar_arbiters_next_3_6_sva | or_tmp_583;
  assign mux_398_nl = MUX_s_1_2_2(or_1276_nl, or_1274_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]);
  assign or_1273_nl = (~ (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[3])) |
      while_mux_1272_tmp | or_tmp_570;
  assign or_1271_nl = while_mux_1271_tmp | or_tmp_580;
  assign mux_397_nl = MUX_s_1_2_2(or_1273_nl, or_1271_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[3]);
  assign mux_399_nl = MUX_s_1_2_2(mux_398_nl, mux_397_nl, while_stage_0_5);
  assign mux_400_nl = MUX_s_1_2_2(mux_399_nl, mux_tmp_392, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[3]);
  assign mux_401_itm = MUX_s_1_2_2(mux_400_nl, mux_tmp_391, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[3]);
  assign nor_425_nl = ~(weight_mem_read_arbxbar_arbiters_next_3_3_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3])));
  assign nor_426_nl = ~(weight_mem_read_arbxbar_arbiters_next_3_1_sva | nor_tmp_149);
  assign mux_405_nl = MUX_s_1_2_2(nor_425_nl, nor_426_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[3]);
  assign nor_427_nl = ~(weight_mem_read_arbxbar_arbiters_next_3_2_sva | or_tmp_574);
  assign mux_406_nl = MUX_s_1_2_2(mux_405_nl, nor_427_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[3]);
  assign nor_428_nl = ~(weight_mem_read_arbxbar_arbiters_next_3_4_sva | or_tmp_575);
  assign mux_407_nl = MUX_s_1_2_2(mux_406_nl, nor_428_nl, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[3]);
  assign nor_429_nl = ~(while_mux_1274_tmp | (~ (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[3])));
  assign nor_430_nl = ~(while_mux_1276_tmp | nor_tmp_143);
  assign mux_402_nl = MUX_s_1_2_2(nor_429_nl, nor_430_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[3]);
  assign nor_431_nl = ~(while_mux_1275_tmp | or_tmp_568);
  assign mux_403_nl = MUX_s_1_2_2(mux_402_nl, nor_431_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[3]);
  assign nor_432_nl = ~(while_mux_1273_tmp | or_tmp_569);
  assign mux_404_nl = MUX_s_1_2_2(mux_403_nl, nor_432_nl, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[3]);
  assign mux_408_nl = MUX_s_1_2_2(mux_407_nl, mux_404_nl, while_stage_0_5);
  assign and_dcpl_642 = mux_408_nl & and_dcpl_550;
  assign and_829_cse = (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]) & while_mux_1264_tmp;
  assign and_830_cse = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2]) & while_mux_1265_tmp;
  assign or_tmp_600 = and_829_cse | and_830_cse;
  assign and_831_cse = (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]) & weight_mem_read_arbxbar_arbiters_next_2_6_sva;
  assign and_832_cse = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2]) & weight_mem_read_arbxbar_arbiters_next_2_5_sva;
  assign or_tmp_602 = and_831_cse | and_832_cse;
  assign mux_411_nl = MUX_s_1_2_2(or_tmp_602, or_tmp_600, while_stage_0_5);
  assign or_1288_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_itm_1
      | or_tmp_602;
  assign or_1286_nl = while_mux_1263_tmp | or_tmp_600;
  assign mux_410_nl = MUX_s_1_2_2(or_1288_nl, or_1286_nl, while_stage_0_5);
  assign mux_tmp_408 = MUX_s_1_2_2(mux_411_nl, mux_410_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2]);
  assign nor_tmp_163 = while_mux_1267_tmp & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2]);
  assign or_tmp_604 = ((weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]) & while_mux_1268_tmp)
      | nor_tmp_163;
  assign or_tmp_605 = ((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[2]) & while_mux_1269_tmp)
      | or_tmp_604;
  assign or_tmp_606 = ((weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2]) & while_mux_1266_tmp)
      | or_tmp_605;
  assign or_tmp_608 = and_829_cse | (~((~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2])
      & while_mux_1265_tmp)) & or_tmp_606));
  assign nor_tmp_169 = weight_mem_read_arbxbar_arbiters_next_2_3_sva & (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2]);
  assign or_tmp_610 = ((weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]) & weight_mem_read_arbxbar_arbiters_next_2_2_sva)
      | nor_tmp_169;
  assign or_tmp_611 = ((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[2]) & weight_mem_read_arbxbar_arbiters_next_2_1_sva)
      | or_tmp_610;
  assign or_tmp_612 = ((weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2]) & weight_mem_read_arbxbar_arbiters_next_2_4_sva)
      | or_tmp_611;
  assign or_tmp_614 = and_831_cse | (~((~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2])
      & weight_mem_read_arbxbar_arbiters_next_2_5_sva)) & or_tmp_612));
  assign mux_414_nl = MUX_s_1_2_2(or_tmp_614, or_tmp_608, while_stage_0_5);
  assign or_1300_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_itm_1
      | or_tmp_614;
  assign or_1294_nl = while_mux_1263_tmp | or_tmp_608;
  assign mux_413_nl = MUX_s_1_2_2(or_1300_nl, or_1294_nl, while_stage_0_5);
  assign mux_415_itm = MUX_s_1_2_2(mux_414_nl, mux_413_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2]);
  assign or_tmp_616 = and_830_cse | or_tmp_606;
  assign or_tmp_617 = and_829_cse | or_tmp_616;
  assign or_tmp_619 = and_832_cse | or_tmp_612;
  assign or_tmp_620 = and_831_cse | or_tmp_619;
  assign or_1306_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_itm_1
      | or_tmp_620;
  assign or_1303_nl = while_mux_1263_tmp | or_tmp_617;
  assign mux_tmp_412 = MUX_s_1_2_2(or_1306_nl, or_1303_nl, while_stage_0_5);
  assign mux_tmp_413 = MUX_s_1_2_2(or_tmp_620, or_tmp_617, while_stage_0_5);
  assign or_1312_nl = (~ (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2])) |
      weight_mem_read_arbxbar_arbiters_next_2_5_sva | or_tmp_612;
  assign or_1310_nl = weight_mem_read_arbxbar_arbiters_next_2_6_sva | or_tmp_619;
  assign mux_419_nl = MUX_s_1_2_2(or_1312_nl, or_1310_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]);
  assign or_1309_nl = (~ (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[2])) |
      while_mux_1265_tmp | or_tmp_606;
  assign or_1307_nl = while_mux_1264_tmp | or_tmp_616;
  assign mux_418_nl = MUX_s_1_2_2(or_1309_nl, or_1307_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[2]);
  assign mux_420_nl = MUX_s_1_2_2(mux_419_nl, mux_418_nl, while_stage_0_5);
  assign mux_421_nl = MUX_s_1_2_2(mux_420_nl, mux_tmp_413, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[2]);
  assign mux_422_itm = MUX_s_1_2_2(mux_421_nl, mux_tmp_412, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[2]);
  assign nor_433_nl = ~(weight_mem_read_arbxbar_arbiters_next_2_3_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2])));
  assign nor_434_nl = ~(weight_mem_read_arbxbar_arbiters_next_2_2_sva | nor_tmp_169);
  assign mux_426_nl = MUX_s_1_2_2(nor_433_nl, nor_434_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]);
  assign nor_435_nl = ~(weight_mem_read_arbxbar_arbiters_next_2_1_sva | or_tmp_610);
  assign mux_427_nl = MUX_s_1_2_2(mux_426_nl, nor_435_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[2]);
  assign nor_436_nl = ~(weight_mem_read_arbxbar_arbiters_next_2_4_sva | or_tmp_611);
  assign mux_428_nl = MUX_s_1_2_2(mux_427_nl, nor_436_nl, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2]);
  assign nor_437_nl = ~(while_mux_1267_tmp | (~ (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[2])));
  assign nor_438_nl = ~(while_mux_1268_tmp | nor_tmp_163);
  assign mux_423_nl = MUX_s_1_2_2(nor_437_nl, nor_438_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[2]);
  assign nor_439_nl = ~(while_mux_1269_tmp | or_tmp_604);
  assign mux_424_nl = MUX_s_1_2_2(mux_423_nl, nor_439_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[2]);
  assign nor_440_nl = ~(while_mux_1266_tmp | or_tmp_605);
  assign mux_425_nl = MUX_s_1_2_2(mux_424_nl, nor_440_nl, weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[2]);
  assign mux_429_nl = MUX_s_1_2_2(mux_428_nl, mux_425_nl, while_stage_0_5);
  assign and_dcpl_643 = mux_429_nl & and_dcpl_557;
  assign and_849_cse = (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]) & while_mux_1257_tmp;
  assign and_850_cse = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1]) & while_mux_1258_tmp;
  assign or_tmp_636 = and_849_cse | and_850_cse;
  assign and_851_cse = (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]) & weight_mem_read_arbxbar_arbiters_next_1_6_sva;
  assign and_852_cse = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1]) & weight_mem_read_arbxbar_arbiters_next_1_5_sva;
  assign or_tmp_638 = and_851_cse | and_852_cse;
  assign mux_432_nl = MUX_s_1_2_2(or_tmp_638, or_tmp_636, while_stage_0_5);
  assign or_1324_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1
      | or_tmp_638;
  assign or_1322_nl = while_mux_1256_tmp | or_tmp_636;
  assign mux_431_nl = MUX_s_1_2_2(or_1324_nl, or_1322_nl, while_stage_0_5);
  assign mux_tmp_429 = MUX_s_1_2_2(mux_432_nl, mux_431_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1]);
  assign and_855_cse = while_mux_1259_tmp & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]);
  assign and_853_cse = (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]) & while_mux_1261_tmp;
  assign or_1325_nl = and_855_cse | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1]);
  assign mux_434_nl = MUX_s_1_2_2(and_855_cse, or_1325_nl, while_mux_1260_tmp);
  assign or_tmp_642 = and_853_cse | ((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1])
      & while_mux_1262_tmp) | mux_434_nl;
  assign or_tmp_644 = and_849_cse | (~((~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1])
      & while_mux_1258_tmp)) & or_tmp_642));
  assign and_861_cse = weight_mem_read_arbxbar_arbiters_next_1_4_sva & (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1]);
  assign and_859_cse = (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]) & weight_mem_read_arbxbar_arbiters_next_1_2_sva;
  assign or_1331_nl = and_861_cse | (weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1]);
  assign mux_435_nl = MUX_s_1_2_2(and_861_cse, or_1331_nl, weight_mem_read_arbxbar_arbiters_next_1_3_sva);
  assign or_tmp_648 = and_859_cse | ((weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1])
      & weight_mem_read_arbxbar_arbiters_next_1_1_sva) | mux_435_nl;
  assign or_tmp_650 = and_851_cse | (~((~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1])
      & weight_mem_read_arbxbar_arbiters_next_1_5_sva)) & or_tmp_648));
  assign mux_437_nl = MUX_s_1_2_2(or_tmp_650, or_tmp_644, while_stage_0_5);
  assign or_1336_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1
      | or_tmp_650;
  assign or_1330_nl = while_mux_1256_tmp | or_tmp_644;
  assign mux_436_nl = MUX_s_1_2_2(or_1336_nl, or_1330_nl, while_stage_0_5);
  assign mux_438_itm = MUX_s_1_2_2(mux_437_nl, mux_436_nl, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1]);
  assign or_tmp_652 = and_850_cse | or_tmp_642;
  assign or_tmp_653 = and_849_cse | or_tmp_652;
  assign or_tmp_655 = and_852_cse | or_tmp_648;
  assign or_tmp_656 = and_851_cse | or_tmp_655;
  assign or_1342_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1
      | or_tmp_656;
  assign or_1339_nl = while_mux_1256_tmp | or_tmp_653;
  assign mux_tmp_435 = MUX_s_1_2_2(or_1342_nl, or_1339_nl, while_stage_0_5);
  assign mux_tmp_436 = MUX_s_1_2_2(or_tmp_656, or_tmp_653, while_stage_0_5);
  assign or_1348_nl = (~ (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1])) |
      weight_mem_read_arbxbar_arbiters_next_1_5_sva | or_tmp_648;
  assign or_1346_nl = weight_mem_read_arbxbar_arbiters_next_1_6_sva | or_tmp_655;
  assign mux_442_nl = MUX_s_1_2_2(or_1348_nl, or_1346_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]);
  assign or_1345_nl = (~ (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[1])) |
      while_mux_1258_tmp | or_tmp_642;
  assign or_1343_nl = while_mux_1257_tmp | or_tmp_652;
  assign mux_441_nl = MUX_s_1_2_2(or_1345_nl, or_1343_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[1]);
  assign mux_443_nl = MUX_s_1_2_2(mux_442_nl, mux_441_nl, while_stage_0_5);
  assign mux_444_nl = MUX_s_1_2_2(mux_443_nl, mux_tmp_436, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[1]);
  assign mux_445_itm = MUX_s_1_2_2(mux_444_nl, mux_tmp_435, weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[1]);
  assign or_tmp_665 = and_853_cse | and_855_cse;
  assign or_tmp_668 = and_859_cse | and_861_cse;
  assign nor_441_nl = ~(weight_mem_read_arbxbar_arbiters_next_1_4_sva | (~ (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1])));
  assign nor_442_nl = ~(weight_mem_read_arbxbar_arbiters_next_1_2_sva | and_861_cse);
  assign mux_451_nl = MUX_s_1_2_2(nor_441_nl, nor_442_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]);
  assign nor_443_nl = ~(while_mux_1259_tmp | (~ (weight_mem_read_arbxbar_xbar_1_for_5_lshift_tmp[1])));
  assign nor_444_nl = ~(while_mux_1261_tmp | and_855_cse);
  assign mux_450_nl = MUX_s_1_2_2(nor_443_nl, nor_444_nl, weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[1]);
  assign mux_452_nl = MUX_s_1_2_2(mux_451_nl, mux_450_nl, while_stage_0_5);
  assign nor_445_nl = ~(weight_mem_read_arbxbar_arbiters_next_1_3_sva | or_tmp_668);
  assign nor_446_nl = ~(while_mux_1260_tmp | or_tmp_665);
  assign mux_449_nl = MUX_s_1_2_2(nor_445_nl, nor_446_nl, while_stage_0_5);
  assign mux_453_nl = MUX_s_1_2_2(mux_452_nl, mux_449_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1]);
  assign nor_447_nl = ~(weight_mem_read_arbxbar_arbiters_next_1_1_sva | or_tmp_668);
  assign nor_448_nl = ~(while_mux_1262_tmp | or_tmp_665);
  assign mux_447_nl = MUX_s_1_2_2(nor_447_nl, nor_448_nl, while_stage_0_5);
  assign nor_449_nl = ~(weight_mem_read_arbxbar_arbiters_next_1_1_sva | weight_mem_read_arbxbar_arbiters_next_1_3_sva
      | or_tmp_668);
  assign nor_450_nl = ~(while_mux_1260_tmp | while_mux_1262_tmp | or_tmp_665);
  assign mux_446_nl = MUX_s_1_2_2(nor_449_nl, nor_450_nl, while_stage_0_5);
  assign mux_448_nl = MUX_s_1_2_2(mux_447_nl, mux_446_nl, weight_mem_read_arbxbar_xbar_1_for_4_lshift_tmp[1]);
  assign mux_454_nl = MUX_s_1_2_2(mux_453_nl, mux_448_nl, weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[1]);
  assign and_dcpl_644 = mux_454_nl & and_dcpl_564;
  assign and_873_cse = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0]) & while_mux_1251_tmp;
  assign and_874_cse = while_mux_1249_tmp & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0]);
  assign or_tmp_678 = and_873_cse | and_874_cse;
  assign and_875_cse = (weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0]) & weight_mem_read_arbxbar_arbiters_next_0_5_sva;
  assign and_876_cse = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1
      & (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0]);
  assign or_tmp_680 = and_875_cse | and_876_cse;
  assign mux_457_nl = MUX_s_1_2_2(or_tmp_680, or_tmp_678, while_stage_0_5);
  assign or_1366_nl = weight_mem_read_arbxbar_arbiters_next_0_6_sva | or_tmp_680;
  assign or_1364_nl = while_mux_1250_tmp | or_tmp_678;
  assign mux_456_nl = MUX_s_1_2_2(or_1366_nl, or_1364_nl, while_stage_0_5);
  assign mux_tmp_454 = MUX_s_1_2_2(mux_457_nl, mux_456_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]);
  assign Arbiter_8U_Roundrobin_pick_1_mux_626_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_0_2_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_30_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1);
  assign while_mux_1254_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_626_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_5_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_879_cse = (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0]) & while_mux_1254_nl;
  assign Arbiter_8U_Roundrobin_pick_1_mux_625_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_arbiters_next_0_1_sva,
      Arbiter_8U_Roundrobin_pick_1_mux_31_itm_1, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1);
  assign while_mux_1255_nl = MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_mux_625_nl,
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_6_mx1w0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_880_cse = while_mux_1255_nl & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[0]);
  assign or_tmp_685 = and_873_cse | and_874_cse | (~(and_879_cse | and_880_cse |
      weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_1_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp));
  assign and_883_cse = (weight_mem_read_arbxbar_xbar_1_for_3_lshift_tmp[0]) & weight_mem_read_arbxbar_arbiters_next_0_2_sva;
  assign and_884_cse = weight_mem_read_arbxbar_arbiters_next_0_1_sva & (weight_mem_read_arbxbar_xbar_1_for_2_lshift_tmp[0]);
  assign or_tmp_690 = and_875_cse | and_876_cse | (~(and_883_cse | and_884_cse |
      weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_1_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp));
  assign mux_460_nl = MUX_s_1_2_2(or_tmp_690, or_tmp_685, while_stage_0_5);
  assign or_1376_nl = weight_mem_read_arbxbar_arbiters_next_0_6_sva | or_tmp_690;
  assign or_1371_nl = while_mux_1250_tmp | or_tmp_685;
  assign mux_459_nl = MUX_s_1_2_2(or_1376_nl, or_1371_nl, while_stage_0_5);
  assign mux_461_itm = MUX_s_1_2_2(mux_460_nl, mux_459_nl, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]);
  assign and_dcpl_645 = ~(weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_2_tmp
      | weight_mem_read_arbxbar_xbar_1_for_3_1_Arbiter_8U_Roundrobin_pick_1_priority_and_1_tmp);
  assign or_tmp_692 = and_879_cse | and_880_cse;
  assign or_tmp_693 = and_874_cse | or_tmp_692;
  assign or_tmp_694 = and_873_cse | or_tmp_693;
  assign or_tmp_696 = and_883_cse | and_884_cse;
  assign or_tmp_697 = and_876_cse | or_tmp_696;
  assign or_tmp_698 = and_875_cse | or_tmp_697;
  assign or_1384_nl = weight_mem_read_arbxbar_arbiters_next_0_6_sva | or_tmp_698;
  assign or_1380_nl = while_mux_1250_tmp | or_tmp_694;
  assign mux_tmp_458 = MUX_s_1_2_2(or_1384_nl, or_1380_nl, while_stage_0_5);
  assign mux_tmp_459 = MUX_s_1_2_2(or_tmp_698, or_tmp_694, while_stage_0_5);
  assign or_1397_nl = Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1
      | (~ (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0])) | or_tmp_696;
  assign or_1386_nl = weight_mem_read_arbxbar_arbiters_next_0_5_sva | or_tmp_697;
  assign mux_465_nl = MUX_s_1_2_2(or_1397_nl, or_1386_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0]);
  assign or_1398_nl = while_mux_1249_tmp | (~ (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0]))
      | or_tmp_692;
  assign or_1385_nl = while_mux_1251_tmp | or_tmp_693;
  assign mux_464_nl = MUX_s_1_2_2(or_1398_nl, or_1385_nl, weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0]);
  assign mux_466_nl = MUX_s_1_2_2(mux_465_nl, mux_464_nl, while_stage_0_5);
  assign mux_467_nl = MUX_s_1_2_2(mux_466_nl, mux_tmp_459, weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0]);
  assign mux_468_nl = MUX_s_1_2_2(mux_467_nl, mux_tmp_458, weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0]);
  assign and_dcpl_646 = (~ mux_468_nl) & and_dcpl_645;
  assign mux_469_nl = MUX_s_1_2_2(or_tmp_696, or_tmp_692, while_stage_0_5);
  assign and_dcpl_651 = (~ mux_469_nl) & and_dcpl_645 & (~ (weight_mem_read_arbxbar_xbar_1_for_8_lshift_tmp[0]))
      & (~((weight_mem_read_arbxbar_xbar_1_for_6_lshift_tmp[0]) | (weight_mem_read_arbxbar_xbar_1_for_1_lshift_tmp[0])
      | (weight_mem_read_arbxbar_xbar_1_for_7_lshift_tmp[0])));
  assign or_dcpl_678 = ~(Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1 & weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs);
  assign PECore_PushAxiRsp_mux_13_itm_1_mx0c1 = and_dcpl_241 & (~ rva_in_reg_rw_sva_5);
  assign ProductSum_for_acc_11_cmp_a = weight_port_read_out_data_7_1_sva_dfm_2;
  assign ProductSum_for_acc_11_cmp_b_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[15:8];
  assign ProductSum_for_acc_11_cmp_load_pff = ProductSum_for_asn_16_itm_5;
  assign ProductSum_for_acc_11_cmp_datavalid_pff = and_dcpl_31;
  assign ProductSum_for_acc_10_cmp_a = weight_port_read_out_data_7_0_sva_dfm_2;
  assign ProductSum_for_acc_10_cmp_b_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[7:0];
  assign ProductSum_for_acc_9_cmp_a0 = weight_port_read_out_data_7_5_sva_dfm_1;
  assign ProductSum_for_acc_9_cmp_a1_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5_63_16[31:24];
  assign ProductSum_for_acc_9_cmp_b0 = weight_port_read_out_data_7_2_sva_dfm_1;
  assign ProductSum_for_acc_9_cmp_b1_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5_63_16[7:0];
  assign ProductSum_for_acc_9_cmp_c0 = weight_port_read_out_data_7_3_sva_dfm_1;
  assign ProductSum_for_acc_9_cmp_c1_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5_63_16[15:8];
  assign ProductSum_for_acc_9_cmp_load_pff = ProductSum_for_asn_12_itm_6;
  assign ProductSum_for_acc_9_cmp_datavalid_pff = and_dcpl_459;
  assign ProductSum_for_acc_8_cmp_a0 = weight_port_read_out_data_7_6_sva_dfm_1;
  assign ProductSum_for_acc_8_cmp_a1_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5_63_16[39:32];
  assign ProductSum_for_acc_8_cmp_b0 = weight_port_read_out_data_7_7_sva_dfm_1;
  assign ProductSum_for_acc_8_cmp_b1_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5_63_16[47:40];
  assign ProductSum_for_acc_8_cmp_c0 = weight_port_read_out_data_7_4_sva_dfm_1;
  assign ProductSum_for_acc_8_cmp_c1_pff = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5_63_16[23:16];
  assign PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_a = MUX_v_8_2_2(weight_port_read_out_data_6_1_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_2_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2,
      weight_mem_run_3_for_land_7_lpi_1_dfm_2);
  assign PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_load_pff = ProductSum_for_asn_25_itm_5;
  assign PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_4_cmp_a = MUX_v_8_2_2(weight_port_read_out_data_6_0_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_1_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2,
      weight_mem_run_3_for_land_7_lpi_1_dfm_2);
  assign PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_a0 = weight_mem_run_3_for_5_mux_53_itm_1;
  assign PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_b0 = weight_mem_run_3_for_5_mux_50_itm_1;
  assign PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_c0 = weight_mem_run_3_for_5_mux_51_itm_1;
  assign PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_load_pff = ProductSum_for_asn_23_itm_6;
  assign PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_a0 = weight_mem_run_3_for_5_mux_54_itm_1;
  assign PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_b0 = weight_mem_run_3_for_5_mux_55_itm_1;
  assign PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_c0 = weight_mem_run_3_for_5_mux_52_itm_1;
  assign PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_a = weight_port_read_out_data_5_1_sva_dfm_2;
  assign PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_load_pff = ProductSum_for_asn_42_itm_5;
  assign PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_4_cmp_a = weight_port_read_out_data_5_0_sva_dfm_2;
  assign PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_a0 = weight_port_read_out_data_5_5_sva_dfm_1;
  assign PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_b0 = weight_port_read_out_data_5_2_sva_dfm_1;
  assign PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_c0 = weight_port_read_out_data_5_3_sva_dfm_1;
  assign PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_load_pff = ProductSum_for_asn_38_itm_6;
  assign PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_a0 = weight_port_read_out_data_5_6_sva_dfm_1;
  assign PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_b0 = weight_port_read_out_data_5_7_sva_dfm_1;
  assign PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_c0 = weight_port_read_out_data_5_4_sva_dfm_1;
  assign PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_a = MUX_v_8_2_2(weight_port_read_out_data_4_1_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_2_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2,
      weight_mem_run_3_for_land_5_lpi_1_dfm_2);
  assign PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_load_pff = ProductSum_for_asn_51_itm_5;
  assign PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_4_cmp_a = MUX_v_8_2_2(weight_port_read_out_data_4_0_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_1_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2,
      weight_mem_run_3_for_land_5_lpi_1_dfm_2);
  assign PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_a0 = weight_mem_run_3_for_5_mux_37_itm_1;
  assign PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_b0 = weight_mem_run_3_for_5_mux_34_itm_1;
  assign PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_c0 = weight_mem_run_3_for_5_mux_35_itm_1;
  assign PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_load_pff = ProductSum_for_asn_49_itm_6;
  assign PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_a0 = weight_mem_run_3_for_5_mux_38_itm_1;
  assign PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_b0 = weight_mem_run_3_for_5_mux_39_itm_1;
  assign PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_c0 = weight_mem_run_3_for_5_mux_36_itm_1;
  assign PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_a = MUX_v_8_2_2(weight_port_read_out_data_3_1_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000000,
      weight_mem_run_3_for_land_4_lpi_1_dfm_2);
  assign PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_load_pff = ProductSum_for_asn_64_itm_5;
  assign PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_4_cmp_a = MUX_v_8_2_2(weight_port_read_out_data_3_0_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000001,
      weight_mem_run_3_for_land_4_lpi_1_dfm_2);
  assign PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_a0 = weight_port_read_out_data_3_5_sva_dfm_1;
  assign PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_b0 = weight_mem_run_3_for_5_mux_26_itm_1;
  assign PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_c0 = weight_mem_run_3_for_5_mux_27_itm_1;
  assign PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_load_pff = ProductSum_for_asn_62_itm_6;
  assign PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_a0 = weight_port_read_out_data_3_6_sva_dfm_1;
  assign PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_b0 = weight_port_read_out_data_3_7_sva_dfm_1;
  assign PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_c0 = weight_port_read_out_data_3_4_sva_dfm_1;
  assign PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_a = MUX_v_8_2_2(weight_port_read_out_data_2_1_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000000,
      weight_mem_run_3_for_land_3_lpi_1_dfm_2);
  assign PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_load = ProductSum_for_asn_73_itm_5;
  assign and_521_nl = fsm_output & (~ weight_mem_run_3_for_land_3_lpi_1_dfm_3);
  assign PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_a = MUX_v_8_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000001,
      weight_port_read_out_data_2_0_sva_dfm_1, and_521_nl);
  assign PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_b = input_mem_banks_read_1_read_data_lpi_1_dfm_1_5_7_0;
  assign PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_load_pff = ProductSum_for_asn_72_itm_6;
  assign PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_a0 = weight_mem_run_3_for_5_mux_21_itm_1;
  assign PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_b0 = weight_mem_run_3_for_5_mux_18_itm_1;
  assign PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_c0 = weight_mem_run_3_for_5_mux_19_itm_1;
  assign PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_a0 = weight_mem_run_3_for_5_mux_22_itm_1;
  assign PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_b0 = weight_mem_run_3_for_5_mux_23_itm_1;
  assign PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_c0 = weight_mem_run_3_for_5_mux_20_itm_1;
  assign PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_a = MUX_v_8_2_2(weight_port_read_out_data_1_1_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000000,
      weight_mem_run_3_for_land_2_lpi_1_dfm_2);
  assign PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_load_pff = ProductSum_for_asn_82_itm_5;
  assign PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_4_cmp_a = MUX_v_8_2_2(weight_port_read_out_data_1_0_sva_dfm_1,
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000001,
      weight_mem_run_3_for_land_2_lpi_1_dfm_2);
  assign PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_a0 = weight_mem_run_3_for_5_mux_13_itm_1;
  assign PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_b0 = {weight_mem_run_3_for_5_mux_10_itm_1_7
      , weight_mem_run_3_for_5_mux_10_itm_1_6_0};
  assign PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_c0 = {weight_mem_run_3_for_5_mux_11_itm_1_7
      , weight_mem_run_3_for_5_mux_11_itm_1_6_0};
  assign PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_load_pff = ProductSum_for_asn_80_itm_6;
  assign PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_a0 = weight_mem_run_3_for_5_mux_14_itm_1;
  assign PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_b0 = weight_mem_run_3_for_5_mux_15_itm_1;
  assign PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_c0 = {weight_mem_run_3_for_5_mux_12_itm_1_7_6
      , weight_mem_run_3_for_5_mux_12_itm_1_5_0};
  assign weight_port_read_out_data_mux_8_nl = MUX_s_1_2_2(weight_port_read_out_data_0_1_sva_dfm_2_7,
      PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_a_mx1_7, fsm_output);
  assign weight_port_read_out_data_mux_22_nl = MUX_v_7_2_2(weight_port_read_out_data_0_1_sva_dfm_2_6_0,
      PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_a_mx1_6_0, fsm_output);
  assign PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_a = {weight_port_read_out_data_mux_8_nl
      , weight_port_read_out_data_mux_22_nl};
  assign PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_load_pff = ProductSum_for_asn_98_itm_5;
  assign PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_a = {weight_port_read_out_data_0_0_sva_dfm_3_7
      , weight_port_read_out_data_0_0_sva_dfm_3_6_0};
  assign PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_a0 = {weight_port_read_out_data_0_3_sva_dfm_1_7
      , weight_port_read_out_data_0_3_sva_dfm_1_6_4 , weight_port_read_out_data_0_3_sva_dfm_1_3_0};
  assign PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_b0 = {weight_port_read_out_data_0_0_sva_dfm_1_7
      , weight_port_read_out_data_0_0_sva_dfm_1_6 , weight_port_read_out_data_0_0_sva_dfm_1_5_0};
  assign PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_c0 = {weight_port_read_out_data_0_1_sva_dfm_1_7
      , weight_port_read_out_data_0_1_sva_dfm_1_6_4 , weight_port_read_out_data_0_1_sva_dfm_1_3_0};
  assign PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_load_pff = ProductSum_for_asn_94_itm_6;
  assign PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_a0 = {weight_mem_run_3_for_5_mux_6_itm_1_7_4
      , weight_mem_run_3_for_5_mux_6_itm_1_3_0};
  assign PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_b0 = {weight_port_read_out_data_0_7_sva_dfm_1_1_rsp_0
      , weight_port_read_out_data_0_7_sva_dfm_1_1_rsp_1};
  assign PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_c0 = {weight_port_read_out_data_0_2_sva_dfm_1_7
      , weight_port_read_out_data_0_2_sva_dfm_1_6 , weight_port_read_out_data_0_2_sva_dfm_1_5_0};
  assign weight_mem_banks_bank_a0_a0_a0_a_rsci_d_d = {weight_write_data_data_0_7_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_6_lpi_1_dfm_1_2_6 , weight_write_data_data_0_5_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_4_lpi_1_dfm_1_2_6 , weight_write_data_data_0_3_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_2_lpi_1_dfm_1_2_6 , weight_write_data_data_0_1_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_0_lpi_1_dfm_1_2_6};
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_5_nl
      = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1
      | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0));
  assign weight_mem_banks_write_if_for_if_and_35_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_36_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_37_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_38_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_39_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_40_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_41_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1 & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_5_nl
      = MUX1HOT_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
      {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_5_nl
      , weight_mem_banks_write_if_for_if_and_35_nl , weight_mem_banks_write_if_for_if_and_36_nl
      , weight_mem_banks_write_if_for_if_and_37_nl , weight_mem_banks_write_if_for_if_and_38_nl
      , weight_mem_banks_write_if_for_if_and_39_nl , weight_mem_banks_write_if_for_if_and_40_nl
      , weight_mem_banks_write_if_for_if_and_41_nl});
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_nl = MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3,
      (weight_read_addrs_1_lpi_1_dfm_1[3]), (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_3_lpi_1_dfm_1[3]), (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]),
      (weight_read_addrs_5_lpi_1_dfm_1[3]), (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_7_lpi_1_dfm_1[3]), {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_2
      , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_1 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_18_0});
  assign weight_mem_banks_write_if_for_if_mux_7_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_nl,
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a0_a0_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_5_nl
      , weight_mem_banks_write_if_for_if_mux_7_nl};
  assign nor_463_nl = ~((~ PECore_PushOutput_PECore_PushOutput_if_and_svs_st_3) |
      PECore_RunFSM_switch_lp_equal_tmp_1_2);
  assign mux_256_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp,
      nor_463_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_pff = mux_256_nl & while_stage_0_5;
  assign weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_pff = weight_write_addrs_lpi_1_dfm_1_2[14:3];
  assign weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_pff = and_dcpl_178;
  assign weight_mem_banks_bank_a0_a0_a1_a_rsci_d_d = {weight_write_data_data_0_7_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_6_lpi_1_dfm_1_2_6 , weight_write_data_data_0_5_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_4_lpi_1_dfm_1_2_6 , weight_write_data_data_0_3_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_2_lpi_1_dfm_1_2_6 , weight_write_data_data_0_1_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_0_lpi_1_dfm_1_2_6};
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_4_nl
      = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1
      | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0));
  assign weight_mem_banks_write_if_for_if_and_28_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_29_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_30_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_31_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_32_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_33_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_34_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1 & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_4_nl
      = MUX1HOT_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
      {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_4_nl
      , weight_mem_banks_write_if_for_if_and_28_nl , weight_mem_banks_write_if_for_if_and_29_nl
      , weight_mem_banks_write_if_for_if_and_30_nl , weight_mem_banks_write_if_for_if_and_31_nl
      , weight_mem_banks_write_if_for_if_and_32_nl , weight_mem_banks_write_if_for_if_and_33_nl
      , weight_mem_banks_write_if_for_if_and_34_nl});
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_1_nl = MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3,
      (weight_read_addrs_1_lpi_1_dfm_1[3]), (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_3_lpi_1_dfm_1[3]), (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]),
      (weight_read_addrs_5_lpi_1_dfm_1[3]), (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_7_lpi_1_dfm_1[3]), {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_2
      , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_1 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_20_0});
  assign weight_mem_banks_write_if_for_if_mux_6_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_1_nl,
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a0_a1_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_4_nl
      , weight_mem_banks_write_if_for_if_mux_6_nl};
  assign nor_462_nl = ~(PECore_UpdateFSM_switch_lp_equal_tmp_2_3 | (~ PECore_RunMac_PECore_RunMac_if_and_svs_st_3));
  assign mux_255_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp,
      nor_462_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_pff = mux_255_nl & while_stage_0_5;
  assign weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_pff = and_dcpl_181;
  assign weight_mem_banks_bank_a0_a1_a0_a_rsci_d_d = {weight_write_data_data_0_7_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_6_lpi_1_dfm_1_2_6 , weight_write_data_data_0_5_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_4_lpi_1_dfm_1_2_6 , weight_write_data_data_0_3_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_2_lpi_1_dfm_1_2_6 , weight_write_data_data_0_1_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_0_lpi_1_dfm_1_2_6};
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_3_nl
      = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1
      | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0));
  assign weight_mem_banks_write_if_for_if_and_21_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_22_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_23_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_24_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_25_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_26_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_27_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1 & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_3_nl
      = MUX1HOT_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
      {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_3_nl
      , weight_mem_banks_write_if_for_if_and_21_nl , weight_mem_banks_write_if_for_if_and_22_nl
      , weight_mem_banks_write_if_for_if_and_23_nl , weight_mem_banks_write_if_for_if_and_24_nl
      , weight_mem_banks_write_if_for_if_and_25_nl , weight_mem_banks_write_if_for_if_and_26_nl
      , weight_mem_banks_write_if_for_if_and_27_nl});
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_2_nl = MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3,
      (weight_read_addrs_1_lpi_1_dfm_1[3]), (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_3_lpi_1_dfm_1[3]), (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]),
      (weight_read_addrs_5_lpi_1_dfm_1[3]), (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_7_lpi_1_dfm_1[3]), {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_2
      , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_1 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_22_0});
  assign weight_mem_banks_write_if_for_if_mux_5_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_2_nl,
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a1_a0_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_3_nl
      , weight_mem_banks_write_if_for_if_mux_5_nl};
  assign nor_461_nl = ~((~ PECore_RunScale_PECore_RunScale_if_and_1_svs_3) | ProductSum_for_asn_16_itm_3);
  assign mux_254_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp,
      nor_461_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_pff = mux_254_nl & while_stage_0_5;
  assign weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_pff = and_dcpl_184;
  assign weight_mem_banks_bank_a0_a1_a1_a_rsci_d_d = {weight_write_data_data_0_7_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_6_lpi_1_dfm_1_2_6 , weight_write_data_data_0_5_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_4_lpi_1_dfm_1_2_6 , weight_write_data_data_0_3_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_2_lpi_1_dfm_1_2_6 , weight_write_data_data_0_1_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_0_lpi_1_dfm_1_2_6};
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_2_nl
      = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1
      | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0));
  assign weight_mem_banks_write_if_for_if_and_14_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_15_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_16_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_17_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_18_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_19_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_20_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1 & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_2_nl
      = MUX1HOT_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
      {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_2_nl
      , weight_mem_banks_write_if_for_if_and_14_nl , weight_mem_banks_write_if_for_if_and_15_nl
      , weight_mem_banks_write_if_for_if_and_16_nl , weight_mem_banks_write_if_for_if_and_17_nl
      , weight_mem_banks_write_if_for_if_and_18_nl , weight_mem_banks_write_if_for_if_and_19_nl
      , weight_mem_banks_write_if_for_if_and_20_nl});
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_3_nl = MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3,
      (weight_read_addrs_1_lpi_1_dfm_1[3]), (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_3_lpi_1_dfm_1[3]), (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]),
      (weight_read_addrs_5_lpi_1_dfm_1[3]), (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_7_lpi_1_dfm_1[3]), {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_2
      , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_1 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_24_0});
  assign weight_mem_banks_write_if_for_if_mux_4_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_3_nl,
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a1_a1_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_2_nl
      , weight_mem_banks_write_if_for_if_mux_4_nl};
  assign nor_460_nl = ~((~ PECore_RunScale_PECore_RunScale_if_and_1_svs_st_3) | ProductSum_for_asn_25_itm_3);
  assign mux_253_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp,
      nor_460_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_pff = mux_253_nl & while_stage_0_5;
  assign weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_pff = and_dcpl_187;
  assign weight_mem_banks_bank_a1_a0_a0_a_rsci_d_d = {weight_write_data_data_0_7_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_6_lpi_1_dfm_1_2_6 , weight_write_data_data_0_5_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_4_lpi_1_dfm_1_2_6 , weight_write_data_data_0_3_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_2_lpi_1_dfm_1_2_6 , weight_write_data_data_0_1_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_0_lpi_1_dfm_1_2_6};
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_1_nl
      = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1
      | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0));
  assign weight_mem_banks_write_if_for_if_and_7_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_8_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_9_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_10_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_11_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_12_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_13_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1 & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_1_nl
      = MUX1HOT_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
      {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_1_nl
      , weight_mem_banks_write_if_for_if_and_7_nl , weight_mem_banks_write_if_for_if_and_8_nl
      , weight_mem_banks_write_if_for_if_and_9_nl , weight_mem_banks_write_if_for_if_and_10_nl
      , weight_mem_banks_write_if_for_if_and_11_nl , weight_mem_banks_write_if_for_if_and_12_nl
      , weight_mem_banks_write_if_for_if_and_13_nl});
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_4_nl = MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3,
      (weight_read_addrs_1_lpi_1_dfm_1[3]), (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_3_lpi_1_dfm_1[3]), (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]),
      (weight_read_addrs_5_lpi_1_dfm_1[3]), (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_7_lpi_1_dfm_1[3]), {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_2
      , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_1 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_26_0});
  assign weight_mem_banks_write_if_for_if_mux_3_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_4_nl,
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a1_a0_a0_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_1_nl
      , weight_mem_banks_write_if_for_if_mux_3_nl};
  assign nor_459_nl = ~((~ weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_1)
      | ProductSum_for_asn_42_itm_3);
  assign mux_252_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp,
      nor_459_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_pff = mux_252_nl & while_stage_0_5;
  assign weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_pff = and_dcpl_190;
  assign weight_mem_banks_bank_a1_a0_a1_a_rsci_d_d = {weight_write_data_data_0_7_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_6_lpi_1_dfm_1_2_6 , weight_write_data_data_0_5_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_4_lpi_1_dfm_1_2_6 , weight_write_data_data_0_3_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_2_lpi_1_dfm_1_2_6 , weight_write_data_data_0_1_lpi_1_dfm_1_2_6
      , weight_write_data_data_0_0_lpi_1_dfm_1_2_6};
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_nl
      = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1
      | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0));
  assign weight_mem_banks_write_if_for_if_and_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_1_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_2_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_3_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2
      & (~(weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1 | weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0))
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_4_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_5_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1 & (~ weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_and_6_nl = weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2
      & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1 & weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_nl
      = MUX1HOT_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
      (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
      {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_or_nl ,
      weight_mem_banks_write_if_for_if_and_nl , weight_mem_banks_write_if_for_if_and_1_nl
      , weight_mem_banks_write_if_for_if_and_2_nl , weight_mem_banks_write_if_for_if_and_3_nl
      , weight_mem_banks_write_if_for_if_and_4_nl , weight_mem_banks_write_if_for_if_and_5_nl
      , weight_mem_banks_write_if_for_if_and_6_nl});
  assign weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_5_nl = MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3,
      (weight_read_addrs_1_lpi_1_dfm_1[3]), (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_3_lpi_1_dfm_1[3]), (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]),
      (weight_read_addrs_5_lpi_1_dfm_1[3]), (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]),
      (weight_read_addrs_7_lpi_1_dfm_1[3]), {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_2
      , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_1 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_28_0});
  assign weight_mem_banks_write_if_for_if_mux_2_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_if_1_mux_5_nl,
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a1_a0_a1_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_weight_mem_banks_write_if_for_if_mux1h_nl
      , weight_mem_banks_write_if_for_if_mux_2_nl};
  assign nor_458_nl = ~((~ weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_1)
      | ProductSum_for_asn_51_itm_3);
  assign mux_251_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp,
      nor_458_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_pff = mux_251_nl & while_stage_0_5;
  assign weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_pff = and_dcpl_193;
  assign weight_mem_banks_bank_a1_a1_a0_a_rsci_d_d = {weight_write_data_data_0_7_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_6_lpi_1_dfm_1_3_2 , weight_write_data_data_0_5_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_4_lpi_1_dfm_1_3_2 , weight_write_data_data_0_3_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_2_lpi_1_dfm_1_3_2 , weight_write_data_data_0_1_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_0_lpi_1_dfm_1_3_2};
  assign weight_mem_banks_write_if_for_if_mux_1_nl = MUX_v_11_2_2(weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_11_1,
      weight_read_addrs_0_14_4_lpi_1_dfm_1_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_banks_write_if_for_if_mux_54_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_0,
      weight_read_addrs_4_14_2_lpi_1_dfm_2_0, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_banks_bank_a1_a1_a0_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_mux_1_nl
      , weight_mem_banks_write_if_for_if_mux_54_nl};
  assign nor_457_nl = ~((~ weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_2)
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_44_itm_1);
  assign mux_250_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1,
      nor_457_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_pff = mux_250_nl & while_stage_0_6;
  assign weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_pff = weight_write_addrs_lpi_1_dfm_1_3_14_3;
  assign weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_pff = and_dcpl_469;
  assign weight_mem_banks_bank_a1_a1_a1_a_rsci_d_d = {weight_write_data_data_0_7_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_6_lpi_1_dfm_1_3_2 , weight_write_data_data_0_5_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_4_lpi_1_dfm_1_3_2 , weight_write_data_data_0_3_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_2_lpi_1_dfm_1_3_2 , weight_write_data_data_0_1_lpi_1_dfm_1_3_2
      , weight_write_data_data_0_0_lpi_1_dfm_1_3_2};
  assign weight_mem_banks_write_if_for_if_mux_nl = MUX_v_11_2_2(weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_11_1,
      weight_read_addrs_0_14_4_lpi_1_dfm_1_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_banks_write_if_for_if_mux_53_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_0,
      weight_read_addrs_slc_weight_read_addrs_0_3_0_3_23_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_banks_bank_a1_a1_a1_a_rsci_radr_d = {weight_mem_banks_write_if_for_if_mux_nl
      , weight_mem_banks_write_if_for_if_mux_53_nl};
  assign nor_456_nl = ~((~ weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_2)
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_54_itm_1);
  assign mux_249_nl = MUX_s_1_2_2(weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1,
      nor_456_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_pff = mux_249_nl & while_stage_0_6;
  assign weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_pff = and_dcpl_467;
  assign or_dcpl_679 = ((weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]) & and_dcpl_580)
      | ((weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]) & and_dcpl_584) | ((weight_mem_write_arbxbar_xbar_for_empty_sva_2[2])
      & and_dcpl_582);
  assign nor_tmp = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0])
      & (weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]);
  assign and_dcpl_664 = (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_1_itm_2[1])
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_62_itm_1;
  assign or_dcpl_683 = and_dcpl_664 | ((pe_manager_base_weight_slc_pe_manager_base_weight_1_0_1_itm_2[0])
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_79_itm_1);
  assign and_dcpl_665 = (pe_manager_base_weight_slc_pe_manager_base_weight_1_0_1_itm_2[0])
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_47_itm_1;
  assign or_dcpl_684 = and_dcpl_664 | and_dcpl_665;
  assign PECore_DecodeAxiRead_switch_lp_mux_23_nl = MUX_s_1_2_2((SC_SRAM_CONFIG[0]),
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_9,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_21_nl
      = PECore_DecodeAxiRead_switch_lp_mux_23_nl & PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign rva_out_reg_data_mux_20_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_21_nl,
      rva_out_reg_data_0_sva_dfm_6, rva_in_reg_rw_sva_9);
  assign PECore_PushAxiRsp_if_else_mux_14_itm = MUX_s_1_2_2(rva_out_reg_data_mux_20_nl,
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_2,
      input_read_req_valid_lpi_1_dfm_1_9);
  assign PECore_DecodeAxiRead_switch_lp_mux_24_nl = MUX_s_1_2_2((SC_SRAM_CONFIG[8]),
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_9,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_22_nl
      = PECore_DecodeAxiRead_switch_lp_mux_24_nl & PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign rva_out_reg_data_mux_21_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_22_nl,
      rva_out_reg_data_8_sva_dfm_6, rva_in_reg_rw_sva_9);
  assign PECore_PushAxiRsp_if_else_mux_15_itm = MUX_s_1_2_2(rva_out_reg_data_mux_21_nl,
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_2,
      input_read_req_valid_lpi_1_dfm_1_9);
  assign PECore_DecodeAxiRead_switch_lp_mux_25_nl = MUX_s_1_2_2((SC_SRAM_CONFIG[16]),
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_7,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_23_nl
      = PECore_DecodeAxiRead_switch_lp_mux_25_nl & PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign rva_out_reg_data_mux_22_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_23_nl,
      rva_out_reg_data_16_sva_dfm_6, rva_in_reg_rw_sva_9);
  assign PECore_PushAxiRsp_if_else_mux_16_itm = MUX_s_1_2_2(rva_out_reg_data_mux_22_nl,
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_2,
      input_read_req_valid_lpi_1_dfm_1_9);
  assign PECore_DecodeAxiRead_switch_lp_mux_26_nl = MUX_s_1_2_2((SC_SRAM_CONFIG[24]),
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_7,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_25_nl
      = PECore_DecodeAxiRead_switch_lp_mux_26_nl & PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign rva_out_reg_data_mux_24_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_25_nl,
      rva_out_reg_data_24_sva_dfm_6, rva_in_reg_rw_sva_9);
  assign PECore_PushAxiRsp_if_else_mux_17_nl = MUX_s_1_2_2(rva_out_reg_data_mux_24_nl,
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_2,
      input_read_req_valid_lpi_1_dfm_1_9);
  assign PECore_PushAxiRsp_if_mux1h_15 = MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_17_nl,
      (reg_weight_port_read_out_data_0_3_sva_dfm_4_ftd_2[0]), crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_24_nl
      = (SC_SRAM_CONFIG[31]) & (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8) &
      PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign rva_out_reg_data_mux_23_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_24_nl,
      rva_out_reg_data_31_sva_dfm_6, rva_in_reg_rw_sva_9);
  assign PECore_PushAxiRsp_if_else_mux_18_nl = MUX_s_1_2_2(rva_out_reg_data_mux_23_nl,
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_2,
      input_read_req_valid_lpi_1_dfm_1_9);
  assign PECore_PushAxiRsp_if_mux1h_17 = MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_18_nl,
      reg_weight_port_read_out_data_0_3_sva_dfm_4_ftd, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7);
  assign or_3652_cse = (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1]) | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_80_itm_1;
  assign or_3651_cse = (~ (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1])) | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_80_itm_1;
  assign or_3650_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_cse
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_80_itm_1;
  assign mux_1254_nl = MUX_s_1_2_2(or_3652_cse, or_3651_cse, reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[2]);
  assign mux_1255_nl = MUX_s_1_2_2(mux_1254_nl, or_3650_cse, reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[0]);
  assign or_3653_cse = or_tmp_2755 | (crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3
      & mux_1255_nl);
  assign or_3659_cse = (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1]) | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_10_itm_1;
  assign or_3658_cse = (~ (reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[1])) | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_10_itm_1;
  assign or_3657_cse = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_cse
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_10_itm_1;
  assign weight_port_read_out_data_and_106_enex5 = weight_port_read_out_data_and_92_cse
      & reg_weight_port_read_out_data_0_2_sva_dfm_2_2_enexo;
  assign weight_port_read_out_data_and_42_ssc = PECoreRun_wen & (while_and_1123_rgt
      | while_and_24_cse) & while_stage_0_7;
  assign mux_1265_nl = MUX_s_1_2_2(not_tmp_1925, or_tmp_2778, or_3652_cse);
  assign mux_1264_nl = MUX_s_1_2_2(not_tmp_1925, or_tmp_2778, or_3651_cse);
  assign mux_1266_nl = MUX_s_1_2_2(mux_1265_nl, mux_1264_nl, reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[2]);
  assign mux_1263_nl = MUX_s_1_2_2(not_tmp_1925, or_tmp_2778, or_3650_cse);
  assign mux_1267_nl = MUX_s_1_2_2(mux_1266_nl, mux_1263_nl, reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[0]);
  assign mux_1268_cse = MUX_s_1_2_2(not_tmp_1925, mux_1267_nl, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign or_3670_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_44_itm_2
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_71_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_60_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_47_itm_1;
  assign mux_1269_nl = MUX_s_1_2_2(mux_1268_cse, or_tmp_2778, or_3670_nl);
  assign and_2218_cse = mux_1269_nl & weight_mem_run_3_for_aelse_and_cse;
  assign weight_port_read_out_data_and_107_enex5 = weight_port_read_out_data_and_92_cse
      & reg_weight_port_read_out_data_0_3_sva_dfm_2_2_enexo;
  assign rva_out_reg_data_and_115_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_46_40_sva_dfm_4_2_1_enexo;
  assign rva_out_reg_data_and_116_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_55_48_sva_dfm_4_2_enexo;
  assign rva_out_reg_data_and_117_enex5 = input_read_req_valid_and_1_cse & reg_rva_out_reg_data_55_48_sva_dfm_4_2_1_enexo;
  assign weight_port_read_out_data_and_96_ssc = PECoreRun_wen & and_dcpl_293 & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_4
      & while_stage_0_8;
  assign weight_port_read_out_data_and_108_enex5 = weight_port_read_out_data_and_96_ssc
      & reg_weight_port_read_out_data_0_0_sva_dfm_1_2_enexo;
  assign weight_port_read_out_data_and_109_enex5 = weight_port_read_out_data_and_96_ssc
      & reg_weight_port_read_out_data_0_1_sva_dfm_1_2_enexo;
  assign weight_port_read_out_data_and_110_enex5 = weight_port_read_out_data_and_96_ssc
      & reg_weight_port_read_out_data_0_2_sva_dfm_1_2_enexo;
  assign weight_port_read_out_data_and_111_enex5 = weight_port_read_out_data_and_96_ssc
      & reg_weight_port_read_out_data_0_3_sva_dfm_1_2_enexo;
  assign rva_out_reg_data_and_118_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_46_40_sva_dfm_4_1_1_enexo;
  assign rva_out_reg_data_and_119_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_55_48_sva_dfm_4_1_enexo;
  assign rva_out_reg_data_and_120_enex5 = input_read_req_valid_and_2_cse & reg_rva_out_reg_data_55_48_sva_dfm_4_1_1_enexo;
  assign mux_174_nl = MUX_s_1_2_2(while_and_24_cse, or_tmp_3, PECore_RunMac_PECore_RunMac_if_and_svs_st_5);
  assign mux_175_nl = MUX_s_1_2_2(mux_174_nl, (~ or_tmp_2), rva_in_reg_rw_sva_st_1_5);
  assign weight_port_read_out_data_and_100_ssc = PECoreRun_wen & mux_175_nl & while_stage_0_7;
  assign weight_port_read_out_data_0_0_sva_dfm_3_7 = MUX1HOT_s_1_9_2(weight_port_read_out_data_0_0_sva_dfm_2_7,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[7]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[7]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[7]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[7]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[7]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[7]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[7]), (BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9[7]),
      {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , weight_mem_run_3_for_5_and_161_cse
      , weight_mem_run_3_for_5_and_162_itm_2 , reg_weight_mem_run_3_for_5_and_163_itm_2_cse
      , weight_mem_run_3_for_5_and_164_itm_2 , reg_weight_mem_run_3_for_5_and_165_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_166_itm_2_cse , reg_weight_mem_run_3_for_5_and_167_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_168_itm_2_cse});
  assign weight_port_read_out_data_0_0_sva_dfm_3_6_0 = MUX1HOT_v_7_9_2(weight_port_read_out_data_0_0_sva_dfm_2_6_0,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[6:0]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[6:0]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[6:0]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[6:0]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[6:0]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[6:0]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[6:0]), (BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9[6:0]),
      {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , weight_mem_run_3_for_5_and_161_cse
      , weight_mem_run_3_for_5_and_162_itm_2 , reg_weight_mem_run_3_for_5_and_163_itm_2_cse
      , weight_mem_run_3_for_5_and_164_itm_2 , reg_weight_mem_run_3_for_5_and_165_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_166_itm_2_cse , reg_weight_mem_run_3_for_5_and_167_itm_2_cse
      , reg_weight_mem_run_3_for_5_and_168_itm_2_cse});
  assign weight_mem_run_3_for_5_and_179_ssc = reg_weight_mem_run_3_for_5_and_166_itm_2_cse
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_a_mx1_7 = MUX1HOT_s_1_9_2(weight_port_read_out_data_0_1_sva_dfm_2_7,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[15]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[15]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[15]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[15]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[15]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[15]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[15]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[7]),
      {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , weight_mem_run_3_for_5_and_161_cse
      , weight_mem_run_3_for_5_and_175_cse , weight_mem_run_3_for_5_and_176_cse ,
      weight_mem_run_3_for_5_and_177_cse , weight_mem_run_3_for_5_and_178_cse , weight_mem_run_3_for_5_and_179_ssc
      , weight_mem_run_3_for_5_and_180_cse , weight_mem_run_3_for_5_and_181_cse});
  assign PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_a_mx1_6_0 = MUX1HOT_v_7_9_2(weight_port_read_out_data_0_1_sva_dfm_2_6_0,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[14:8]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[14:8]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[14:8]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[14:8]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[14:8]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[14:8]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[14:8]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[6:0]),
      {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , weight_mem_run_3_for_5_and_161_cse
      , weight_mem_run_3_for_5_and_175_cse , weight_mem_run_3_for_5_and_176_cse ,
      weight_mem_run_3_for_5_and_177_cse , weight_mem_run_3_for_5_and_178_cse , weight_mem_run_3_for_5_and_179_ssc
      , weight_mem_run_3_for_5_and_180_cse , weight_mem_run_3_for_5_and_181_cse});
  assign weight_mem_run_3_for_5_and_182_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_3
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_mem_run_3_for_5_and_187_ssc = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_itm_2
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign weight_port_read_out_data_0_7_sva_dfm_1_1_mx0_7 = MUX1HOT_s_1_9_2(weight_port_read_out_data_0_7_sva_dfm_2_7,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[63]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[63]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[63]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[63]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[63]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[63]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[63]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[55]),
      {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , weight_mem_run_3_for_5_and_182_ssc
      , weight_mem_run_3_for_5_and_175_cse , weight_mem_run_3_for_5_and_176_cse ,
      weight_mem_run_3_for_5_and_177_cse , weight_mem_run_3_for_5_and_178_cse , weight_mem_run_3_for_5_and_187_ssc
      , weight_mem_run_3_for_5_and_180_cse , weight_mem_run_3_for_5_and_181_cse});
  assign weight_port_read_out_data_0_7_sva_dfm_1_1_mx0_6_0 = MUX1HOT_v_7_9_2(weight_port_read_out_data_0_7_sva_dfm_2_6_0,
      (input_mem_banks_read_read_data_lpi_1_dfm_1_4[62:56]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[62:56]),
      (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[62:56]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[62:56]),
      (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[62:56]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[62:56]),
      (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[62:56]), (weight_mem_banks_read_1_read_data_lpi_1_dfm_63_8_mx0[54:48]),
      {(~ weight_mem_run_3_for_land_1_lpi_1_dfm_3) , weight_mem_run_3_for_5_and_182_ssc
      , weight_mem_run_3_for_5_and_175_cse , weight_mem_run_3_for_5_and_176_cse ,
      weight_mem_run_3_for_5_and_177_cse , weight_mem_run_3_for_5_and_178_cse , weight_mem_run_3_for_5_and_187_ssc
      , weight_mem_run_3_for_5_and_180_cse , weight_mem_run_3_for_5_and_181_cse});
  assign rva_out_reg_data_55_48_sva_dfm_6_mx1_7_4 = MUX_v_4_2_2(rva_out_reg_data_55_48_sva_dfm_4_1_7_4,
      rva_out_reg_data_55_48_sva_dfm_6_rsp_0, or_dcpl_665);
  assign rva_out_reg_data_55_48_sva_dfm_6_mx1_3_0 = MUX_v_4_2_2(rva_out_reg_data_55_48_sva_dfm_4_1_3_0,
      rva_out_reg_data_55_48_sva_dfm_6_rsp_1, or_dcpl_665);
  assign rva_out_reg_data_46_40_sva_dfm_6_mx1_6_4 = MUX_v_3_2_2(rva_out_reg_data_46_40_sva_dfm_4_1_6_4,
      rva_out_reg_data_46_40_sva_dfm_6_rsp_0, or_dcpl_665);
  assign rva_out_reg_data_46_40_sva_dfm_6_mx1_3_0 = MUX_v_4_2_2(rva_out_reg_data_46_40_sva_dfm_4_1_3_0,
      rva_out_reg_data_46_40_sva_dfm_6_rsp_1, or_dcpl_665);
  assign rva_out_reg_data_39_36_sva_dfm_6_mx1_3 = MUX_s_1_2_2(rva_out_reg_data_39_36_sva_dfm_4_1_3,
      rva_out_reg_data_39_36_sva_dfm_6_rsp_0, or_dcpl_665);
  assign rva_out_reg_data_39_36_sva_dfm_6_mx1_2 = MUX_s_1_2_2(rva_out_reg_data_39_36_sva_dfm_4_1_2,
      rva_out_reg_data_39_36_sva_dfm_6_rsp_1, or_dcpl_665);
  assign rva_out_reg_data_39_36_sva_dfm_6_mx1_1_0 = MUX_v_2_2_2(rva_out_reg_data_39_36_sva_dfm_4_1_1_0,
      rva_out_reg_data_39_36_sva_dfm_6_rsp_2, or_dcpl_665);
  assign weight_port_read_out_data_and_112_enex5 = weight_port_read_out_data_and_68_cse
      & reg_weight_port_read_out_data_0_0_sva_dfm_3_2_enexo;
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_16_nl
      = (SC_SRAM_CONFIG[7]) & (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8) &
      PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign PECore_PushAxiRsp_if_mux1h_10_6 = MUX1HOT_s_1_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_16_nl,
      rva_out_reg_data_7_1_sva_dfm_6_rsp_0, (input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2[6]),
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_1_ftd,
      {PECore_PushAxiRsp_if_asn_55 , PECore_PushAxiRsp_if_asn_57 , PECore_PushAxiRsp_if_asn_59
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7});
  assign PECore_DecodeAxiRead_switch_lp_mux_20_nl = MUX_s_1_2_2((SC_SRAM_CONFIG[15]),
      (rva_out_reg_data_15_9_sva_dfm_9[6]), PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_14_nl
      = PECore_DecodeAxiRead_switch_lp_mux_20_nl & PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign PECore_PushAxiRsp_if_mux1h_12_6 = MUX1HOT_s_1_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_14_nl,
      rva_out_reg_data_15_9_sva_dfm_6_rsp_0, (input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2[6]),
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_1_ftd,
      {PECore_PushAxiRsp_if_asn_55 , PECore_PushAxiRsp_if_asn_57 , PECore_PushAxiRsp_if_asn_59
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7});
  assign PECore_DecodeAxiRead_switch_lp_mux_21_nl = MUX_s_1_2_2((SC_SRAM_CONFIG[23]),
      (rva_out_reg_data_23_17_sva_dfm_7[6]), PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_11_nl
      = PECore_DecodeAxiRead_switch_lp_mux_21_nl & PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign PECore_PushAxiRsp_if_mux1h_14_6 = MUX1HOT_s_1_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_11_nl,
      rva_out_reg_data_23_17_sva_dfm_6_rsp_0, (input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2[6]),
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_ftd,
      {PECore_PushAxiRsp_if_asn_55 , PECore_PushAxiRsp_if_asn_57 , PECore_PushAxiRsp_if_asn_59
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7});
  assign PECore_DecodeAxiRead_switch_lp_mux_28_nl = MUX_s_1_2_2((SC_SRAM_CONFIG[22]),
      (rva_out_reg_data_23_17_sva_dfm_7[5]), PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_28_nl
      = PECore_DecodeAxiRead_switch_lp_mux_28_nl & PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign PECore_PushAxiRsp_if_mux1h_14_5 = MUX1HOT_s_1_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_28_nl,
      rva_out_reg_data_23_17_sva_dfm_6_rsp_1, (input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2[5]),
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_ftd_1,
      {PECore_PushAxiRsp_if_asn_55 , PECore_PushAxiRsp_if_asn_57 , PECore_PushAxiRsp_if_asn_59
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7});
  assign PECore_DecodeAxiRead_switch_lp_mux_29_nl = MUX_v_5_2_2((SC_SRAM_CONFIG[21:17]),
      (rva_out_reg_data_23_17_sva_dfm_7[4:0]), PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_29_nl
      = MUX_v_5_2_2(5'b00000, PECore_DecodeAxiRead_switch_lp_mux_29_nl, PECore_DecodeAxiRead_switch_lp_nor_9_cse_1);
  assign PECore_PushAxiRsp_if_mux1h_14_4_0 = MUX1HOT_v_5_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_29_nl,
      rva_out_reg_data_23_17_sva_dfm_6_rsp_2, (input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2[4:0]),
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_ftd_2,
      {PECore_PushAxiRsp_if_asn_55 , PECore_PushAxiRsp_if_asn_57 , PECore_PushAxiRsp_if_asn_59
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7});
  assign PECore_DecodeAxiRead_switch_lp_mux_22_nl = MUX_v_3_2_2((SC_SRAM_CONFIG[30:28]),
      (rva_out_reg_data_30_25_sva_dfm_7[5:3]), PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_8_nl =
      MUX_v_3_2_2(3'b000, PECore_DecodeAxiRead_switch_lp_mux_22_nl, PECore_DecodeAxiRead_switch_lp_nor_9_cse_1);
  assign PECore_PushAxiRsp_if_mux1h_16_5_3 = MUX1HOT_v_3_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_8_nl,
      rva_out_reg_data_30_25_sva_dfm_6_rsp_0, (input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2[5:3]),
      reg_weight_port_read_out_data_0_3_sva_dfm_4_ftd_1, {PECore_PushAxiRsp_if_asn_55
      , PECore_PushAxiRsp_if_asn_57 , PECore_PushAxiRsp_if_asn_59 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7});
  assign PECore_DecodeAxiRead_switch_lp_mux_30_nl = MUX_v_3_2_2((SC_SRAM_CONFIG[27:25]),
      (rva_out_reg_data_30_25_sva_dfm_7[2:0]), PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_30_nl
      = MUX_v_3_2_2(3'b000, PECore_DecodeAxiRead_switch_lp_mux_30_nl, PECore_DecodeAxiRead_switch_lp_nor_9_cse_1);
  assign PECore_PushAxiRsp_if_mux1h_16_2_0 = MUX1HOT_v_3_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_30_nl,
      rva_out_reg_data_30_25_sva_dfm_6_rsp_1, (input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2[2:0]),
      (reg_weight_port_read_out_data_0_3_sva_dfm_4_ftd_2[3:1]), {PECore_PushAxiRsp_if_asn_55
      , PECore_PushAxiRsp_if_asn_57 , PECore_PushAxiRsp_if_asn_59 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7});
  assign weight_port_read_out_data_and_113_enex5 = weight_port_read_out_data_and_92_cse
      & reg_weight_port_read_out_data_0_0_sva_dfm_2_2_enexo;
  assign weight_port_read_out_data_and_114_enex5 = weight_port_read_out_data_and_92_cse
      & reg_weight_port_read_out_data_0_1_sva_dfm_2_2_enexo;
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_26_nl
      = (SC_SRAM_CONFIG[6]) & (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8) &
      PECore_DecodeAxiRead_switch_lp_nor_9_cse_1;
  assign PECore_PushAxiRsp_if_mux1h_10_5 = MUX1HOT_s_1_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_26_nl,
      rva_out_reg_data_7_1_sva_dfm_6_rsp_1_rsp_0, (input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2[5]),
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_1_ftd_1_rsp_0,
      {PECore_PushAxiRsp_if_asn_55 , PECore_PushAxiRsp_if_asn_57 , PECore_PushAxiRsp_if_asn_59
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7});
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_31_nl
      = (SC_SRAM_CONFIG[5:1]) & (signext_5_1(~ PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8))
      & ({{4{PECore_DecodeAxiRead_switch_lp_nor_9_cse_1}}, PECore_DecodeAxiRead_switch_lp_nor_9_cse_1});
  assign PECore_PushAxiRsp_if_mux1h_10_4_0 = MUX1HOT_v_5_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_31_nl,
      rva_out_reg_data_7_1_sva_dfm_6_rsp_1_rsp_1, (input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2[4:0]),
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_1_ftd_1_rsp_1,
      {PECore_PushAxiRsp_if_asn_55 , PECore_PushAxiRsp_if_asn_57 , PECore_PushAxiRsp_if_asn_59
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7});
  assign PECore_DecodeAxiRead_switch_lp_mux_27_nl = MUX_v_3_2_2((SC_SRAM_CONFIG[14:12]),
      (rva_out_reg_data_15_9_sva_dfm_9[5:3]), PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_27_nl
      = MUX_v_3_2_2(3'b000, PECore_DecodeAxiRead_switch_lp_mux_27_nl, PECore_DecodeAxiRead_switch_lp_nor_9_cse_1);
  assign PECore_PushAxiRsp_if_mux1h_12_5_3 = MUX1HOT_v_3_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_27_nl,
      rva_out_reg_data_15_9_sva_dfm_6_rsp_1_rsp_0, (input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2[5:3]),
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_1_ftd_1_rsp_0,
      {PECore_PushAxiRsp_if_asn_55 , PECore_PushAxiRsp_if_asn_57 , PECore_PushAxiRsp_if_asn_59
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7});
  assign PECore_DecodeAxiRead_switch_lp_mux_31_nl = MUX_v_3_2_2((SC_SRAM_CONFIG[11:9]),
      (rva_out_reg_data_15_9_sva_dfm_9[2:0]), PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_32_nl
      = MUX_v_3_2_2(3'b000, PECore_DecodeAxiRead_switch_lp_mux_31_nl, PECore_DecodeAxiRead_switch_lp_nor_9_cse_1);
  assign PECore_PushAxiRsp_if_mux1h_12_2_0 = MUX1HOT_v_3_4_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_32_nl,
      rva_out_reg_data_15_9_sva_dfm_6_rsp_1_rsp_1, (input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2[2:0]),
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_1_ftd_1_rsp_1,
      {PECore_PushAxiRsp_if_asn_55 , PECore_PushAxiRsp_if_asn_57 , PECore_PushAxiRsp_if_asn_59
      , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7});
  assign or_dcpl_717 = weight_mem_run_3_for_5_and_108_itm_1 | weight_mem_run_3_for_5_and_112_itm_1;
  assign or_dcpl_718 = weight_mem_run_3_for_5_and_111_itm_1 | weight_mem_run_3_for_5_and_110_itm_1;
  assign or_dcpl_727 = weight_mem_run_3_for_5_and_44_itm_2 | weight_mem_run_3_for_5_and_48_itm_1;
  assign or_tmp_720 = ((reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_cse
      | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_5_cse | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_cse
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_3 | Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_2
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_0)
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1) | ((reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_6_cse
      | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_5_cse | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_4_cse
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_3 | Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_2
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_0)
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1) | ((reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_cse
      | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_5_cse | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_cse
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_3 | Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_2
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_0)
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1) | ((Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_6
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_5 | Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_4
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_3 | Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_2
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_0)
      & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1);
  assign or_1480_nl = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_cse
      | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_5_cse | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_cse
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_3 | Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_2
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_0
      | or_tmp_720;
  assign mux_tmp_481 = MUX_s_1_2_2(or_tmp_720, or_1480_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1);
  assign or_1481_nl = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_cse
      | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_5_cse | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_cse
      | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_3_cse | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_2_cse
      | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_1_cse | Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_0
      | mux_tmp_481;
  assign mux_tmp_482 = MUX_s_1_2_2(mux_tmp_481, or_1481_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1);
  assign or_1482_nl = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_cse
      | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_5_cse | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4_cse
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_3 | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_2
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_0
      | mux_tmp_482;
  assign mux_tmp_483 = MUX_s_1_2_2(mux_tmp_482, or_1482_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1);
  assign and_dcpl_759 = while_stage_0_3 & fsm_output;
  assign or_dcpl_751 = weight_mem_run_3_for_5_and_111_itm_1 | weight_mem_run_3_for_5_and_102_itm_2;
  assign or_dcpl_779 = weight_mem_run_3_for_5_and_39_itm_2 | weight_mem_run_3_for_5_and_46_itm_2;
  assign or_dcpl_801 = weight_mem_run_3_for_5_and_31_itm_2 | weight_mem_run_3_for_5_and_30_itm_2;
  assign or_dcpl_824 = accum_vector_operator_1_for_asn_64_itm_7 | reg_PECore_RunMac_PECore_RunMac_if_and_svs_st_8_cse;
  assign and_dcpl_885 = fsm_output & while_stage_0_10;
  assign or_tmp_745 = PECore_RunMac_PECore_RunMac_if_and_svs_st_7 | accum_vector_operator_1_for_asn_70_itm_6;
  assign or_dcpl_826 = accum_vector_operator_1_for_asn_55_itm_7 | reg_PECore_RunMac_PECore_RunMac_if_and_svs_st_8_cse;
  assign or_tmp_762 = PECore_RunMac_PECore_RunMac_if_and_svs_st_7 | accum_vector_operator_1_for_asn_61_itm_6;
  assign or_dcpl_828 = reg_PECore_RunMac_PECore_RunMac_if_and_svs_st_8_cse | accum_vector_operator_1_for_asn_46_itm_7;
  assign or_tmp_779 = PECore_RunMac_PECore_RunMac_if_and_svs_st_7 | accum_vector_operator_1_for_asn_52_itm_6;
  assign or_tmp_796 = PECore_RunMac_PECore_RunMac_if_and_svs_st_7 | accum_vector_operator_1_for_asn_43_itm_6;
  assign or_tmp_830 = PECore_RunMac_PECore_RunMac_if_and_svs_st_7 | accum_vector_operator_1_for_asn_34_itm_6;
  assign or_tmp_864 = PECore_RunMac_PECore_RunMac_if_and_svs_st_7 | accum_vector_operator_1_for_asn_25_itm_6;
  assign or_tmp_915 = PECore_RunMac_PECore_RunMac_if_and_svs_st_7 | accum_vector_operator_1_for_asn_16_itm_6;
  assign or_tmp_949 = PECore_RunMac_PECore_RunMac_if_and_svs_st_7 | accum_vector_operator_1_for_asn_7_itm_6;
  assign and_dcpl_964 = fsm_output & while_stage_0_9;
  assign and_2590_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b11111111) & mux_773_cse;
  assign and_2591_nl = input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4==8'b11111111);
  assign mux_tmp_1225 = MUX_s_1_2_2(and_2590_nl, and_2591_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign or_tmp_2755 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_60_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_48_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_62_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_47_itm_1;
  assign or_tmp_2762 = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_72_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_48_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_62_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_79_itm_1;
  assign or_tmp_2778 = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      | weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign not_tmp_1925 = ~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
      | (~ weight_mem_run_3_for_land_1_lpi_1_dfm_3));
  assign data_in_tmp_operator_2_for_and_tmp = PECoreRun_wen & and_dcpl_32 & weight_mem_run_3_for_land_3_lpi_1_dfm_2;
  assign pe_manager_base_input_and_tmp = PECoreRun_wen & ((or_dcpl_87 & while_stage_0_3)
      | and_692_cse);
  assign rva_in_reg_data_and_tmp = PECoreRun_wen & and_dcpl_312 & (and_321_cse |
      (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  assign and_2435_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10100111))) & mux_773_cse;
  assign nor_1421_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:3]!=5'b10100)
      | nand_408_cse);
  assign mux_1076_nl = MUX_s_1_2_2(and_2435_nl, nor_1421_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1920_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1076_nl & and_dcpl_759
      & PECoreRun_wen;
  assign and_2337_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01010110))) & mux_773_cse;
  assign nor_1193_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01010110));
  assign mux_914_nl = MUX_s_1_2_2(and_2337_nl, nor_1193_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1677_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_914_nl & and_dcpl_759
      & PECoreRun_wen;
  assign and_2547_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11110010))) & mux_773_cse;
  assign nor_1638_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11110010));
  assign mux_1226_nl = MUX_s_1_2_2(and_2547_nl, nor_1638_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2145_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1226_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1414_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b1010010) |
      mux_799_cse);
  assign nor_1415_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10100101));
  assign mux_1072_nl = MUX_s_1_2_2(nor_1414_nl, nor_1415_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1914_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1072_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_277_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10111010))) &
      mux_773_cse);
  assign or_3244_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10111010);
  assign mux_1114_nl = MUX_s_1_2_2(nand_277_nl, or_3244_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1977_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_1114_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nand_184_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01101110))) &
      mux_773_cse);
  assign or_2782_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01101110);
  assign mux_962_nl = MUX_s_1_2_2(nand_184_nl, or_2782_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1749_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_962_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nand_278_nl = ~((PEManager_15U_GetInputAddr_acc_tmp==8'b10111011) & mux_773_cse);
  assign or_3250_nl = (~(input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]==6'b101110)))
      | nand_407_cse;
  assign mux_1116_nl = MUX_s_1_2_2(nand_278_nl, or_3250_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1980_tmp = (~((reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_return_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) | mux_1116_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign and_2560_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b11110110) & mux_773_cse;
  assign and_2561_nl = input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4==8'b11110110);
  assign mux_1234_nl = MUX_s_1_2_2(and_2560_nl, and_2561_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2157_tmp = (~(reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_return_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) & mux_1234_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1315_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10000001) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1316_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10000001));
  assign mux_1000_nl = MUX_s_1_2_2(nor_1315_nl, nor_1316_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1806_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1000_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_259_nl = ~((PEManager_15U_GetInputAddr_acc_tmp==8'b10101111) & mux_773_cse);
  assign or_3180_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:4]!=4'b1010)
      | nand_410_cse;
  assign mux_1092_nl = MUX_s_1_2_2(nand_259_nl, or_3180_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1944_tmp = (~((reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_return_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) | mux_1092_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nand_347_nl = ~((PEManager_15U_GetInputAddr_acc_tmp==8'b11101111) & mux_773_cse);
  assign or_3555_nl = (~(input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:4]==4'b1110)))
      | nand_410_cse;
  assign mux_1220_nl = MUX_s_1_2_2(nand_347_nl, or_3555_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2136_tmp = (~((reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_return_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) | mux_1220_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign and_2521_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11100011))) & mux_773_cse;
  assign nor_1593_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b111000)
      | nand_407_cse);
  assign mux_1196_nl = MUX_s_1_2_2(and_2521_nl, nor_1593_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2100_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1196_nl & and_dcpl_759
      & PECoreRun_wen;
  assign or_2952_nl = (PEManager_15U_GetInputAddr_acc_tmp!=8'b10001010) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse);
  assign or_2948_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10001010);
  assign mux_1018_nl = MUX_s_1_2_2(or_2952_nl, or_2948_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1833_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_1018_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nand_258_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10101110))) &
      mux_773_cse);
  assign or_3174_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10101110);
  assign mux_1090_nl = MUX_s_1_2_2(nand_258_nl, or_3174_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1941_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_1090_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign or_2162_nl = (PEManager_15U_GetInputAddr_acc_tmp!=8'b00001011) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse);
  assign or_2158_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b000010)
      | nand_407_cse;
  assign mux_764_nl = MUX_s_1_2_2(or_2162_nl, or_2158_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1452_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_764_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nand_147_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01001111))) &
      mux_773_cse);
  assign or_2590_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:4]!=4'b0100)
      | nand_410_cse;
  assign mux_900_nl = MUX_s_1_2_2(nand_147_nl, or_2590_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1656_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_900_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1153_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01000111) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1154_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:3]!=5'b01000)
      | nand_408_cse);
  assign mux_884_nl = MUX_s_1_2_2(nor_1153_nl, nor_1154_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1632_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_884_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1181_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01010010) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1182_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01010010));
  assign mux_906_nl = MUX_s_1_2_2(nor_1181_nl, nor_1182_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1665_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_906_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1223_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01100001) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1224_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01100001));
  assign mux_936_nl = MUX_s_1_2_2(nor_1223_nl, nor_1224_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1710_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_936_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_279_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10111100))) &
      mux_773_cse);
  assign or_3255_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10111100);
  assign mux_1118_nl = MUX_s_1_2_2(nand_279_nl, or_3255_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1983_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_1118_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1406_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10100010) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1407_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10100010));
  assign mux_1066_nl = MUX_s_1_2_2(nor_1406_nl, nor_1407_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1905_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1066_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_299_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11001101))) &
      mux_773_cse);
  assign or_3360_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11001101);
  assign mux_1152_nl = MUX_s_1_2_2(nand_299_nl, or_3360_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2034_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_1152_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nand_164_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01011101))) &
      mux_773_cse);
  assign or_2678_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01011101);
  assign mux_928_nl = MUX_s_1_2_2(nand_164_nl, or_2678_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1698_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_928_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign and_2306_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00110110))) & mux_773_cse;
  assign nor_1105_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00110110));
  assign mux_850_nl = MUX_s_1_2_2(and_2306_nl, nor_1105_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1581_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_850_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1062_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00100110) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1063_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00100110));
  assign mux_818_nl = MUX_s_1_2_2(nor_1062_nl, nor_1063_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1533_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_818_nl & and_dcpl_759
      & PECoreRun_wen;
  assign and_2469_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11000000))) & mux_773_cse;
  assign nor_1493_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11000000));
  assign mux_1126_nl = MUX_s_1_2_2(and_2469_nl, nor_1493_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1995_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1126_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1539_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b1101000) |
      mux_799_cse);
  assign nor_1540_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11010001));
  assign mux_1160_nl = MUX_s_1_2_2(nor_1539_nl, nor_1540_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2046_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1160_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_321_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11011100))) &
      mux_773_cse);
  assign or_3446_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11011100);
  assign mux_1182_nl = MUX_s_1_2_2(nand_321_nl, or_3446_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2079_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_1182_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign or_2959_nl = (PEManager_15U_GetInputAddr_acc_tmp!=8'b10001011) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse);
  assign or_2955_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b100010)
      | nand_407_cse;
  assign mux_1020_nl = MUX_s_1_2_2(or_2959_nl, or_2955_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1836_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_1020_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign and_2475_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11000100))) & mux_773_cse;
  assign nor_1505_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11000100));
  assign mux_1134_nl = MUX_s_1_2_2(and_2475_nl, nor_1505_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2007_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1134_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_301_nl = ~((PEManager_15U_GetInputAddr_acc_tmp==8'b11001111) & mux_773_cse);
  assign or_3371_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:4]!=4'b1100)
      | nand_410_cse;
  assign mux_1156_nl = MUX_s_1_2_2(nand_301_nl, or_3371_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2040_tmp = (~((reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_return_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) | mux_1156_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign and_2515_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11100000))) & mux_773_cse;
  assign nor_1585_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11100000));
  assign mux_1190_nl = MUX_s_1_2_2(and_2515_nl, nor_1585_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2091_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1190_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_298_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11001100))) &
      mux_773_cse);
  assign or_3354_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11001100);
  assign mux_1150_nl = MUX_s_1_2_2(nand_298_nl, or_3354_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2031_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_1150_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1096_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00110011) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1097_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b001100)
      | nand_407_cse);
  assign mux_844_nl = MUX_s_1_2_2(nor_1096_nl, nor_1097_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1572_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_844_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_144_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01001000))) &
      mux_773_cse);
  assign or_2544_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01001000);
  assign mux_886_nl = MUX_s_1_2_2(nand_144_nl, or_2544_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1635_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_886_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nand_185_nl = ~((PEManager_15U_GetInputAddr_acc_tmp==8'b01101111) & mux_773_cse);
  assign or_2788_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:4]!=4'b0110)
      | nand_410_cse;
  assign mux_964_nl = MUX_s_1_2_2(nand_185_nl, or_2788_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1752_tmp = (~((reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_return_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) | mux_964_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nor_967_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00000010) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_968_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00000010));
  assign mux_746_nl = MUX_s_1_2_2(nor_967_nl, nor_968_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1425_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_746_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1229_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01100011) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1230_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b011000)
      | nand_407_cse);
  assign mux_940_nl = MUX_s_1_2_2(nor_1229_nl, nor_1230_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1716_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_940_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1135_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01000001) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1136_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01000001));
  assign mux_872_nl = MUX_s_1_2_2(nor_1135_nl, nor_1136_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1614_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_872_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1234_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b0110010) |
      mux_799_cse);
  assign nor_1235_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01100101));
  assign mux_944_nl = MUX_s_1_2_2(nor_1234_nl, nor_1235_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1722_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_944_nl & and_dcpl_759
      & PECoreRun_wen;
  assign and_2303_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00110100))) & mux_773_cse;
  assign nor_1100_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00110100));
  assign mux_846_nl = MUX_s_1_2_2(and_2303_nl, nor_1100_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1575_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_846_nl & and_dcpl_759
      & PECoreRun_wen;
  assign and_2453_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10110110))) & mux_773_cse;
  assign nor_1463_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10110110));
  assign mux_1106_nl = MUX_s_1_2_2(and_2453_nl, nor_1463_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1965_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1106_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_183_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01101101))) &
      mux_773_cse);
  assign or_2777_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01101101);
  assign mux_960_nl = MUX_s_1_2_2(nand_183_nl, or_2777_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1746_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_960_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nand_131_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00111100))) &
      mux_773_cse);
  assign or_2471_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00111100);
  assign mux_862_nl = MUX_s_1_2_2(nand_131_nl, or_2471_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1599_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_862_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1184_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01010011) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1185_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b010100)
      | nand_407_cse);
  assign mux_908_nl = MUX_s_1_2_2(nor_1184_nl, nor_1185_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1668_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_908_nl & and_dcpl_759
      & PECoreRun_wen;
  assign and_2499_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11010110))) & mux_773_cse;
  assign nor_1555_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11010110));
  assign mux_1170_nl = MUX_s_1_2_2(and_2499_nl, nor_1555_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2061_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1170_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1047_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00100001) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1048_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00100001));
  assign mux_808_nl = MUX_s_1_2_2(nor_1047_nl, nor_1048_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1518_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_808_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1022_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00010111) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1023_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:3]!=5'b00010)
      | nand_408_cse);
  assign mux_788_nl = MUX_s_1_2_2(nor_1022_nl, nor_1023_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1488_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_788_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_257_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10101101))) &
      mux_773_cse);
  assign or_3169_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10101101);
  assign mux_1088_nl = MUX_s_1_2_2(nand_257_nl, or_3169_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1938_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_1088_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign or_2974_nl = (PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b1000110) | mux_799_cse;
  assign or_2967_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10001101);
  assign mux_1024_nl = MUX_s_1_2_2(or_2974_nl, or_2967_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1842_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_1024_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign and_2367_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01110010))) & mux_773_cse;
  assign nor_1271_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01110010));
  assign mux_970_nl = MUX_s_1_2_2(and_2367_nl, nor_1271_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1761_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_970_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_344_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11101100))) &
      mux_773_cse);
  assign or_3538_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11101100);
  assign mux_1214_nl = MUX_s_1_2_2(nand_344_nl, or_3538_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2127_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_1214_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nand_346_nl = ~((PEManager_15U_GetInputAddr_acc_tmp==8'b11101110) & mux_773_cse);
  assign nand_486_nl = ~(input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4==8'b11101110));
  assign mux_1218_nl = MUX_s_1_2_2(nand_346_nl, nand_486_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2133_tmp = (~((reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_return_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) | mux_1218_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign and_2417_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10010111))) & mux_773_cse;
  assign nor_1376_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:3]!=5'b10010)
      | nand_408_cse);
  assign mux_1044_nl = MUX_s_1_2_2(and_2417_nl, nor_1376_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1872_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1044_nl & and_dcpl_759
      & PECoreRun_wen;
  assign and_2551_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b11110011) & mux_773_cse;
  assign nor_1641_nl = ~((~(input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]==6'b111100)))
      | nand_407_cse);
  assign mux_1228_nl = MUX_s_1_2_2(and_2551_nl, nor_1641_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2148_tmp = (~(reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_return_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) & mux_1228_nl & and_dcpl_759
      & PECoreRun_wen;
  assign and_2556_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b11110101) & mux_773_cse;
  assign and_2557_nl = input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4==8'b11110101);
  assign mux_1232_nl = MUX_s_1_2_2(and_2556_nl, and_2557_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2154_tmp = (~(reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_return_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) & mux_1232_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1321_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10000011) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1322_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b100000)
      | nand_407_cse);
  assign mux_1004_nl = MUX_s_1_2_2(nor_1321_nl, nor_1322_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1812_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1004_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_165_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01011110))) &
      mux_773_cse);
  assign or_2683_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01011110);
  assign mux_930_nl = MUX_s_1_2_2(nand_165_nl, or_2683_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1701_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_930_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign and_2518_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11100010))) & mux_773_cse;
  assign nor_1590_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11100010));
  assign mux_1194_nl = MUX_s_1_2_2(and_2518_nl, nor_1590_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2097_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1194_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_253_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10101000))) &
      mux_773_cse);
  assign or_3137_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10101000);
  assign mux_1078_nl = MUX_s_1_2_2(nand_253_nl, or_3137_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1923_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_1078_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign or_2257_nl = (PEManager_15U_GetInputAddr_acc_tmp!=8'b00011010) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse);
  assign or_2253_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00011010);
  assign mux_794_nl = MUX_s_1_2_2(or_2257_nl, or_2253_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1497_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_794_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nand_205_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01111100))) &
      mux_773_cse);
  assign or_2863_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01111100);
  assign mux_990_nl = MUX_s_1_2_2(nand_205_nl, or_2863_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1791_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_990_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign or_2381_nl = (PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b0010110) | mux_799_cse;
  assign or_2374_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00101101);
  assign mux_832_nl = MUX_s_1_2_2(or_2381_nl, or_2374_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1554_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_832_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign or_2659_nl = (PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b0101100) | mux_799_cse;
  assign or_2652_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01011001);
  assign mux_920_nl = MUX_s_1_2_2(or_2659_nl, or_2652_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1686_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_920_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign or_2567_nl = (PEManager_15U_GetInputAddr_acc_tmp!=8'b01001011) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse);
  assign or_2563_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b010010)
      | nand_407_cse;
  assign mux_892_nl = MUX_s_1_2_2(or_2567_nl, or_2563_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1644_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_892_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1409_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10100011) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1410_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b101000)
      | nand_407_cse);
  assign mux_1068_nl = MUX_s_1_2_2(nor_1409_nl, nor_1410_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1908_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1068_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_132_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00111101))) &
      mux_773_cse);
  assign or_2477_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00111101);
  assign mux_864_nl = MUX_s_1_2_2(nand_132_nl, or_2477_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1602_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_864_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign or_2175_nl = (PEManager_15U_GetInputAddr_acc_tmp!=8'b00001101) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse);
  assign or_2171_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00001101);
  assign mux_768_nl = MUX_s_1_2_2(or_2175_nl, or_2171_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1458_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_768_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nand_133_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00111110))) &
      mux_773_cse);
  assign or_2482_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00111110);
  assign mux_866_nl = MUX_s_1_2_2(nand_133_nl, or_2482_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1605_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_866_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign and_2284_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00100000))) & mux_773_cse;
  assign nor_1045_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00100000));
  assign mux_806_nl = MUX_s_1_2_2(and_2284_nl, nor_1045_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1515_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_806_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nor_979_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00000110) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_980_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00000110));
  assign mux_754_nl = MUX_s_1_2_2(nor_979_nl, nor_980_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1437_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_754_nl & and_dcpl_759
      & PECoreRun_wen;
  assign and_2490_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11010010))) & mux_773_cse;
  assign nor_1543_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11010010));
  assign mux_1162_nl = MUX_s_1_2_2(and_2490_nl, nor_1543_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2049_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1162_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_102_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00011111))) &
      mux_773_cse);
  assign or_2287_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:5]!=3'b000)
      | nand_414_cse;
  assign mux_804_nl = MUX_s_1_2_2(nand_102_nl, or_2287_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1512_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_804_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign and_2376_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01110110))) & mux_773_cse;
  assign nor_1283_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01110110));
  assign mux_978_nl = MUX_s_1_2_2(and_2376_nl, nor_1283_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1773_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_978_nl & and_dcpl_759
      & PECoreRun_wen;
  assign and_2527_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11100110))) & mux_773_cse;
  assign nor_1602_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11100110));
  assign mux_1202_nl = MUX_s_1_2_2(and_2527_nl, nor_1602_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2109_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1202_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_366_nl = ~((PEManager_15U_GetInputAddr_acc_tmp==8'b11111010) & mux_773_cse);
  assign nand_502_nl = ~(input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4==8'b11111010));
  assign mux_1242_nl = MUX_s_1_2_2(nand_366_nl, nand_502_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2169_tmp = (~((reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_return_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) | mux_1242_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nand_318_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11011001))) &
      mux_773_cse);
  assign or_3430_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11011001);
  assign mux_1176_nl = MUX_s_1_2_2(nand_318_nl, or_3430_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2070_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_1176_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nand_369_nl = ~((PEManager_15U_GetInputAddr_acc_tmp==8'b11111101) & mux_773_cse);
  assign nand_507_nl = ~(input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4==8'b11111101));
  assign mux_1248_nl = MUX_s_1_2_2(nand_369_nl, nand_507_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2178_tmp = (~((reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_return_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) | mux_1248_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign and_2495_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11010100))) & mux_773_cse;
  assign nor_1549_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11010100));
  assign mux_1166_nl = MUX_s_1_2_2(and_2495_nl, nor_1549_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2055_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1166_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1324_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10000100) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1325_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10000100));
  assign mux_1006_nl = MUX_s_1_2_2(nor_1324_nl, nor_1325_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1815_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1006_nl & and_dcpl_759
      & PECoreRun_wen;
  assign or_2366_nl = (PEManager_15U_GetInputAddr_acc_tmp!=8'b00101011) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse);
  assign or_2362_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b001010)
      | nand_407_cse;
  assign mux_828_nl = MUX_s_1_2_2(or_2366_nl, or_2362_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1548_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_828_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign and_2423_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10100000))) & mux_773_cse;
  assign nor_1401_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10100000));
  assign mux_1062_nl = MUX_s_1_2_2(and_2423_nl, nor_1401_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1899_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1062_nl & and_dcpl_759
      & PECoreRun_wen;
  assign or_2359_nl = (PEManager_15U_GetInputAddr_acc_tmp!=8'b00101010) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse);
  assign or_2355_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00101010);
  assign mux_826_nl = MUX_s_1_2_2(or_2359_nl, or_2355_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1545_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_826_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1189_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b0101010) |
      mux_799_cse);
  assign nor_1190_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01010101));
  assign mux_912_nl = MUX_s_1_2_2(nor_1189_nl, nor_1190_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1674_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_912_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nor_973_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00000100) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_974_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00000100));
  assign mux_750_nl = MUX_s_1_2_2(nor_973_nl, nor_974_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1431_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_750_nl & and_dcpl_759
      & PECoreRun_wen;
  assign and_2271_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00010000))) & mux_773_cse;
  assign nor_1002_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00010000));
  assign mux_774_nl = MUX_s_1_2_2(and_2271_nl, nor_1002_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1467_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_774_nl & and_dcpl_759
      & PECoreRun_wen;
  assign or_2251_nl = (PEManager_15U_GetInputAddr_acc_tmp!=8'b00011001) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse);
  assign or_2247_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00011001);
  assign mux_792_nl = MUX_s_1_2_2(or_2251_nl, or_2247_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1494_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_792_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nand_114_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00101110))) &
      mux_773_cse);
  assign or_2383_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00101110);
  assign mux_834_nl = MUX_s_1_2_2(nand_114_nl, or_2383_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1557_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_834_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1093_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00110010) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1094_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00110010));
  assign mux_842_nl = MUX_s_1_2_2(nor_1093_nl, nor_1094_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1569_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_842_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_112_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00101000))) &
      mux_773_cse);
  assign or_2343_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00101000);
  assign mux_822_nl = MUX_s_1_2_2(nand_112_nl, or_2343_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1539_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_822_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign and_2374_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01110101))) & mux_773_cse;
  assign nor_1280_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01110101));
  assign mux_976_nl = MUX_s_1_2_2(and_2374_nl, nor_1280_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1770_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_976_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1330_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10000110) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1331_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10000110));
  assign mux_1010_nl = MUX_s_1_2_2(nor_1330_nl, nor_1331_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1821_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1010_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_236_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10011011))) &
      mux_773_cse);
  assign or_3059_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b100110)
      | nand_407_cse;
  assign mux_1052_nl = MUX_s_1_2_2(nand_236_nl, or_3059_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1884_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_1052_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nand_370_nl = ~((PEManager_15U_GetInputAddr_acc_tmp==8'b11111110) & mux_773_cse);
  assign nand_508_nl = ~(input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4==8'b11111110));
  assign mux_1250_nl = MUX_s_1_2_2(nand_370_nl, nand_508_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2181_tmp = (~((reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_return_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) | mux_1250_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1004_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00010001) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1005_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00010001));
  assign mux_776_nl = MUX_s_1_2_2(nor_1004_nl, nor_1005_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1470_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_776_nl & and_dcpl_759
      & PECoreRun_wen;
  assign and_2487_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11010000))) & mux_773_cse;
  assign nor_1538_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11010000));
  assign mux_1158_nl = MUX_s_1_2_2(and_2487_nl, nor_1538_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2043_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1158_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_276_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10111001))) &
      mux_773_cse);
  assign or_3239_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10111001);
  assign mux_1112_nl = MUX_s_1_2_2(nand_276_nl, or_3239_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1974_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_1112_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nand_320_nl = ~((PEManager_15U_GetInputAddr_acc_tmp==8'b11011011) & mux_773_cse);
  assign or_3441_nl = (~(input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]==6'b110110)))
      | nand_407_cse;
  assign mux_1180_nl = MUX_s_1_2_2(nand_320_nl, or_3441_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2076_tmp = (~((reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_return_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) | mux_1180_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nand_206_nl = ~((PEManager_15U_GetInputAddr_acc_tmp==8'b01111101) & mux_773_cse);
  assign nand_441_nl = ~(input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4==8'b01111101));
  assign mux_992_nl = MUX_s_1_2_2(nand_206_nl, nand_441_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1794_tmp = (~((reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_return_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) | mux_992_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1144_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01000100) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1145_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01000100));
  assign mux_878_nl = MUX_s_1_2_2(nor_1144_nl, nor_1145_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1623_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_878_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_99_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00011000))) &
      mux_773_cse);
  assign or_2241_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00011000);
  assign mux_790_nl = MUX_s_1_2_2(nand_99_nl, or_2241_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1491_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_790_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign or_2168_nl = (PEManager_15U_GetInputAddr_acc_tmp!=8'b00001100) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse);
  assign or_2164_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00001100);
  assign mux_766_nl = MUX_s_1_2_2(or_2168_nl, or_2164_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1455_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_766_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nand_130_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00111011))) &
      mux_773_cse);
  assign or_2466_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b001110)
      | nand_407_cse;
  assign mux_860_nl = MUX_s_1_2_2(nand_130_nl, or_2466_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1596_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_860_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign and_2481_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11000111))) & mux_773_cse;
  assign nor_1513_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:3]!=5'b11000)
      | nand_408_cse);
  assign mux_1140_nl = MUX_s_1_2_2(and_2481_nl, nor_1513_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2016_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1140_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_237_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10011100))) &
      mux_773_cse);
  assign or_3064_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10011100);
  assign mux_1054_nl = MUX_s_1_2_2(nand_237_nl, or_3064_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1887_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_1054_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign or_2582_nl = (PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b0100110) | mux_799_cse;
  assign or_2575_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01001101);
  assign mux_896_nl = MUX_s_1_2_2(or_2582_nl, or_2575_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1650_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_896_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nand_317_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11011000))) &
      mux_773_cse);
  assign or_3424_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11011000);
  assign mux_1174_nl = MUX_s_1_2_2(nand_317_nl, or_3424_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2067_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_1174_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1050_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00100010) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1051_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00100010));
  assign mux_810_nl = MUX_s_1_2_2(nor_1050_nl, nor_1051_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1521_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_810_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_367_nl = ~((PEManager_15U_GetInputAddr_acc_tmp==8'b11111011) & mux_773_cse);
  assign or_3621_nl = (~(input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]==6'b111110)))
      | nand_407_cse;
  assign mux_1244_nl = MUX_s_1_2_2(nand_367_nl, or_3621_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2172_tmp = (~((reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_return_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) | mux_1244_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign and_2523_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11100100))) & mux_773_cse;
  assign nor_1596_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11100100));
  assign mux_1198_nl = MUX_s_1_2_2(and_2523_nl, nor_1596_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2103_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1198_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_146_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01001110))) &
      mux_773_cse);
  assign or_2584_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01001110);
  assign mux_898_nl = MUX_s_1_2_2(nand_146_nl, or_2584_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1653_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_898_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1141_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01000011) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1142_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b010000)
      | nand_407_cse);
  assign mux_876_nl = MUX_s_1_2_2(nor_1141_nl, nor_1142_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1620_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_876_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1010_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00010011) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1011_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b000100)
      | nand_407_cse);
  assign mux_780_nl = MUX_s_1_2_2(nor_1010_nl, nor_1011_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1476_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_780_nl & and_dcpl_759
      & PECoreRun_wen;
  assign or_2264_nl = (PEManager_15U_GetInputAddr_acc_tmp!=8'b00011011) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse);
  assign or_2260_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b000110)
      | nand_407_cse;
  assign mux_796_nl = MUX_s_1_2_2(or_2264_nl, or_2260_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1500_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_796_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1178_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01010001) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1179_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01010001));
  assign mux_904_nl = MUX_s_1_2_2(nor_1178_nl, nor_1179_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1662_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_904_nl & and_dcpl_759
      & PECoreRun_wen;
  assign and_2429_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10100100))) & mux_773_cse;
  assign nor_1413_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10100100));
  assign mux_1070_nl = MUX_s_1_2_2(and_2429_nl, nor_1413_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1911_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1070_nl & and_dcpl_759
      & PECoreRun_wen;
  assign and_2457_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b10110111) & mux_773_cse;
  assign nor_1466_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:3]!=5'b10110)
      | nand_408_cse);
  assign mux_1108_nl = MUX_s_1_2_2(and_2457_nl, nor_1466_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1968_tmp = (~(reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_return_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) & mux_1108_nl & and_dcpl_759
      & PECoreRun_wen;
  assign and_2447_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10110011))) & mux_773_cse;
  assign nor_1454_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b101100)
      | nand_407_cse);
  assign mux_1100_nl = MUX_s_1_2_2(and_2447_nl, nor_1454_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1956_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1100_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_280_nl = ~((PEManager_15U_GetInputAddr_acc_tmp==8'b10111101) & mux_773_cse);
  assign nand_462_nl = ~(input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4==8'b10111101));
  assign mux_1120_nl = MUX_s_1_2_2(nand_280_nl, nand_462_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1986_tmp = (~((reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_return_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) | mux_1120_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign and_2497_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11010101))) & mux_773_cse;
  assign nor_1552_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11010101));
  assign mux_1168_nl = MUX_s_1_2_2(and_2497_nl, nor_1552_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2058_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1168_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_342_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11101010))) &
      mux_773_cse);
  assign or_3527_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11101010);
  assign mux_1210_nl = MUX_s_1_2_2(nand_342_nl, or_3527_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2121_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_1210_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nand_364_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11111000))) &
      mux_773_cse);
  assign or_3604_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11111000);
  assign mux_1238_nl = MUX_s_1_2_2(nand_364_nl, or_3604_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2163_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_1238_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nand_365_nl = ~((PEManager_15U_GetInputAddr_acc_tmp==8'b11111001) & mux_773_cse);
  assign nand_501_nl = ~(input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4==8'b11111001));
  assign mux_1240_nl = MUX_s_1_2_2(nand_365_nl, nand_501_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2166_tmp = (~((reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_return_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) | mux_1240_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign and_2364_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01110000))) & mux_773_cse;
  assign nor_1266_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01110000));
  assign mux_966_nl = MUX_s_1_2_2(and_2364_nl, nor_1266_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1755_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_966_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_340_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11101000))) &
      mux_773_cse);
  assign or_3516_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11101000);
  assign mux_1206_nl = MUX_s_1_2_2(nand_340_nl, or_3516_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2115_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_1206_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign and_2451_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10110101))) & mux_773_cse;
  assign nor_1460_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10110101));
  assign mux_1104_nl = MUX_s_1_2_2(and_2451_nl, nor_1460_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1962_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1104_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1007_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00010010) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1008_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00010010));
  assign mux_778_nl = MUX_s_1_2_2(nor_1007_nl, nor_1008_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1473_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_778_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_319_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11011010))) &
      mux_773_cse);
  assign or_3435_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11011010);
  assign mux_1178_nl = MUX_s_1_2_2(nand_319_nl, or_3435_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2073_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_1178_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign and_2328_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01010000))) & mux_773_cse;
  assign nor_1176_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01010000));
  assign mux_902_nl = MUX_s_1_2_2(and_2328_nl, nor_1176_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1659_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_902_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_202_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01111001))) &
      mux_773_cse);
  assign or_2847_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01111001);
  assign mux_984_nl = MUX_s_1_2_2(nand_202_nl, or_2847_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1782_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_984_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign or_2188_nl = (PEManager_15U_GetInputAddr_acc_tmp!=8'b00001111) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse);
  assign or_2184_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:4]!=4'b0000)
      | nand_410_cse;
  assign mux_772_nl = MUX_s_1_2_2(or_2188_nl, or_2184_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1464_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_772_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nand_163_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01011100))) &
      mux_773_cse);
  assign or_2672_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01011100);
  assign mux_926_nl = MUX_s_1_2_2(nand_163_nl, or_2672_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1695_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_926_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nand_234_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10011000))) &
      mux_773_cse);
  assign or_3038_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10011000);
  assign mux_1046_nl = MUX_s_1_2_2(nand_234_nl, or_3038_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1875_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_1046_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nand_297_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11001011))) &
      mux_773_cse);
  assign or_3349_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b110010)
      | nand_407_cse;
  assign mux_1148_nl = MUX_s_1_2_2(nand_297_nl, or_3349_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2028_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_1148_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign or_2090_nl = (state_2_1_sva[0]) | (~ input_port_PopNB_mioi_return_rsc_z_mxwt)
      | PECore_RunFSM_switch_lp_nor_tmp_1;
  assign or_2089_nl = (~ PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva)
      | PECore_RunFSM_switch_lp_nor_tmp_1;
  assign mux_741_nl = MUX_s_1_2_2(or_2090_nl, or_2089_nl, or_2088_cse);
  assign nor_961_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00000000) | mux_741_nl);
  assign nor_962_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00000000));
  assign mux_742_nl = MUX_s_1_2_2(nor_961_nl, nor_962_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1419_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_742_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_113_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00101100))) &
      mux_773_cse);
  assign or_2368_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00101100);
  assign mux_830_nl = MUX_s_1_2_2(nand_113_nl, or_2368_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1551_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_830_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nand_345_nl = ~((PEManager_15U_GetInputAddr_acc_tmp==8'b11101101) & mux_773_cse);
  assign nand_485_nl = ~(input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4==8'b11101101));
  assign mux_1216_nl = MUX_s_1_2_2(nand_345_nl, nand_485_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2130_tmp = (~((reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_return_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) | mux_1216_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign or_2758_nl = (PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b0110100) | mux_799_cse;
  assign or_2751_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01101001);
  assign mux_952_nl = MUX_s_1_2_2(or_2758_nl, or_2751_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1734_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_952_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign and_2334_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01010100))) & mux_773_cse;
  assign nor_1188_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01010100));
  assign mux_910_nl = MUX_s_1_2_2(and_2334_nl, nor_1188_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1671_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_910_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1495_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11000001) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1496_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11000001));
  assign mux_1128_nl = MUX_s_1_2_2(nor_1495_nl, nor_1496_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1998_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1128_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1586_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b1110000) |
      mux_799_cse);
  assign nor_1587_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11100001));
  assign mux_1192_nl = MUX_s_1_2_2(nor_1586_nl, nor_1587_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2094_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1192_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1016_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00010101) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1017_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00010101));
  assign mux_784_nl = MUX_s_1_2_2(nor_1016_nl, nor_1017_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1482_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_784_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_221_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10001111))) &
      mux_773_cse);
  assign or_2982_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:4]!=4'b1000)
      | nand_410_cse;
  assign mux_1028_nl = MUX_s_1_2_2(nand_221_nl, or_2982_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1848_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_1028_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign or_2458_nl = (PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b0011100) | mux_799_cse;
  assign or_2451_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00111001);
  assign mux_856_nl = MUX_s_1_2_2(or_2458_nl, or_2451_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1590_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_856_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nand_235_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10011010))) &
      mux_773_cse);
  assign or_3053_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10011010);
  assign mux_1050_nl = MUX_s_1_2_2(nand_235_nl, or_3053_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1881_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_1050_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nand_134_nl = ~((PEManager_15U_GetInputAddr_acc_tmp==8'b00111111) & mux_773_cse);
  assign or_2488_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:6]!=2'b00)
      | nand_422_cse;
  assign mux_868_nl = MUX_s_1_2_2(nand_134_nl, or_2488_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1608_tmp = (~((reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_return_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) | mux_868_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nand_180_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01101010))) &
      mux_773_cse);
  assign or_2760_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01101010);
  assign mux_954_nl = MUX_s_1_2_2(nand_180_nl, or_2760_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1737_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_954_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign and_2340_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01010111))) & mux_773_cse;
  assign nor_1196_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:3]!=5'b01010)
      | nand_408_cse);
  assign mux_916_nl = MUX_s_1_2_2(and_2340_nl, nor_1196_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1680_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_916_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1447_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b1011000) |
      mux_799_cse);
  assign nor_1448_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10110001));
  assign mux_1096_nl = MUX_s_1_2_2(nor_1447_nl, nor_1448_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1950_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1096_nl & and_dcpl_759
      & PECoreRun_wen;
  assign or_3341_nl = (PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b1100100) | mux_799_cse;
  assign or_3334_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11001001);
  assign mux_1144_nl = MUX_s_1_2_2(or_3341_nl, or_3334_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2022_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_1144_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nand_203_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01111010))) &
      mux_773_cse);
  assign or_2852_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01111010);
  assign mux_986_nl = MUX_s_1_2_2(nand_203_nl, or_2852_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1785_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_986_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1267_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b0111000) |
      mux_799_cse);
  assign nor_1268_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01110001));
  assign mux_968_nl = MUX_s_1_2_2(nor_1267_nl, nor_1268_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1758_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_968_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_160_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01011000))) &
      mux_773_cse);
  assign or_2646_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01011000);
  assign mux_918_nl = MUX_s_1_2_2(nand_160_nl, or_2646_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1683_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_918_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign or_2560_nl = (PEManager_15U_GetInputAddr_acc_tmp!=8'b01001010) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse);
  assign or_2556_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01001010);
  assign mux_890_nl = MUX_s_1_2_2(or_2560_nl, or_2556_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1641_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_890_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nand_161_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01011010))) &
      mux_773_cse);
  assign or_2661_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01011010);
  assign mux_922_nl = MUX_s_1_2_2(nand_161_nl, or_2661_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1689_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_922_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign or_2353_nl = (PEManager_15U_GetInputAddr_acc_tmp!=8'b00101001) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse);
  assign or_2349_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00101001);
  assign mux_824_nl = MUX_s_1_2_2(or_2353_nl, or_2349_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1542_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_824_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nor_982_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00000111) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_983_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:3]!=5'b00000)
      | nand_408_cse);
  assign mux_756_nl = MUX_s_1_2_2(nor_982_nl, nor_983_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1440_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_756_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_343_nl = ~((PEManager_15U_GetInputAddr_acc_tmp==8'b11101011) & mux_773_cse);
  assign or_3533_nl = (~(input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]==6'b111010)))
      | nand_407_cse;
  assign mux_1212_nl = MUX_s_1_2_2(nand_343_nl, or_3533_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2124_tmp = (~((reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_return_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) | mux_1212_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nand_207_nl = ~((PEManager_15U_GetInputAddr_acc_tmp==8'b01111110) & mux_773_cse);
  assign nand_442_nl = ~(input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4==8'b01111110));
  assign mux_994_nl = MUX_s_1_2_2(nand_207_nl, nand_442_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1797_tmp = (~((reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_return_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) | mux_994_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1361_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10010010) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1362_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10010010));
  assign mux_1034_nl = MUX_s_1_2_2(nor_1361_nl, nor_1362_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1857_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1034_nl & and_dcpl_759
      & PECoreRun_wen;
  assign and_2525_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11100101))) & mux_773_cse;
  assign nor_1599_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11100101));
  assign mux_1200_nl = MUX_s_1_2_2(and_2525_nl, nor_1599_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2106_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1200_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_324_nl = ~((PEManager_15U_GetInputAddr_acc_tmp==8'b11011111) & mux_773_cse);
  assign or_3463_nl = (~(input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:5]==3'b110)))
      | nand_414_cse;
  assign mux_1188_nl = MUX_s_1_2_2(nand_324_nl, or_3463_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2088_tmp = (~((reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_return_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) | mux_1188_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1403_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10100001) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1404_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10100001));
  assign mux_1064_nl = MUX_s_1_2_2(nor_1403_nl, nor_1404_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1902_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1064_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_300_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11001110))) &
      mux_773_cse);
  assign or_3365_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11001110);
  assign mux_1154_nl = MUX_s_1_2_2(nand_300_nl, or_3365_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2037_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_1154_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1318_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10000010) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1319_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10000010));
  assign mux_1002_nl = MUX_s_1_2_2(nor_1318_nl, nor_1319_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1809_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1002_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1501_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11000011) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1502_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b110000)
      | nand_407_cse);
  assign mux_1132_nl = MUX_s_1_2_2(nor_1501_nl, nor_1502_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2004_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1132_nl & and_dcpl_759
      & PECoreRun_wen;
  assign input_mem_banks_read_read_data_and_21_tmp = PECoreRun_wen & and_dcpl_219;
  assign and_2358_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01100111))) & mux_773_cse;
  assign nor_1241_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:3]!=5'b01100)
      | nand_408_cse);
  assign mux_948_nl = MUX_s_1_2_2(and_2358_nl, nor_1241_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1728_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_948_nl & and_dcpl_759
      & PECoreRun_wen;
  assign and_2352_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01100100))) & mux_773_cse;
  assign nor_1233_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01100100));
  assign mux_942_nl = MUX_s_1_2_2(and_2352_nl, nor_1233_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1719_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_942_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_238_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10011101))) &
      mux_773_cse);
  assign or_3070_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10011101);
  assign mux_1056_nl = MUX_s_1_2_2(nand_238_nl, or_3070_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1890_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_1056_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nand_208_nl = ~((PEManager_15U_GetInputAddr_acc_tmp==8'b01111111) & mux_773_cse);
  assign or_2880_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01111111);
  assign mux_996_nl = MUX_s_1_2_2(nand_208_nl, or_2880_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1800_tmp = (~((reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_return_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) | mux_996_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1090_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00110001) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1091_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00110001));
  assign mux_840_nl = MUX_s_1_2_2(nor_1090_nl, nor_1091_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1566_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_840_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_115_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00101111))) &
      mux_773_cse);
  assign or_2389_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:4]!=4'b0010)
      | nand_410_cse;
  assign mux_836_nl = MUX_s_1_2_2(nand_115_nl, or_2389_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1560_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_836_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign and_2543_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11110000))) & mux_773_cse;
  assign nor_1632_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11110000));
  assign mux_1222_nl = MUX_s_1_2_2(and_2543_nl, nor_1632_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2139_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1222_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_323_nl = ~((PEManager_15U_GetInputAddr_acc_tmp==8'b11011110) & mux_773_cse);
  assign nand_476_nl = ~(input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4==8'b11011110));
  assign mux_1186_nl = MUX_s_1_2_2(nand_323_nl, nand_476_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2085_tmp = (~((reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_return_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) | mux_1186_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nand_201_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01111000))) &
      mux_773_cse);
  assign or_2841_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01111000);
  assign mux_982_nl = MUX_s_1_2_2(nand_201_nl, or_2841_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1779_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_982_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1138_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01000010) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1139_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01000010));
  assign mux_874_nl = MUX_s_1_2_2(nor_1138_nl, nor_1139_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1617_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_874_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1053_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00100011) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1054_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b001000)
      | nand_407_cse);
  assign mux_812_nl = MUX_s_1_2_2(nor_1053_nl, nor_1054_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1524_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_812_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1327_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10000101) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1328_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10000101));
  assign mux_1008_nl = MUX_s_1_2_2(nor_1327_nl, nor_1328_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1818_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1008_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_256_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10101100))) &
      mux_773_cse);
  assign or_3163_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10101100);
  assign mux_1086_nl = MUX_s_1_2_2(nand_256_nl, or_3163_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1935_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_1086_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1147_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01000101) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1148_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01000101));
  assign mux_880_nl = MUX_s_1_2_2(nor_1147_nl, nor_1148_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1626_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_880_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_182_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01101100))) &
      mux_773_cse);
  assign or_2771_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01101100);
  assign mux_958_nl = MUX_s_1_2_2(nand_182_nl, or_2771_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1743_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_958_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign or_2181_nl = (PEManager_15U_GetInputAddr_acc_tmp!=8'b00001110) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse);
  assign or_2177_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00001110);
  assign mux_770_nl = MUX_s_1_2_2(or_2181_nl, or_2177_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1461_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_770_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nand_240_nl = ~((PEManager_15U_GetInputAddr_acc_tmp==8'b10011111) & mux_773_cse);
  assign or_3081_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:5]!=3'b100)
      | nand_414_cse;
  assign mux_1060_nl = MUX_s_1_2_2(nand_240_nl, or_3081_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1896_tmp = (~((reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_return_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) | mux_1060_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nand_145_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01001100))) &
      mux_773_cse);
  assign or_2569_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01001100);
  assign mux_894_nl = MUX_s_1_2_2(nand_145_nl, or_2569_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1647_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_894_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign and_2545_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11110001))) & mux_773_cse;
  assign nor_1635_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11110001));
  assign mux_1224_nl = MUX_s_1_2_2(and_2545_nl, nor_1635_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2142_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1224_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_255_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10101011))) &
      mux_773_cse);
  assign or_3158_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b101010)
      | nand_407_cse;
  assign mux_1084_nl = MUX_s_1_2_2(nand_255_nl, or_3158_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1932_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_1084_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nand_295_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11001000))) &
      mux_773_cse);
  assign or_3328_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11001000);
  assign mux_1142_nl = MUX_s_1_2_2(nand_295_nl, or_3328_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2019_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_1142_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1226_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01100010) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1227_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01100010));
  assign mux_938_nl = MUX_s_1_2_2(nor_1226_nl, nor_1227_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1713_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_938_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_341_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11101001))) &
      mux_773_cse);
  assign or_3522_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11101001);
  assign mux_1208_nl = MUX_s_1_2_2(nand_341_nl, or_3522_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2118_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_1208_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign and_2411_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10010100))) & mux_773_cse;
  assign nor_1368_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10010100));
  assign mux_1038_nl = MUX_s_1_2_2(and_2411_nl, nor_1368_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1863_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1038_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_179_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01101000))) &
      mux_773_cse);
  assign or_2745_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01101000);
  assign mux_950_nl = MUX_s_1_2_2(nand_179_nl, or_2745_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1731_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_950_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign and_2309_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00110111))) & mux_773_cse;
  assign nor_1108_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:3]!=5'b00110)
      | nand_408_cse);
  assign mux_852_nl = MUX_s_1_2_2(and_2309_nl, nor_1108_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1584_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_852_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_204_nl = ~((PEManager_15U_GetInputAddr_acc_tmp==8'b01111011) & mux_773_cse);
  assign or_2858_nl = (~(input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]==6'b011110)))
      | nand_407_cse;
  assign mux_988_nl = MUX_s_1_2_2(nand_204_nl, or_2858_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1788_tmp = (~((reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_return_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) | mux_988_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign and_2380_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b01110111) & mux_773_cse;
  assign nor_1286_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:3]!=5'b01110)
      | nand_408_cse);
  assign mux_980_nl = MUX_s_1_2_2(and_2380_nl, nor_1286_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1776_tmp = (~(reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_return_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) & mux_980_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1333_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10000111) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1334_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:3]!=5'b10000)
      | nand_408_cse);
  assign mux_1012_nl = MUX_s_1_2_2(nor_1333_nl, nor_1334_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1824_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1012_nl & and_dcpl_759
      & PECoreRun_wen;
  assign and_2372_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01110100))) & mux_773_cse;
  assign nor_1277_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01110100));
  assign mux_974_nl = MUX_s_1_2_2(and_2372_nl, nor_1277_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1767_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_974_nl & and_dcpl_759
      & PECoreRun_wen;
  assign and_2392_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10000000))) & mux_773_cse;
  assign nor_1313_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10000000));
  assign mux_998_nl = MUX_s_1_2_2(and_2392_nl, nor_1313_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1803_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_998_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1498_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11000010) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1499_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11000010));
  assign mux_1130_nl = MUX_s_1_2_2(nor_1498_nl, nor_1499_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2001_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1130_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_101_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00011110))) &
      mux_773_cse);
  assign or_2281_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00011110);
  assign mux_802_nl = MUX_s_1_2_2(nand_101_nl, or_2281_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1509_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_802_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nand_218_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10001000))) &
      mux_773_cse);
  assign or_2936_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10001000);
  assign mux_1014_nl = MUX_s_1_2_2(nand_218_nl, or_2936_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1827_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_1014_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign and_2581_nl = (~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3]))) & mux_tmp_1225;
  assign nand_511_nl = ~(reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_return_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:18]==2'b01));
  assign mux_1253_nl = MUX_s_1_2_2(and_2581_nl, mux_tmp_1225, nand_511_nl);
  assign and_2184_tmp = mux_1253_nl & and_dcpl_759 & PECoreRun_wen;
  assign nand_322_nl = ~((PEManager_15U_GetInputAddr_acc_tmp==8'b11011101) & mux_773_cse);
  assign nand_475_nl = ~(input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4==8'b11011101));
  assign mux_1184_nl = MUX_s_1_2_2(nand_322_nl, nand_475_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2082_tmp = (~((reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_return_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) | mux_1184_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign and_2553_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11110100))) & mux_773_cse;
  assign nor_1644_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11110100));
  assign mux_1230_nl = MUX_s_1_2_2(and_2553_nl, nor_1644_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2151_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1230_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_100_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00011100))) &
      mux_773_cse);
  assign or_2266_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00011100);
  assign mux_798_nl = MUX_s_1_2_2(nand_100_nl, or_2266_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1503_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_798_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign and_2531_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b11100111) & mux_773_cse;
  assign nor_1605_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:3]!=5'b11100)
      | nand_408_cse);
  assign mux_1204_nl = MUX_s_1_2_2(and_2531_nl, nor_1605_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2112_tmp = (~(reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_return_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) & mux_1204_nl & and_dcpl_759
      & PECoreRun_wen;
  assign and_2449_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10110100))) & mux_773_cse;
  assign nor_1457_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10110100));
  assign mux_1102_nl = MUX_s_1_2_2(and_2449_nl, nor_1457_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1959_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1102_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1358_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10010001) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1359_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10010001));
  assign mux_1032_nl = MUX_s_1_2_2(nor_1358_nl, nor_1359_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1854_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1032_nl & and_dcpl_759
      & PECoreRun_wen;
  assign and_2414_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10010110))) & mux_773_cse;
  assign nor_1373_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10010110));
  assign mux_1042_nl = MUX_s_1_2_2(and_2414_nl, nor_1373_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1869_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1042_nl & and_dcpl_759
      & PECoreRun_wen;
  assign and_2346_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01100000))) & mux_773_cse;
  assign nor_1221_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01100000));
  assign mux_934_nl = MUX_s_1_2_2(and_2346_nl, nor_1221_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1707_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_934_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_219_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10001100))) &
      mux_773_cse);
  assign or_2961_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10001100);
  assign mux_1022_nl = MUX_s_1_2_2(nand_219_nl, or_2961_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1839_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_1022_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign or_2142_nl = (PEManager_15U_GetInputAddr_acc_tmp!=8'b00001000) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse);
  assign or_2138_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00001000);
  assign mux_758_nl = MUX_s_1_2_2(or_2142_nl, or_2138_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1443_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_758_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nand_162_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01011011))) &
      mux_773_cse);
  assign or_2667_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b010110)
      | nand_407_cse;
  assign mux_924_nl = MUX_s_1_2_2(nand_162_nl, or_2667_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1692_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_924_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nand_296_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11001010))) &
      mux_773_cse);
  assign or_3343_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11001010);
  assign mux_1146_nl = MUX_s_1_2_2(nand_296_nl, or_3343_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2025_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_1146_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1013_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00010100) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1014_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00010100));
  assign mux_782_nl = MUX_s_1_2_2(nor_1013_nl, nor_1014_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1479_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_782_nl & and_dcpl_759
      & PECoreRun_wen;
  assign or_3150_nl = (PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b1010100) | mux_799_cse;
  assign or_3143_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10101001);
  assign mux_1080_nl = MUX_s_1_2_2(or_3150_nl, or_3143_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1926_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_1080_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign and_2441_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10110000))) & mux_773_cse;
  assign nor_1446_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10110000));
  assign mux_1094_nl = MUX_s_1_2_2(and_2441_nl, nor_1446_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1947_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1094_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_239_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10011110))) &
      mux_773_cse);
  assign or_3075_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10011110);
  assign mux_1058_nl = MUX_s_1_2_2(nand_239_nl, or_3075_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1893_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_1058_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1369_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b1001010) |
      mux_799_cse);
  assign nor_1370_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10010101));
  assign mux_1040_nl = MUX_s_1_2_2(nor_1369_nl, nor_1370_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1866_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1040_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1364_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10010011) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1365_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b100100)
      | nand_407_cse);
  assign mux_1036_nl = MUX_s_1_2_2(nor_1364_nl, nor_1365_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1860_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1036_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1101_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b0011010) |
      mux_799_cse);
  assign nor_1102_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00110101));
  assign mux_848_nl = MUX_s_1_2_2(nor_1101_nl, nor_1102_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1578_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_848_nl & and_dcpl_759
      & PECoreRun_wen;
  assign or_2279_nl = (PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b0001110) | mux_799_cse;
  assign or_2272_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00011101);
  assign mux_800_nl = MUX_s_1_2_2(or_2279_nl, or_2272_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1506_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_800_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign or_3051_nl = (PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b1001100) | mux_799_cse;
  assign or_3044_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10011001);
  assign mux_1048_nl = MUX_s_1_2_2(or_3051_nl, or_3044_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1878_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_1048_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nand_368_nl = ~((PEManager_15U_GetInputAddr_acc_tmp==8'b11111100) & mux_773_cse);
  assign nand_505_nl = ~(input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4==8'b11111100));
  assign mux_1246_nl = MUX_s_1_2_2(nand_368_nl, nand_505_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2175_tmp = (~((reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_return_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) | mux_1246_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nor_970_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00000011) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_971_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b000000)
      | nand_407_cse);
  assign mux_748_nl = MUX_s_1_2_2(nor_970_nl, nor_971_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1428_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_748_nl & and_dcpl_759
      & PECoreRun_wen;
  assign and_2355_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01100110))) & mux_773_cse;
  assign nor_1238_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01100110));
  assign mux_946_nl = MUX_s_1_2_2(and_2355_nl, nor_1238_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1725_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_946_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_181_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01101011))) &
      mux_773_cse);
  assign or_2766_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b011010)
      | nand_407_cse;
  assign mux_956_nl = MUX_s_1_2_2(nand_181_nl, or_2766_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1740_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_956_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign or_2149_nl = (PEManager_15U_GetInputAddr_acc_tmp!=8'b00001001) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse);
  assign or_2145_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00001001);
  assign mux_760_nl = MUX_s_1_2_2(or_2149_nl, or_2145_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1446_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_760_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign or_2946_nl = (PEManager_15U_GetInputAddr_acc_tmp!=8'b10001001) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse);
  assign or_2942_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10001001);
  assign mux_1016_nl = MUX_s_1_2_2(or_2946_nl, or_2942_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1830_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_1016_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign and_2370_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01110011))) & mux_773_cse;
  assign nor_1274_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b011100)
      | nand_407_cse);
  assign mux_972_nl = MUX_s_1_2_2(and_2370_nl, nor_1274_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1764_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_972_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_254_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10101010))) &
      mux_773_cse);
  assign or_3152_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10101010);
  assign mux_1082_nl = MUX_s_1_2_2(nand_254_nl, or_3152_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1929_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_1082_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign and_2493_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11010011))) & mux_773_cse;
  assign nor_1546_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:2]!=6'b110100)
      | nand_407_cse);
  assign mux_1164_nl = MUX_s_1_2_2(and_2493_nl, nor_1546_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2052_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1164_nl & and_dcpl_759
      & PECoreRun_wen;
  assign or_2155_nl = (PEManager_15U_GetInputAddr_acc_tmp!=8'b00001010) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse);
  assign or_2151_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00001010);
  assign mux_762_nl = MUX_s_1_2_2(or_2155_nl, or_2151_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1449_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_762_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1506_nl = ~((PEManager_15U_GetInputAddr_acc_tmp[7:1]!=7'b1100010) |
      mux_799_cse);
  assign nor_1507_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11000101));
  assign mux_1136_nl = MUX_s_1_2_2(nor_1506_nl, nor_1507_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2010_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1136_nl & and_dcpl_759
      & PECoreRun_wen;
  assign and_2315_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01000000))) & mux_773_cse;
  assign nor_1133_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01000000));
  assign mux_870_nl = MUX_s_1_2_2(and_2315_nl, nor_1133_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1611_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_870_nl & and_dcpl_759
      & PECoreRun_wen;
  assign and_2432_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10100110))) & mux_773_cse;
  assign nor_1418_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10100110));
  assign mux_1074_nl = MUX_s_1_2_2(and_2432_nl, nor_1418_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1917_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1074_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_282_nl = ~((PEManager_15U_GetInputAddr_acc_tmp==8'b10111111) & mux_773_cse);
  assign or_3272_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:6]!=2'b10)
      | nand_422_cse;
  assign mux_1124_nl = MUX_s_1_2_2(nand_282_nl, or_3272_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1992_tmp = (~((reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_return_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) | mux_1124_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign and_2478_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b11000110))) & mux_773_cse;
  assign nor_1510_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b11000110));
  assign mux_1138_nl = MUX_s_1_2_2(and_2478_nl, nor_1510_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2013_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1138_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_281_nl = ~((PEManager_15U_GetInputAddr_acc_tmp==8'b10111110) & mux_773_cse);
  assign nand_463_nl = ~(input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4==8'b10111110));
  assign mux_1122_nl = MUX_s_1_2_2(nand_281_nl, nand_463_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1989_tmp = (~((reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_return_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) | mux_1122_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nor_976_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00000101) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_977_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00000101));
  assign mux_752_nl = MUX_s_1_2_2(nor_976_nl, nor_977_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1434_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_752_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_275_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10111000))) &
      mux_773_cse);
  assign or_3233_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10111000);
  assign mux_1110_nl = MUX_s_1_2_2(nand_275_nl, or_3233_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1971_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_1110_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign and_2503_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b11010111) & mux_773_cse;
  assign nor_1558_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:3]!=5'b11010)
      | nand_408_cse);
  assign mux_1172_nl = MUX_s_1_2_2(and_2503_nl, nor_1558_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2064_tmp = (~(reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_return_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) & mux_1172_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1059_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00100101) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1060_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00100101));
  assign mux_816_nl = MUX_s_1_2_2(nor_1059_nl, nor_1060_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1530_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_816_nl & and_dcpl_759
      & PECoreRun_wen;
  assign and_2565_nl = (PEManager_15U_GetInputAddr_acc_tmp==8'b11110111) & mux_773_cse;
  assign nor_1651_nl = ~((~(input_write_req_valid_lpi_1_dfm_1_1 & (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:3]==5'b11110)))
      | nand_408_cse);
  assign mux_1236_nl = MUX_s_1_2_2(and_2565_nl, nor_1651_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_2160_tmp = (~(reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_return_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) & mux_1236_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1056_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00100100) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1057_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00100100));
  assign mux_814_nl = MUX_s_1_2_2(nor_1056_nl, nor_1057_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1527_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_814_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_220_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10001110))) &
      mux_773_cse);
  assign or_2976_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10001110);
  assign mux_1026_nl = MUX_s_1_2_2(nand_220_nl, or_2976_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1845_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_1026_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign and_2444_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10110010))) & mux_773_cse;
  assign nor_1451_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10110010));
  assign mux_1098_nl = MUX_s_1_2_2(and_2444_nl, nor_1451_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1953_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1098_nl & and_dcpl_759
      & PECoreRun_wen;
  assign or_2554_nl = (PEManager_15U_GetInputAddr_acc_tmp!=8'b01001001) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse);
  assign or_2550_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01001001);
  assign mux_888_nl = MUX_s_1_2_2(or_2554_nl, or_2550_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1638_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_888_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign and_2405_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b10010000))) & mux_773_cse;
  assign nor_1356_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b10010000));
  assign mux_1030_nl = MUX_s_1_2_2(and_2405_nl, nor_1356_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1851_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_1030_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1019_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00010110) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1020_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00010110));
  assign mux_786_nl = MUX_s_1_2_2(nor_1019_nl, nor_1020_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1485_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_786_nl & and_dcpl_759
      & PECoreRun_wen;
  assign and_2297_nl = (~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00110000))) & mux_773_cse;
  assign nor_1088_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00110000));
  assign mux_838_nl = MUX_s_1_2_2(and_2297_nl, nor_1088_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1563_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_838_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_128_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00111000))) &
      mux_773_cse);
  assign or_2445_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00111000);
  assign mux_854_nl = MUX_s_1_2_2(nand_128_nl, or_2445_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1587_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_854_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1065_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00100111) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1066_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:3]!=5'b00100)
      | nand_408_cse);
  assign mux_820_nl = MUX_s_1_2_2(nor_1065_nl, nor_1066_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1536_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_820_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_129_nl = ~((~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00111010))) &
      mux_773_cse);
  assign or_2460_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00111010);
  assign mux_858_nl = MUX_s_1_2_2(nand_129_nl, or_2460_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1593_tmp = (~((~((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]))
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])))) | mux_858_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nor_964_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b00000001) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_965_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b00000001));
  assign mux_744_nl = MUX_s_1_2_2(nor_964_nl, nor_965_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1422_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_744_nl & and_dcpl_759
      & PECoreRun_wen;
  assign nand_166_nl = ~((PEManager_15U_GetInputAddr_acc_tmp==8'b01011111) & mux_773_cse);
  assign or_2689_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4[7:5]!=3'b010)
      | nand_414_cse;
  assign mux_932_nl = MUX_s_1_2_2(nand_166_nl, or_2689_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1704_tmp = (~((reg_rva_in_PopNB_mioi_iswt0_cse & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_return_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]))
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]) & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) | mux_932_nl)) & and_dcpl_759
      & PECoreRun_wen;
  assign nor_1150_nl = ~((PEManager_15U_GetInputAddr_acc_tmp!=8'b01000110) | PECore_RunFSM_switch_lp_nor_tmp_1
      | (~ mux_743_cse));
  assign nor_1151_nl = ~((~ input_write_req_valid_lpi_1_dfm_1_1) | (while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4!=8'b01000110));
  assign mux_882_nl = MUX_s_1_2_2(nor_1150_nl, nor_1151_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign and_1629_tmp = ((~ reg_rva_in_PopNB_mioi_iswt0_cse) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3])) & mux_882_nl & and_dcpl_759
      & PECoreRun_wen;
  assign input_mem_banks_read_read_data_and_20_tmp = PECoreRun_wen & (~((~((~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2)
      & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_17_itm_1 & (~ rva_in_reg_rw_sva_st_1_4)))
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4))
      & while_stage_0_6;
  assign nor_927_nl = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt));
  assign or_1587_nl = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[15:1]!=15'b000000000000000);
  assign mux_529_nl = MUX_s_1_2_2(nor_927_nl, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt,
      or_1587_nl);
  assign or_1590_nl = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]) | (~((~ while_stage_0_3)
      | (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1)
      | PECore_DecodeAxiWrite_switch_lp_equal_tmp_1 | PECore_DecodeAxiWrite_switch_lp_equal_tmp_2
      | PECore_DecodeAxiWrite_switch_lp_nor_tmp_1 | (~(reg_rva_in_reg_rw_sva_st_1_1_cse
      & mux_529_nl))));
  assign mux_530_nl = MUX_s_1_2_2(rva_in_PopNB_mioi_data_rw_rsc_z_mxwt, or_1590_nl,
      nor_536_cse);
  assign and_1217_tmp = (~ mux_530_nl) & and_692_cse & PECoreRun_wen;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_cgo_ir_cse <=
          1'b0;
      reg_PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_cgo_ir_cse <=
          1'b0;
      reg_weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_cse <= 1'b0;
      reg_weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_cse <= 1'b0;
      reg_rva_out_Push_mioi_iswt0_cse <= 1'b0;
      reg_start_PopNB_mioi_iswt0_cse <= 1'b0;
      reg_act_port_Push_mioi_iswt0_cse <= 1'b0;
      reg_rva_in_PopNB_mioi_iswt0_cse <= 1'b0;
      pe_config_manager_counter_sva_dfm_3_1 <= 4'b0000;
      pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_nor_mdf_sva_st_1
          <= 1'b0;
      pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1
          <= 1'b0;
      while_stage_0_3 <= 1'b0;
      while_stage_0_4 <= 1'b0;
      while_stage_0_5 <= 1'b0;
      while_stage_0_6 <= 1'b0;
      while_stage_0_7 <= 1'b0;
      while_stage_0_8 <= 1'b0;
      while_stage_0_9 <= 1'b0;
      while_stage_0_10 <= 1'b0;
      while_stage_0_11 <= 1'b0;
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_122_itm_1 <= 1'b0;
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_95_itm_1 <= 1'b0;
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_93_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_1_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_1
          <= 1'b0;
      input_read_addrs_sva_1_1 <= 8'b00000000;
      ProductSum_for_asn_64_itm_1 <= 1'b0;
      ProductSum_for_asn_73_itm_1 <= 1'b0;
      ProductSum_for_asn_82_itm_1 <= 1'b0;
      ProductSum_for_asn_98_itm_1 <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1 <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_1 <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1 <= 1'b0;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_1_1 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_1 <= 1'b0;
    end
    else if ( PECoreRun_wen ) begin
      reg_PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_cgo_ir_cse <=
          and_480_rmff;
      reg_PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_cgo_ir_cse <=
          and_483_rmff;
      reg_weight_mem_banks_bank_a1_a1_a1_a_rsci_cgo_ir_cse <= and_487_rmff;
      reg_weight_mem_banks_bank_a1_a1_a0_a_rsci_cgo_ir_cse <= and_490_rmff;
      reg_weight_mem_banks_bank_a1_a0_a1_a_rsci_cgo_ir_cse <= and_494_rmff;
      reg_weight_mem_banks_bank_a1_a0_a0_a_rsci_cgo_ir_cse <= and_498_rmff;
      reg_weight_mem_banks_bank_a0_a1_a1_a_rsci_cgo_ir_cse <= and_502_rmff;
      reg_weight_mem_banks_bank_a0_a1_a0_a_rsci_cgo_ir_cse <= and_506_rmff;
      reg_weight_mem_banks_bank_a0_a0_a1_a_rsci_cgo_ir_cse <= and_510_rmff;
      reg_weight_mem_banks_bank_a0_a0_a0_a_rsci_cgo_ir_cse <= and_514_rmff;
      reg_rva_out_Push_mioi_iswt0_cse <= and_516_cse;
      reg_start_PopNB_mioi_iswt0_cse <= and_518_rmff;
      reg_act_port_Push_mioi_iswt0_cse <= and_520_rmff;
      reg_rva_in_PopNB_mioi_iswt0_cse <= fsm_output;
      pe_config_manager_counter_sva_dfm_3_1 <= MUX_v_4_2_2(4'b0000, operator_4_false_acc_nl,
          pe_config_UpdateManagerCounter_if_not_7_nl);
      pe_config_UpdateInputCounter_pe_config_UpdateInputCounter_if_nor_mdf_sva_st_1
          <= ~((pe_config_input_counter_sva_mx1 != (operator_16_false_acc_sdt_sva_1[7:0]))
          | (operator_16_false_acc_sdt_sva_1[8]));
      pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1
          <= pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1_1;
      while_stage_0_3 <= reg_rva_in_PopNB_mioi_iswt0_cse;
      while_stage_0_4 <= while_stage_0_3;
      while_stage_0_5 <= while_stage_0_4;
      while_stage_0_6 <= while_stage_0_5;
      while_stage_0_7 <= while_stage_0_6;
      while_stage_0_8 <= while_stage_0_7;
      while_stage_0_9 <= while_stage_0_8;
      while_stage_0_10 <= while_stage_0_9;
      while_stage_0_11 <= while_stage_0_10;
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_122_itm_1 <= pe_manager_base_weight_sva_mx1_3_0[1];
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_95_itm_1 <= pe_manager_base_weight_sva_mx2[2];
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_93_itm_1 <= pe_manager_base_weight_sva_mx1_3_0[0];
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_1_itm_1 <= ~ (pe_manager_base_weight_sva_mx1_3_0[1]);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_1 <= (pe_manager_base_weight_sva_mx2[2])
          & (pe_manager_base_weight_sva_mx1_3_0[1:0]==2'b01) & weight_mem_run_3_for_land_1_lpi_1_dfm_1_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_1
          <= ~((pe_manager_base_weight_sva_mx2[2]) | (pe_manager_base_weight_sva_mx1_3_0[1:0]!=2'b00));
      input_read_addrs_sva_1_1 <= nl_input_read_addrs_sva_1_1[7:0];
      ProductSum_for_asn_64_itm_1 <= MUX1HOT_s_1_3_2(accum_vector_data_3_sva_1_load_mx0w0,
          accum_vector_data_3_sva_1_load, while_if_while_if_and_12_nl, {and_dcpl_611
          , and_dcpl_612 , rva_in_PopNB_mioi_return_rsc_z_mxwt});
      ProductSum_for_asn_73_itm_1 <= MUX_s_1_2_2(accum_vector_data_2_sva_1_load_mx0w0,
          accum_vector_data_2_sva_1_load, or_dcpl_616);
      ProductSum_for_asn_82_itm_1 <= MUX_s_1_2_2(accum_vector_data_1_sva_1_load_mx0w0,
          accum_vector_data_1_sva_1_load, or_dcpl_616);
      ProductSum_for_asn_98_itm_1 <= MUX_s_1_2_2(accum_vector_data_0_sva_1_load_mx0w0,
          accum_vector_data_0_sva_1_load, or_dcpl_616);
      PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1 <= MUX1HOT_s_1_3_2(PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_mx0w0,
          accum_vector_data_6_sva_1_load_mx0w1, accum_vector_data_6_sva_1_load, {rva_in_PopNB_mioi_return_rsc_z_mxwt
          , and_dcpl_611 , and_dcpl_612});
      PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_1 <= MUX1HOT_s_1_3_2(and_321_cse,
          accum_vector_data_7_sva_1_load_mx0w1, accum_vector_data_7_sva_1_load, {rva_in_PopNB_mioi_return_rsc_z_mxwt
          , and_dcpl_611 , and_dcpl_612});
      PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1 <= MUX1HOT_s_1_3_2(PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_mx0w0,
          accum_vector_data_5_sva_1_load_mx0w1, accum_vector_data_5_sva_1_load, {rva_in_PopNB_mioi_return_rsc_z_mxwt
          , and_dcpl_611 , and_dcpl_612});
      PECore_RunScale_PECore_RunScale_if_and_1_svs_1_1 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_1;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_1 <= MUX1HOT_s_1_3_2(PECore_DecodeAxiRead_switch_lp_nor_tmp_mx0w0,
          accum_vector_data_4_sva_1_load_mx0w1, accum_vector_data_4_sva_1_load, {rva_in_PopNB_mioi_return_rsc_z_mxwt
          , and_dcpl_611 , and_dcpl_612});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_9 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_9 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_9 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_2_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_8 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_1_7;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_9 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_8;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_9 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_8;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_9 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_9 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_78_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_9 <= rva_out_reg_data_15_9_sva_dfm_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_23_17_sva_dfm_7 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_79_enex5 ) begin
      rva_out_reg_data_23_17_sva_dfm_7 <= rva_out_reg_data_23_17_sva_dfm_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_7 <= 6'b000000;
    end
    else if ( rva_out_reg_data_and_80_enex5 ) begin
      rva_out_reg_data_30_25_sva_dfm_7 <= rva_out_reg_data_30_25_sva_dfm_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_63_sva_dfm_4_4 <= 1'b0;
      rva_out_reg_data_47_sva_dfm_4_4 <= 1'b0;
      reg_rva_out_reg_data_46_40_sva_dfm_4_4_ftd <= 3'b000;
      reg_rva_out_reg_data_39_36_sva_dfm_4_4_ftd <= 1'b0;
      reg_rva_out_reg_data_39_36_sva_dfm_4_4_ftd_1 <= 1'b0;
      reg_rva_out_reg_data_39_36_sva_dfm_4_4_ftd_2 <= 2'b00;
      input_read_req_valid_lpi_1_dfm_1_9 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( rva_out_reg_data_and_17_cse ) begin
      rva_out_reg_data_63_sva_dfm_4_4 <= reg_PECore_RunMac_PECore_RunMac_if_and_svs_st_8_cse;
      rva_out_reg_data_47_sva_dfm_4_4 <= PECore_PushOutput_PECore_PushOutput_if_and_svs_st_8;
      reg_rva_out_reg_data_46_40_sva_dfm_4_4_ftd <= rva_out_reg_data_46_40_sva_dfm_4_3_rsp_0;
      reg_rva_out_reg_data_39_36_sva_dfm_4_4_ftd <= rva_out_reg_data_39_36_sva_dfm_4_3_rsp_0;
      reg_rva_out_reg_data_39_36_sva_dfm_4_4_ftd_1 <= rva_out_reg_data_39_36_sva_dfm_4_3_rsp_1;
      reg_rva_out_reg_data_39_36_sva_dfm_4_4_ftd_2 <= rva_out_reg_data_39_36_sva_dfm_4_3_rsp_2;
      input_read_req_valid_lpi_1_dfm_1_9 <= input_read_req_valid_lpi_1_dfm_1_8;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_56_sva_dfm_4_4 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_81_enex5 ) begin
      rva_out_reg_data_62_56_sva_dfm_4_4 <= rva_out_reg_data_62_56_sva_dfm_4_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_4_ftd <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_82_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_4_ftd <= rva_out_reg_data_55_48_sva_dfm_4_3_rsp_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_4_ftd_1 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_83_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_4_ftd_1 <= rva_out_reg_data_55_48_sva_dfm_4_3_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_4_ftd_1 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_84_enex5 ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_4_ftd_1 <= rva_out_reg_data_46_40_sva_dfm_4_3_rsp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_4_4 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_85_enex5 ) begin
      rva_out_reg_data_35_32_sva_dfm_4_4 <= rva_out_reg_data_35_32_sva_dfm_4_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_2 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_2 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_2
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_2
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_2
          <= 1'b0;
    end
    else if ( input_mem_banks_read_read_data_and_cse ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_2 <=
          input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_1;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_2 <=
          input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_1;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_2
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_1;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_2
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_1;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_2
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_slc_weight_port_read_out_data_0_0_0_itm_1 <= 1'b0;
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_1_ftd
          <= 1'b0;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_1_0_itm_1 <= 1'b0;
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_1_ftd
          <= 1'b0;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_0_itm_1 <= 1'b0;
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_ftd
          <= 1'b0;
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_ftd_1
          <= 1'b0;
      reg_weight_port_read_out_data_0_3_sva_dfm_4_ftd <= 1'b0;
      reg_weight_port_read_out_data_0_3_sva_dfm_4_ftd_1 <= 3'b000;
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_1_ftd_1_rsp_0
          <= 1'b0;
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_1_ftd_1_rsp_0
          <= 3'b000;
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_1_ftd_1_rsp_1
          <= 3'b000;
    end
    else if ( weight_port_read_out_data_and_68_cse ) begin
      weight_port_read_out_data_slc_weight_port_read_out_data_0_0_0_itm_1 <= weight_port_read_out_data_0_0_sva_dfm_3_rsp_1_5_0[0];
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_1_ftd
          <= weight_port_read_out_data_0_0_sva_dfm_3_rsp_0;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_1_0_itm_1 <= weight_port_read_out_data_0_1_sva_dfm_3_rsp_1_3_0[0];
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_1_ftd
          <= weight_port_read_out_data_0_1_sva_dfm_3_rsp_0;
      weight_port_read_out_data_slc_weight_port_read_out_data_0_2_0_itm_1 <= weight_port_read_out_data_0_2_sva_dfm_3_rsp_2[0];
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_ftd
          <= weight_port_read_out_data_0_2_sva_dfm_3_rsp_0;
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_ftd_1
          <= weight_port_read_out_data_0_2_sva_dfm_3_rsp_1;
      reg_weight_port_read_out_data_0_3_sva_dfm_4_ftd <= weight_port_read_out_data_0_3_sva_dfm_3_rsp_0;
      reg_weight_port_read_out_data_0_3_sva_dfm_4_ftd_1 <= weight_port_read_out_data_0_3_sva_dfm_3_rsp_1;
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_1_ftd_1_rsp_0
          <= weight_port_read_out_data_0_0_sva_dfm_3_rsp_1_6;
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_1_ftd_1_rsp_0
          <= weight_port_read_out_data_0_1_sva_dfm_3_rsp_1_6_4;
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_1_7_1_itm_1_ftd_1_rsp_1
          <= weight_port_read_out_data_0_1_sva_dfm_3_rsp_1_3_0[3:1];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_22_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_2
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_23_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_2
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_24_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_2
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_ftd_2
          <= 5'b00000;
    end
    else if ( weight_port_read_out_data_and_104_enex5 ) begin
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_2_7_1_itm_1_ftd_2
          <= weight_port_read_out_data_0_2_sva_dfm_3_rsp_2[5:1];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_4_ftd_2 <= 4'b0000;
    end
    else if ( weight_port_read_out_data_and_105_enex5 ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_4_ftd_2 <= weight_port_read_out_data_0_3_sva_dfm_3_rsp_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2
          <= 6'b000000;
    end
    else if ( input_mem_banks_read_read_data_and_25_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_2
          <= input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_9 <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_9
          <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_cse ) begin
      rva_in_reg_rw_sva_9 <= rva_in_reg_rw_sva_8;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_9
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_st_1_9 <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_4 ) begin
      rva_in_reg_rw_sva_st_1_9 <= rva_in_reg_rw_sva_st_1_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_9
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_9
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_7
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_7
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_9
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_8;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_9
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_8;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_7
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_6;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_7
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_0_sva_dfm_6 <= 1'b0;
      rva_out_reg_data_8_sva_dfm_6 <= 1'b0;
      rva_out_reg_data_16_sva_dfm_6 <= 1'b0;
      rva_out_reg_data_31_sva_dfm_6 <= 1'b0;
      rva_out_reg_data_24_sva_dfm_6 <= 1'b0;
      rva_out_reg_data_7_1_sva_dfm_6_rsp_0 <= 1'b0;
      rva_out_reg_data_15_9_sva_dfm_6_rsp_0 <= 1'b0;
      rva_out_reg_data_23_17_sva_dfm_6_rsp_0 <= 1'b0;
      rva_out_reg_data_23_17_sva_dfm_6_rsp_1 <= 1'b0;
      rva_out_reg_data_23_17_sva_dfm_6_rsp_2 <= 5'b00000;
      rva_out_reg_data_30_25_sva_dfm_6_rsp_0 <= 3'b000;
      rva_out_reg_data_30_25_sva_dfm_6_rsp_1 <= 3'b000;
      rva_out_reg_data_7_1_sva_dfm_6_rsp_1_rsp_0 <= 1'b0;
      rva_out_reg_data_7_1_sva_dfm_6_rsp_1_rsp_1 <= 5'b00000;
      rva_out_reg_data_15_9_sva_dfm_6_rsp_1_rsp_0 <= 3'b000;
      rva_out_reg_data_15_9_sva_dfm_6_rsp_1_rsp_1 <= 3'b000;
    end
    else if ( rva_out_reg_data_and_cse ) begin
      rva_out_reg_data_0_sva_dfm_6 <= MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_14_itm,
          weight_port_read_out_data_slc_weight_port_read_out_data_0_0_0_itm_1, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7);
      rva_out_reg_data_8_sva_dfm_6 <= MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_15_itm,
          weight_port_read_out_data_slc_weight_port_read_out_data_0_1_0_itm_1, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7);
      rva_out_reg_data_16_sva_dfm_6 <= MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_16_itm,
          weight_port_read_out_data_slc_weight_port_read_out_data_0_2_0_itm_1, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_7);
      rva_out_reg_data_31_sva_dfm_6 <= PECore_PushAxiRsp_if_mux1h_17;
      rva_out_reg_data_24_sva_dfm_6 <= PECore_PushAxiRsp_if_mux1h_15;
      rva_out_reg_data_7_1_sva_dfm_6_rsp_0 <= PECore_PushAxiRsp_if_mux1h_10_6;
      rva_out_reg_data_15_9_sva_dfm_6_rsp_0 <= PECore_PushAxiRsp_if_mux1h_12_6;
      rva_out_reg_data_23_17_sva_dfm_6_rsp_0 <= PECore_PushAxiRsp_if_mux1h_14_6;
      rva_out_reg_data_23_17_sva_dfm_6_rsp_1 <= PECore_PushAxiRsp_if_mux1h_14_5;
      rva_out_reg_data_23_17_sva_dfm_6_rsp_2 <= PECore_PushAxiRsp_if_mux1h_14_4_0;
      rva_out_reg_data_30_25_sva_dfm_6_rsp_0 <= PECore_PushAxiRsp_if_mux1h_16_5_3;
      rva_out_reg_data_30_25_sva_dfm_6_rsp_1 <= PECore_PushAxiRsp_if_mux1h_16_2_0;
      rva_out_reg_data_7_1_sva_dfm_6_rsp_1_rsp_0 <= PECore_PushAxiRsp_if_mux1h_10_5;
      rva_out_reg_data_7_1_sva_dfm_6_rsp_1_rsp_1 <= PECore_PushAxiRsp_if_mux1h_10_4_0;
      rva_out_reg_data_15_9_sva_dfm_6_rsp_1_rsp_0 <= PECore_PushAxiRsp_if_mux1h_12_5_3;
      rva_out_reg_data_15_9_sva_dfm_6_rsp_1_rsp_1 <= PECore_PushAxiRsp_if_mux1h_12_2_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_reg_data_243_224_sva_dfm_1_1 <= 20'b00000000000000000000;
      act_port_reg_data_19_0_sva_dfm_1_1 <= 20'b00000000000000000000;
      act_port_reg_data_211_192_sva_dfm_1_1 <= 20'b00000000000000000000;
      act_port_reg_data_51_32_sva_dfm_1_1 <= 20'b00000000000000000000;
      act_port_reg_data_179_160_sva_dfm_1_1 <= 20'b00000000000000000000;
      act_port_reg_data_83_64_sva_dfm_1_1 <= 20'b00000000000000000000;
      act_port_reg_data_147_128_sva_dfm_1_1 <= 20'b00000000000000000000;
      act_port_reg_data_115_96_sva_dfm_1_1 <= 20'b00000000000000000000;
    end
    else if ( and_1002_cse ) begin
      act_port_reg_data_243_224_sva_dfm_1_1 <= MUX_v_20_2_2((readslicef_31_20_11(PECore_RunScale_if_for_8_mul_1_nl)),
          act_port_reg_data_243_224_sva_mx1, or_dcpl_603);
      act_port_reg_data_19_0_sva_dfm_1_1 <= MUX_v_20_2_2((readslicef_31_20_11(PECore_RunScale_if_for_1_mul_1_nl)),
          act_port_reg_data_19_0_sva_mx1, or_dcpl_603);
      act_port_reg_data_211_192_sva_dfm_1_1 <= MUX_v_20_2_2((readslicef_31_20_11(PECore_RunScale_if_for_7_mul_1_nl)),
          act_port_reg_data_211_192_sva_mx1, or_dcpl_603);
      act_port_reg_data_51_32_sva_dfm_1_1 <= MUX_v_20_2_2((readslicef_31_20_11(PECore_RunScale_if_for_2_mul_1_nl)),
          act_port_reg_data_51_32_sva_mx1, or_dcpl_603);
      act_port_reg_data_179_160_sva_dfm_1_1 <= MUX_v_20_2_2((readslicef_31_20_11(PECore_RunScale_if_for_6_mul_1_nl)),
          act_port_reg_data_179_160_sva_mx1, or_dcpl_603);
      act_port_reg_data_83_64_sva_dfm_1_1 <= MUX_v_20_2_2((readslicef_31_20_11(PECore_RunScale_if_for_3_mul_1_nl)),
          act_port_reg_data_83_64_sva_mx1, or_dcpl_603);
      act_port_reg_data_147_128_sva_dfm_1_1 <= MUX_v_20_2_2((readslicef_31_20_11(PECore_RunScale_if_for_5_mul_1_nl)),
          act_port_reg_data_147_128_sva_mx1, or_dcpl_603);
      act_port_reg_data_115_96_sva_dfm_1_1 <= MUX_v_20_2_2((readslicef_31_20_11(PECore_RunScale_if_for_4_mul_1_nl)),
          act_port_reg_data_115_96_sva_mx1, or_dcpl_603);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_9 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_9 <= 1'b0;
    end
    else if ( PECore_PushOutput_if_and_cse ) begin
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_9 <= PECore_PushOutput_PECore_PushOutput_if_and_svs_st_8;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_9 <= PECore_UpdateFSM_switch_lp_equal_tmp_2_8;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_st_1_8 <= 1'b0;
      rva_in_reg_rw_sva_st_8 <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_2_cse ) begin
      rva_in_reg_rw_sva_st_1_8 <= rva_in_reg_rw_sva_st_1_7;
      rva_in_reg_rw_sva_st_8 <= rva_in_reg_rw_sva_st_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_PECore_RunMac_PECore_RunMac_if_and_svs_st_8_cse <= 1'b0;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_8 <= 1'b0;
    end
    else if ( PECore_RunMac_if_and_cse ) begin
      reg_PECore_RunMac_PECore_RunMac_if_and_svs_st_8_cse <= PECore_RunMac_PECore_RunMac_if_and_svs_st_7;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_8 <= PECore_PushOutput_PECore_PushOutput_if_and_svs_st_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8
          <= 1'b0;
      rva_in_reg_rw_sva_8 <= 1'b0;
      accum_vector_data_acc_30_itm_1 <= 23'b00000000000000000000000;
      accum_vector_data_acc_28_itm_1 <= 23'b00000000000000000000000;
      accum_vector_data_acc_25_itm_1 <= 23'b00000000000000000000000;
      accum_vector_data_acc_22_itm_1 <= 23'b00000000000000000000000;
      accum_vector_data_acc_19_itm_1 <= 23'b00000000000000000000000;
      accum_vector_data_acc_13_itm_1 <= 23'b00000000000000000000000;
      accum_vector_data_acc_10_itm_1 <= 23'b00000000000000000000000;
    end
    else if ( while_if_and_6_cse ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7;
      rva_in_reg_rw_sva_8 <= rva_in_reg_rw_sva_7;
      accum_vector_data_acc_30_itm_1 <= nl_accum_vector_data_acc_30_itm_1[22:0];
      accum_vector_data_acc_28_itm_1 <= nl_accum_vector_data_acc_28_itm_1[22:0];
      accum_vector_data_acc_25_itm_1 <= nl_accum_vector_data_acc_25_itm_1[22:0];
      accum_vector_data_acc_22_itm_1 <= nl_accum_vector_data_acc_22_itm_1[22:0];
      accum_vector_data_acc_19_itm_1 <= nl_accum_vector_data_acc_19_itm_1[22:0];
      accum_vector_data_acc_13_itm_1 <= nl_accum_vector_data_acc_13_itm_1[22:0];
      accum_vector_data_acc_10_itm_1 <= nl_accum_vector_data_acc_10_itm_1[22:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_st_1_7 <= 1'b0;
      rva_in_reg_rw_sva_st_7 <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_3_cse ) begin
      rva_in_reg_rw_sva_st_1_7 <= rva_in_reg_rw_sva_st_1_6;
      rva_in_reg_rw_sva_st_7 <= rva_in_reg_rw_sva_st_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_7 <= 1'b0;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_7 <= 1'b0;
    end
    else if ( PECore_RunMac_if_and_1_cse ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_7 <= PECore_RunMac_PECore_RunMac_if_and_svs_st_6;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_7 <= PECore_PushOutput_PECore_PushOutput_if_and_svs_st_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7
          <= 1'b0;
      rva_in_reg_rw_sva_7 <= 1'b0;
    end
    else if ( while_if_and_7_cse ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6;
      rva_in_reg_rw_sva_7 <= rva_in_reg_rw_sva_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ProductSum_for_asn_12_itm_6 <= 1'b0;
      weight_port_read_out_data_7_3_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_7_2_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_7_5_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_7_4_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_7_7_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_7_6_sva_dfm_1 <= 8'b00000000;
      ProductSum_for_asn_23_itm_6 <= 1'b0;
      weight_mem_run_3_for_5_mux_51_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_50_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_53_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_52_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_55_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_54_itm_1 <= 8'b00000000;
      ProductSum_for_asn_38_itm_6 <= 1'b0;
      weight_port_read_out_data_5_3_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_5_2_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_5_5_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_5_4_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_5_7_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_5_6_sva_dfm_1 <= 8'b00000000;
      ProductSum_for_asn_49_itm_6 <= 1'b0;
      weight_mem_run_3_for_5_mux_35_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_34_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_37_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_36_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_39_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_38_itm_1 <= 8'b00000000;
      ProductSum_for_asn_62_itm_6 <= 1'b0;
      weight_mem_run_3_for_5_mux_27_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_26_itm_1 <= 8'b00000000;
      weight_port_read_out_data_3_5_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_3_4_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_3_7_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_3_6_sva_dfm_1 <= 8'b00000000;
      ProductSum_for_asn_72_itm_6 <= 1'b0;
      weight_mem_run_3_for_5_mux_19_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_18_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_21_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_20_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_23_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_22_itm_1 <= 8'b00000000;
      ProductSum_for_asn_80_itm_6 <= 1'b0;
      weight_mem_run_3_for_5_mux_13_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_15_itm_1 <= 8'b00000000;
      weight_mem_run_3_for_5_mux_14_itm_1 <= 8'b00000000;
      ProductSum_for_asn_94_itm_6 <= 1'b0;
      weight_port_read_out_data_0_7_sva_dfm_1_1_rsp_0 <= 1'b0;
      weight_port_read_out_data_0_7_sva_dfm_1_1_rsp_1 <= 7'b0000000;
      weight_mem_run_3_for_5_mux_6_itm_1_7_4 <= 4'b0000;
      weight_mem_run_3_for_5_mux_6_itm_1_3_0 <= 4'b0000;
    end
    else if ( ProductSum_for_and_cse ) begin
      ProductSum_for_asn_12_itm_6 <= ProductSum_for_asn_16_itm_5;
      weight_port_read_out_data_7_3_sva_dfm_1 <= weight_port_read_out_data_7_3_sva_dfm_2;
      weight_port_read_out_data_7_2_sva_dfm_1 <= weight_port_read_out_data_7_2_sva_dfm_2;
      weight_port_read_out_data_7_5_sva_dfm_1 <= weight_port_read_out_data_7_5_sva_dfm_2;
      weight_port_read_out_data_7_4_sva_dfm_1 <= weight_port_read_out_data_7_4_sva_dfm_2;
      weight_port_read_out_data_7_7_sva_dfm_1 <= weight_port_read_out_data_7_7_sva_dfm_2;
      weight_port_read_out_data_7_6_sva_dfm_1 <= weight_port_read_out_data_7_6_sva_dfm_2;
      ProductSum_for_asn_23_itm_6 <= ProductSum_for_asn_25_itm_5;
      weight_mem_run_3_for_5_mux_51_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_6_3_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2,
          weight_mem_run_3_for_land_7_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_50_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_6_2_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_3_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2,
          weight_mem_run_3_for_land_7_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_53_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_6_5_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_6_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2,
          weight_mem_run_3_for_land_7_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_52_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_6_4_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_5_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2,
          weight_mem_run_3_for_land_7_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_55_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_6_7_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2,
          weight_mem_run_3_for_land_7_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_54_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_6_6_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2,
          weight_mem_run_3_for_land_7_lpi_1_dfm_2);
      ProductSum_for_asn_38_itm_6 <= ProductSum_for_asn_42_itm_5;
      weight_port_read_out_data_5_3_sva_dfm_1 <= weight_port_read_out_data_5_3_sva_dfm_2;
      weight_port_read_out_data_5_2_sva_dfm_1 <= weight_port_read_out_data_5_2_sva_dfm_2;
      weight_port_read_out_data_5_5_sva_dfm_1 <= weight_port_read_out_data_5_5_sva_dfm_2;
      weight_port_read_out_data_5_4_sva_dfm_1 <= weight_port_read_out_data_5_4_sva_dfm_2;
      weight_port_read_out_data_5_7_sva_dfm_1 <= weight_port_read_out_data_5_7_sva_dfm_2;
      weight_port_read_out_data_5_6_sva_dfm_1 <= weight_port_read_out_data_5_6_sva_dfm_2;
      ProductSum_for_asn_49_itm_6 <= ProductSum_for_asn_51_itm_5;
      weight_mem_run_3_for_5_mux_35_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_4_3_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2,
          weight_mem_run_3_for_land_5_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_34_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_4_2_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_3_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2,
          weight_mem_run_3_for_land_5_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_37_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_4_5_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_6_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2,
          weight_mem_run_3_for_land_5_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_36_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_4_4_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_5_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2,
          weight_mem_run_3_for_land_5_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_39_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_4_7_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2,
          weight_mem_run_3_for_land_5_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_38_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_4_6_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2,
          weight_mem_run_3_for_land_5_lpi_1_dfm_2);
      ProductSum_for_asn_62_itm_6 <= ProductSum_for_asn_64_itm_5;
      weight_mem_run_3_for_5_mux_27_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_3_3_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000002,
          weight_mem_run_3_for_land_4_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_26_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_3_2_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000003,
          weight_mem_run_3_for_land_4_lpi_1_dfm_2);
      weight_port_read_out_data_3_5_sva_dfm_1 <= weight_port_read_out_data_3_5_sva_dfm_2;
      weight_port_read_out_data_3_4_sva_dfm_1 <= weight_port_read_out_data_3_4_sva_dfm_2;
      weight_port_read_out_data_3_7_sva_dfm_1 <= weight_port_read_out_data_3_7_sva_dfm_2;
      weight_port_read_out_data_3_6_sva_dfm_1 <= weight_port_read_out_data_3_6_sva_dfm_2;
      ProductSum_for_asn_72_itm_6 <= ProductSum_for_asn_73_itm_5;
      weight_mem_run_3_for_5_mux_19_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_2_3_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000006,
          weight_mem_run_3_for_land_3_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_18_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_2_2_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000005,
          weight_mem_run_3_for_land_3_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_21_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_2_5_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000003,
          weight_mem_run_3_for_land_3_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_20_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_2_4_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000004,
          weight_mem_run_3_for_land_3_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_23_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_2_7_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_pmx_sva_1,
          weight_mem_run_3_for_land_3_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_22_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_2_6_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000002,
          weight_mem_run_3_for_land_3_lpi_1_dfm_2);
      ProductSum_for_asn_80_itm_6 <= ProductSum_for_asn_82_itm_5;
      weight_mem_run_3_for_5_mux_13_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_1_5_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000004,
          weight_mem_run_3_for_land_2_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_15_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_1_7_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_pmx_000000,
          weight_mem_run_3_for_land_2_lpi_1_dfm_2);
      weight_mem_run_3_for_5_mux_14_itm_1 <= MUX_v_8_2_2(weight_port_read_out_data_1_6_sva_dfm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000006,
          weight_mem_run_3_for_land_2_lpi_1_dfm_2);
      ProductSum_for_asn_94_itm_6 <= ProductSum_for_asn_98_itm_5;
      weight_port_read_out_data_0_7_sva_dfm_1_1_rsp_0 <= weight_port_read_out_data_0_7_sva_dfm_1_1_mx0_7;
      weight_port_read_out_data_0_7_sva_dfm_1_1_rsp_1 <= weight_port_read_out_data_0_7_sva_dfm_1_1_mx0_6_0;
      weight_mem_run_3_for_5_mux_6_itm_1_7_4 <= MUX_v_4_2_2(weight_port_read_out_data_0_6_sva_dfm_2_7_4,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000000[7:4]),
          weight_mem_run_3_for_land_1_lpi_1_dfm_3);
      weight_mem_run_3_for_5_mux_6_itm_1_3_0 <= MUX_v_4_2_2(weight_port_read_out_data_0_6_sva_dfm_2_3_0,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000000[3:0]),
          weight_mem_run_3_for_land_1_lpi_1_dfm_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_5_63_16 <= 48'b000000000000000000000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_1_read_data_and_enex5 ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_5_63_16 <= input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[63:16];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_5_7_0 <= 8'b00000000;
    end
    else if ( input_mem_banks_read_1_read_data_and_6_enex5 ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_5_7_0 <= input_mem_banks_read_1_read_data_lpi_1_dfm_1_4[7:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_0_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_enex5 ) begin
      weight_port_read_out_data_2_0_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000001;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000001
          <= 8'b00000000;
    end
    else if ( data_in_tmp_operator_2_for_and_tmp ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000001
          <= MUX_v_8_8_2((input_mem_banks_read_read_data_lpi_1_dfm_1_4[7:0]), (weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1[7:0]),
          (weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1[7:0]),
          (weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1[7:0]), (weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1[7:0]),
          (weight_mem_banks_read_1_read_data_7_lpi_1_dfm_mx0[7:0]), BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9,
          {weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 , pe_manager_base_weight_slc_pe_manager_base_weight_0_12_itm_2});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_run_3_for_land_3_lpi_1_dfm_3 <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6
          <= 1'b0;
      rva_in_reg_rw_sva_6 <= 1'b0;
    end
    else if ( weight_mem_run_3_for_aelse_and_cse ) begin
      weight_mem_run_3_for_land_3_lpi_1_dfm_3 <= weight_mem_run_3_for_land_3_lpi_1_dfm_2;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5;
      rva_in_reg_rw_sva_6 <= rva_in_reg_rw_sva_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_run_3_for_5_mux_11_itm_1_7 <= 1'b0;
      weight_mem_run_3_for_5_mux_11_itm_1_6_0 <= 7'b0000000;
      weight_mem_run_3_for_5_mux_10_itm_1_7 <= 1'b0;
      weight_mem_run_3_for_5_mux_10_itm_1_6_0 <= 7'b0000000;
      weight_mem_run_3_for_5_mux_12_itm_1_7_6 <= 2'b00;
      weight_mem_run_3_for_5_mux_12_itm_1_5_0 <= 6'b000000;
    end
    else if ( weight_mem_run_3_for_5_and_209_ssc ) begin
      weight_mem_run_3_for_5_mux_11_itm_1_7 <= MUX_s_1_2_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000002[7]),
          (weight_port_read_out_data_1_3_sva_dfm_1[7]), and_dcpl_505);
      weight_mem_run_3_for_5_mux_11_itm_1_6_0 <= MUX1HOT_v_7_3_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000002[6:0]),
          (weight_port_read_out_data_1_3_sva_dfm_1[6:0]), weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1_6_0,
          {and_dcpl_504 , and_dcpl_505 , while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5});
      weight_mem_run_3_for_5_mux_10_itm_1_7 <= MUX_s_1_2_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000003[7]),
          (weight_port_read_out_data_1_2_sva_dfm_1[7]), and_dcpl_505);
      weight_mem_run_3_for_5_mux_10_itm_1_6_0 <= MUX1HOT_v_7_3_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000003[6:0]),
          (weight_port_read_out_data_1_2_sva_dfm_1[6:0]), weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_itm_1_6_0,
          {and_dcpl_504 , and_dcpl_505 , while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5});
      weight_mem_run_3_for_5_mux_12_itm_1_7_6 <= MUX_v_2_2_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000005[7:6]),
          (weight_port_read_out_data_1_4_sva_dfm_1[7:6]), and_dcpl_505);
      weight_mem_run_3_for_5_mux_12_itm_1_5_0 <= MUX1HOT_v_6_3_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000005[5:0]),
          (weight_port_read_out_data_1_4_sva_dfm_1[5:0]), weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_itm_1_5_0,
          {and_dcpl_504 , and_dcpl_505 , while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_6 <= 1'b0;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_6 <= 1'b0;
    end
    else if ( PECore_RunMac_if_and_2_cse ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_6 <= MUX1HOT_s_1_3_2(PECore_RunMac_PECore_RunMac_if_and_svs_st_5,
          weight_port_read_out_data_0_7_sva_dfm_3_7, PECore_PushAxiRsp_if_else_mux_13_mx0w2,
          {(~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
          , while_and_24_cse , while_and_23_cse});
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_6 <= MUX1HOT_s_1_3_2(PECore_PushOutput_PECore_PushOutput_if_and_svs_st_5,
          (weight_port_read_out_data_0_5_sva_dfm_3_7_4[3]), PECore_PushAxiRsp_if_else_mux_10_mx0w2,
          {(~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
          , while_and_24_cse , while_and_23_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_3
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_44_itm_1)
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
        & while_stage_0_6 ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_3
          <= weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_3
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_54_itm_1)
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
        & while_stage_0_6 ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_3
          <= weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_st_1_5 <= 1'b0;
      rva_in_reg_rw_sva_st_5 <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_4_cse ) begin
      rva_in_reg_rw_sva_st_1_5 <= rva_in_reg_rw_sva_st_1_4;
      rva_in_reg_rw_sva_st_5 <= rva_in_reg_rw_sva_st_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      PECore_RunMac_PECore_RunMac_if_and_svs_st_5 <= 1'b0;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_13_itm_2 <= 1'b0;
      weight_mem_run_3_for_land_lpi_1_dfm_2 <= 1'b0;
      weight_mem_run_3_for_5_and_110_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_111_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_112_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_12_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_102_itm_2 <= 1'b0;
      weight_mem_run_3_for_5_and_103_itm_2 <= 1'b0;
      weight_read_addrs_7_lpi_1_dfm_3_2_0 <= 3'b000;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_5_itm_2 <= 1'b0;
      weight_mem_run_3_for_land_6_lpi_1_dfm_2 <= 1'b0;
      weight_mem_run_3_for_5_and_44_itm_2 <= 1'b0;
      weight_mem_run_3_for_5_and_46_itm_2 <= 1'b0;
      weight_mem_run_3_for_5_and_47_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_48_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_38_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_39_itm_2 <= 1'b0;
      weight_read_addrs_5_lpi_1_dfm_3_2_0 <= 3'b000;
      reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_20_itm_2_cse <= 1'b0;
      weight_mem_run_3_for_5_and_162_itm_2 <= 1'b0;
      reg_weight_mem_run_3_for_5_and_163_itm_2_cse <= 1'b0;
      weight_mem_run_3_for_5_and_164_itm_2 <= 1'b0;
      reg_weight_mem_run_3_for_5_and_165_itm_2_cse <= 1'b0;
      reg_weight_mem_run_3_for_5_and_166_itm_2_cse <= 1'b0;
      reg_weight_mem_run_3_for_5_and_167_itm_2_cse <= 1'b0;
      reg_weight_mem_run_3_for_5_and_168_itm_2_cse <= 1'b0;
      weight_read_addrs_3_lpi_1_dfm_3_2_0 <= 3'b000;
      weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      weight_mem_run_3_for_5_and_156_itm_2 <= 1'b0;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_10_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_84_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_3_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_28_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_30_itm_2 <= 1'b0;
      weight_mem_run_3_for_5_and_31_itm_2 <= 1'b0;
      weight_mem_run_3_for_5_and_20_itm_2 <= 1'b0;
      weight_mem_run_3_for_5_and_22_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_23_itm_1 <= 1'b0;
      reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_2_cse <= 1'b0;
      weight_mem_run_3_for_5_and_8_itm_1 <= 1'b0;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_5 <= 1'b0;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_5 <= 1'b0;
      accum_vector_operator_1_for_asn_70_itm_4 <= 1'b0;
      accum_vector_operator_1_for_asn_61_itm_4 <= 1'b0;
      accum_vector_operator_1_for_asn_52_itm_4 <= 1'b0;
      accum_vector_operator_1_for_asn_43_itm_4 <= 1'b0;
      accum_vector_operator_1_for_asn_34_itm_4 <= 1'b0;
      accum_vector_operator_1_for_asn_25_itm_4 <= 1'b0;
      accum_vector_operator_1_for_asn_16_itm_4 <= 1'b0;
      accum_vector_operator_1_for_asn_7_itm_4 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_5 <= 1'b0;
    end
    else if ( weight_mem_banks_read_1_read_data_and_8_cse ) begin
      weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1 <= MUX_v_64_2_2(weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1_1,
          weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d, weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
      weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1 <= MUX_v_64_2_2(weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1_1,
          weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d, weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
      weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1 <= MUX_v_64_2_2(weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1_1,
          weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d, weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
      weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1 <= MUX_v_64_2_2(weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1_1,
          weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d, weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
      weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1 <= MUX_v_64_2_2(weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1_1,
          weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d, weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
      PECore_RunMac_PECore_RunMac_if_and_svs_st_5 <= reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_13_itm_2 <= weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_13_itm_1;
      weight_mem_run_3_for_land_lpi_1_dfm_2 <= weight_mem_run_3_for_land_lpi_1_dfm_1;
      weight_mem_run_3_for_5_and_110_itm_1 <= (weight_read_addrs_7_lpi_1_dfm_2_2_0==3'b101)
          & weight_mem_run_3_for_land_lpi_1_dfm_1;
      weight_mem_run_3_for_5_and_111_itm_1 <= (weight_read_addrs_7_lpi_1_dfm_2_2_0==3'b110)
          & weight_mem_run_3_for_land_lpi_1_dfm_1;
      weight_mem_run_3_for_5_and_112_itm_1 <= (weight_read_addrs_7_lpi_1_dfm_2_2_0==3'b111)
          & weight_mem_run_3_for_land_lpi_1_dfm_1;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_12_itm_1 <= ~((weight_read_addrs_7_lpi_1_dfm_2_2_0!=3'b000));
      weight_mem_run_3_for_5_and_102_itm_2 <= weight_mem_run_3_for_5_and_102_itm_1;
      weight_mem_run_3_for_5_and_103_itm_2 <= weight_mem_run_3_for_5_and_103_itm_1;
      weight_read_addrs_7_lpi_1_dfm_3_2_0 <= weight_read_addrs_7_lpi_1_dfm_2_2_0;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_5_itm_2 <= weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_5_itm_1;
      weight_mem_run_3_for_land_6_lpi_1_dfm_2 <= weight_mem_run_3_for_land_6_lpi_1_dfm_1;
      weight_mem_run_3_for_5_and_44_itm_2 <= weight_mem_run_3_for_5_and_44_itm_1;
      weight_mem_run_3_for_5_and_46_itm_2 <= weight_mem_run_3_for_5_and_46_itm_1;
      weight_mem_run_3_for_5_and_47_itm_1 <= (weight_read_addrs_5_lpi_1_dfm_2_2_0==3'b110)
          & weight_mem_run_3_for_land_6_lpi_1_dfm_1;
      weight_mem_run_3_for_5_and_48_itm_1 <= (weight_read_addrs_5_lpi_1_dfm_2_2_0==3'b111)
          & weight_mem_run_3_for_land_6_lpi_1_dfm_1;
      weight_mem_run_3_for_5_and_38_itm_1 <= (weight_read_addrs_5_lpi_1_dfm_2_2_0==3'b101)
          & weight_mem_run_3_for_land_6_lpi_1_dfm_1;
      weight_mem_run_3_for_5_and_39_itm_2 <= weight_mem_run_3_for_5_and_39_itm_1;
      weight_read_addrs_5_lpi_1_dfm_3_2_0 <= weight_read_addrs_5_lpi_1_dfm_2_2_0;
      reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_20_itm_2_cse <= weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_20_itm_1;
      weight_mem_run_3_for_5_and_162_itm_2 <= weight_mem_run_3_for_5_and_162_itm_1;
      reg_weight_mem_run_3_for_5_and_163_itm_2_cse <= weight_mem_run_3_for_5_and_163_itm_1;
      weight_mem_run_3_for_5_and_164_itm_2 <= weight_mem_run_3_for_5_and_164_itm_1;
      reg_weight_mem_run_3_for_5_and_165_itm_2_cse <= weight_mem_run_3_for_5_and_165_itm_1;
      reg_weight_mem_run_3_for_5_and_166_itm_2_cse <= weight_mem_run_3_for_5_and_166_itm_1;
      reg_weight_mem_run_3_for_5_and_167_itm_2_cse <= weight_mem_run_3_for_5_and_167_itm_1;
      reg_weight_mem_run_3_for_5_and_168_itm_2_cse <= weight_mem_run_3_for_5_and_168_itm_1;
      weight_read_addrs_3_lpi_1_dfm_3_2_0 <= weight_read_addrs_3_lpi_1_dfm_2_2_0;
      weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      weight_mem_run_3_for_5_and_156_itm_2 <= weight_mem_run_3_for_5_and_156_itm_1;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_10_itm_1 <= ~((weight_read_addrs_5_lpi_1_dfm_2_2_0!=3'b000));
      weight_mem_run_3_for_5_and_84_itm_1 <= (weight_read_addrs_5_lpi_1_dfm_2_2_0==3'b011)
          & weight_mem_run_3_for_land_6_lpi_1_dfm_1;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_3_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_10_itm_mx0w0;
      weight_mem_run_3_for_5_and_28_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_84_itm_mx0w0;
      weight_mem_run_3_for_5_and_30_itm_2 <= weight_mem_run_3_for_5_and_30_itm_1;
      weight_mem_run_3_for_5_and_31_itm_2 <= weight_mem_run_3_for_5_and_31_itm_1;
      weight_mem_run_3_for_5_and_20_itm_2 <= weight_mem_run_3_for_5_and_20_itm_1;
      weight_mem_run_3_for_5_and_22_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_94_itm_1;
      weight_mem_run_3_for_5_and_23_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_71_itm_1_1;
      reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_2_cse <= weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_1;
      weight_mem_run_3_for_5_and_8_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_72_itm_1_1;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_5 <= reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_0_1_itm_2_cse;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_5 <= reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_2_1_itm_2_cse;
      accum_vector_operator_1_for_asn_70_itm_4 <= accum_vector_operator_1_for_asn_70_itm_3;
      accum_vector_operator_1_for_asn_61_itm_4 <= accum_vector_operator_1_for_asn_61_itm_3;
      accum_vector_operator_1_for_asn_52_itm_4 <= accum_vector_operator_1_for_asn_52_itm_3;
      accum_vector_operator_1_for_asn_43_itm_4 <= accum_vector_operator_1_for_asn_43_itm_3;
      accum_vector_operator_1_for_asn_34_itm_4 <= accum_vector_operator_1_for_asn_34_itm_3;
      accum_vector_operator_1_for_asn_25_itm_4 <= accum_vector_operator_1_for_asn_25_itm_3;
      accum_vector_operator_1_for_asn_16_itm_4 <= accum_vector_operator_1_for_asn_16_itm_3;
      accum_vector_operator_1_for_asn_7_itm_4 <= accum_vector_operator_1_for_asn_7_itm_3;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_5 <= PECore_UpdateFSM_switch_lp_equal_tmp_2_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 <= 2'b00;
    end
    else if ( PECoreRun_wen & and_dcpl_41 & weight_mem_run_3_for_land_3_lpi_1_dfm_1
        ) begin
      weight_read_addrs_2_14_1_lpi_1_dfm_3_1_0 <= weight_read_addrs_2_14_1_lpi_1_dfm_2_1_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_base_weight_slc_pe_manager_base_weight_0_12_itm_2 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ mux_6_nl) & while_stage_0_6 ) begin
      pe_manager_base_weight_slc_pe_manager_base_weight_0_12_itm_2 <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_4_14_2_lpi_1_dfm_3_0 <= 1'b0;
    end
    else if ( PECoreRun_wen & weight_mem_run_3_for_land_5_lpi_1_dfm_1 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
        & while_stage_0_6 ) begin
      weight_read_addrs_4_14_2_lpi_1_dfm_3_0 <= weight_read_addrs_4_14_2_lpi_1_dfm_2_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_base_weight_slc_pe_manager_base_weight_1_0_1_itm_2 <= 2'b00;
    end
    else if ( PECoreRun_wen & mux_7_nl & while_stage_0_6 ) begin
      pe_manager_base_weight_slc_pe_manager_base_weight_1_0_1_itm_2 <= MUX_v_2_2_2(pe_manager_base_weight_slc_pe_manager_base_weight_1_0_1_itm_1,
          (weight_mem_write_arbxbar_xbar_for_empty_sva_2[7:6]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 <= 2'b00;
    end
    else if ( PECoreRun_wen & and_dcpl_41 & weight_mem_run_3_for_land_7_lpi_1_dfm_1
        ) begin
      weight_read_addrs_6_14_1_lpi_1_dfm_3_1_0 <= weight_read_addrs_6_14_1_lpi_1_dfm_2_1_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_2_itm_2_cse <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ mux_9_nl) & while_stage_0_6 ) begin
      reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_2_itm_2_cse <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ProductSum_for_asn_16_itm_5 <= 1'b0;
      ProductSum_for_asn_25_itm_5 <= 1'b0;
      ProductSum_for_asn_42_itm_5 <= 1'b0;
      ProductSum_for_asn_51_itm_5 <= 1'b0;
      ProductSum_for_asn_64_itm_5 <= 1'b0;
      ProductSum_for_asn_73_itm_5 <= 1'b0;
      ProductSum_for_asn_82_itm_5 <= 1'b0;
      ProductSum_for_asn_98_itm_5 <= 1'b0;
    end
    else if ( ProductSum_for_and_8_cse ) begin
      ProductSum_for_asn_16_itm_5 <= ProductSum_for_asn_16_itm_4;
      ProductSum_for_asn_25_itm_5 <= ProductSum_for_asn_25_itm_4;
      ProductSum_for_asn_42_itm_5 <= ProductSum_for_asn_42_itm_4;
      ProductSum_for_asn_51_itm_5 <= ProductSum_for_asn_51_itm_4;
      ProductSum_for_asn_64_itm_5 <= ProductSum_for_asn_64_itm_4;
      ProductSum_for_asn_73_itm_5 <= ProductSum_for_asn_73_itm_4;
      ProductSum_for_asn_82_itm_5 <= ProductSum_for_asn_82_itm_4;
      ProductSum_for_asn_98_itm_5 <= ProductSum_for_asn_98_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_4 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_1_read_data_and_7_enex5 ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_4 <= input_mem_banks_read_1_read_data_lpi_1_dfm_1_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_6_1_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_6_0_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_6_3_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_6_2_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_6_5_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_6_4_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_6_7_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_6_6_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_1_cse ) begin
      weight_port_read_out_data_6_1_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_2_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
      weight_port_read_out_data_6_0_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_1_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
      weight_port_read_out_data_6_3_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
      weight_port_read_out_data_6_2_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_3_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
      weight_port_read_out_data_6_5_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_6_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
      weight_port_read_out_data_6_4_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_5_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
      weight_port_read_out_data_6_7_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
      weight_port_read_out_data_6_6_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_7_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_run_3_for_land_7_lpi_1_dfm_2 <= 1'b0;
      weight_mem_run_3_for_land_5_lpi_1_dfm_2 <= 1'b0;
      weight_mem_run_3_for_land_4_lpi_1_dfm_2 <= 1'b0;
      weight_mem_run_3_for_land_3_lpi_1_dfm_2 <= 1'b0;
      weight_mem_run_3_for_land_2_lpi_1_dfm_2 <= 1'b0;
      weight_mem_run_3_for_5_and_108_itm_1 <= 1'b0;
      weight_mem_run_3_for_land_1_lpi_1_dfm_3 <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3 <= 1'b0;
      rva_in_reg_rw_sva_5 <= 1'b0;
    end
    else if ( weight_mem_run_3_for_aelse_and_1_cse ) begin
      weight_mem_run_3_for_land_7_lpi_1_dfm_2 <= weight_mem_run_3_for_land_7_lpi_1_dfm_1;
      weight_mem_run_3_for_land_5_lpi_1_dfm_2 <= weight_mem_run_3_for_land_5_lpi_1_dfm_1;
      weight_mem_run_3_for_land_4_lpi_1_dfm_2 <= weight_mem_run_3_for_land_4_lpi_1_dfm_1;
      weight_mem_run_3_for_land_3_lpi_1_dfm_2 <= weight_mem_run_3_for_land_3_lpi_1_dfm_1;
      weight_mem_run_3_for_land_2_lpi_1_dfm_2 <= weight_mem_run_3_for_land_2_lpi_1_dfm_1;
      weight_mem_run_3_for_5_and_108_itm_1 <= MUX_s_1_2_2(weight_mem_run_3_for_5_and_100_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_54_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      weight_mem_run_3_for_land_1_lpi_1_dfm_3 <= weight_mem_run_3_for_land_1_lpi_1_dfm_2;
      weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
          <= weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2;
      rva_in_reg_rw_sva_5 <= rva_in_reg_rw_sva_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_4_1_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_4_0_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_4_3_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_4_2_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_4_5_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_4_4_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_4_7_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_4_6_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_3_cse ) begin
      weight_port_read_out_data_4_1_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_2_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
      weight_port_read_out_data_4_0_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_1_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
      weight_port_read_out_data_4_3_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
      weight_port_read_out_data_4_2_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_3_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
      weight_port_read_out_data_4_5_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_6_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
      weight_port_read_out_data_4_4_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_5_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
      weight_port_read_out_data_4_7_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
      weight_port_read_out_data_4_6_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_5_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_ncse_sva_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_3_1_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_3_0_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_3_3_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_3_2_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_5_cse ) begin
      weight_port_read_out_data_3_1_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000000;
      weight_port_read_out_data_3_0_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000001;
      weight_port_read_out_data_3_3_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000002;
      weight_port_read_out_data_3_2_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_4_data_in_tmp_operator_2_for_4_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000003;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_2_1_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_2_3_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_2_2_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_2_5_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_2_4_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_2_7_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_2_6_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_7_cse ) begin
      weight_port_read_out_data_2_1_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000000;
      weight_port_read_out_data_2_3_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000006;
      weight_port_read_out_data_2_2_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000005;
      weight_port_read_out_data_2_5_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000003;
      weight_port_read_out_data_2_4_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000004;
      weight_port_read_out_data_2_7_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_pmx_sva_1;
      weight_port_read_out_data_2_6_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000002;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_1_1_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_1_0_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_1_3_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_1_2_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_1_5_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_1_4_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_1_7_sva_dfm_1 <= 8'b00000000;
      weight_port_read_out_data_1_6_sva_dfm_1 <= 8'b00000000;
    end
    else if ( weight_port_read_out_data_and_8_cse ) begin
      weight_port_read_out_data_1_1_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000000;
      weight_port_read_out_data_1_0_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000001;
      weight_port_read_out_data_1_3_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000002;
      weight_port_read_out_data_1_2_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000003;
      weight_port_read_out_data_1_5_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000004;
      weight_port_read_out_data_1_4_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000005;
      weight_port_read_out_data_1_7_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_pmx_000000;
      weight_port_read_out_data_1_6_sva_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_2_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000006;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_1_sva_dfm_1 <= 8'b00000000;
    end
    else if ( (and_1040_cse | or_dcpl_718 | or_dcpl_717) & while_stage_0_7 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & PECoreRun_wen ) begin
      weight_port_read_out_data_7_1_sva_dfm_1 <= weight_port_read_out_data_7_1_sva_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_0_sva_dfm_1 <= 8'b00000000;
    end
    else if ( (and_1044_cse | weight_mem_run_3_for_5_and_112_itm_1 | weight_mem_run_3_for_5_and_103_itm_2
        | weight_mem_run_3_for_5_and_102_itm_2 | weight_mem_run_3_for_5_and_108_itm_1)
        & while_stage_0_7 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & PECoreRun_wen ) begin
      weight_port_read_out_data_7_0_sva_dfm_1 <= weight_port_read_out_data_7_0_sva_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_5_1_sva_dfm_1 <= 8'b00000000;
    end
    else if ( (and_1048_cse | weight_mem_run_3_for_5_and_47_itm_1 | weight_mem_run_3_for_5_and_46_itm_2
        | or_dcpl_727) & while_stage_0_7 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & PECoreRun_wen ) begin
      weight_port_read_out_data_5_1_sva_dfm_1 <= weight_port_read_out_data_5_1_sva_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_5_0_sva_dfm_1 <= 8'b00000000;
    end
    else if ( (and_1048_cse | weight_mem_run_3_for_5_and_48_itm_1 | weight_mem_run_3_for_5_and_39_itm_2
        | weight_mem_run_3_for_5_and_38_itm_1 | weight_mem_run_3_for_5_and_44_itm_2)
        & while_stage_0_7 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & PECoreRun_wen ) begin
      weight_port_read_out_data_5_0_sva_dfm_1 <= weight_port_read_out_data_5_0_sva_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_11_itm_1
          <= 1'b0;
    end
    else if ( PECoreRun_wen & mux_10_nl & while_stage_0_6 ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_11_itm_1
          <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_10_itm_mx0w0,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_17_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_95_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_86_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_76_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_78_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_2 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_101_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_95_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_95_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_86_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_86_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_76_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_76_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_78_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_78_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_10_itm_1
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_84_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_79_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_80_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_71_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_72_itm_1 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_102_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_10_itm_1
          <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_10_itm_mx0w0,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_tmp,
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_84_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_84_itm_mx0w0,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_95_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_79_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_71_itm_1_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_78_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_80_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_72_itm_1_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_86_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_71_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_71_itm_1_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_72_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_72_itm_1_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_76_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_7_itm_1
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_60_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_62_itm_1 <= 1'b0;
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse <= 3'b000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_44_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_47_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_48_itm_1 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_105_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_7_itm_1
          <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_for_crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_tmp,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_44_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_60_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_20_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_46_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_62_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_6_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse <= crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_44_itm_2 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_44_itm_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_and_49_tmp, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_47_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_15_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_48_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_16_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_44_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_6_itm_2
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_46_itm_2 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_108_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_6_itm_2
          <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_6_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_46_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_46_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_54_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_56_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_44_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_34_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_35_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_2_itm_2
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_14_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_15_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_17_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_3 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_19_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_20_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_3
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_itm_2 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_54_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_54_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_56_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_56_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_44_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_44_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_34_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_34_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_35_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_35_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_2_itm_2
          <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_2_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_14_itm_2 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_4;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_15_itm_2 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_4;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_itm_2 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_4;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_17_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_17_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_3 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_2;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_19_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_19_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_20_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_20_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_3
          <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_2;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_itm_2 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_8 <= 8'b00000000;
    end
    else if ( (weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
        | weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
        | weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
        | weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
        | weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
        | weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
        | weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2
        | weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2)
        & mux_512_nl & fsm_output & while_stage_0_7 & PECoreRun_wen & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        ) begin
      BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_8 <= BitsToType_spec_PE_Weight_WordType_return_data_2_0_lpi_1_dfm_9;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_1_for_3_result_val_Marshall_64U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1
          <= 8'b00000000;
    end
    else if ( PECoreRun_wen & mux_12_nl & while_stage_0_6 ) begin
      weight_mem_banks_load_store_1_for_3_result_val_Marshall_64U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1
          <= MUX_v_8_2_2((weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[7:0]), weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_24_nl,
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_1_for_5_result_val_Marshall_64U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1
          <= 8'b00000000;
    end
    else if ( PECoreRun_wen & mux_13_nl & while_stage_0_6 ) begin
      weight_mem_banks_load_store_1_for_5_result_val_Marshall_64U_2_for_1_marshaller_AddField_ac_int_8_false_8_15_else_bits_slc_BitsToType_spec_PE_Weight_WordType_2_marshaller_glob_1_7_0_1_itm_1
          <= MUX_v_8_2_2((weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[7:0]), weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_40_nl,
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_lpi_1_dfm_1_63_8 <= 56'b00000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & (~(or_dcpl_606 | (~ weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2)
        | (~ fsm_output))) & mux_14_nl ) begin
      weight_mem_banks_read_1_read_data_lpi_1_dfm_1_63_8 <= weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d[63:8];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_7_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & (~(or_dcpl_606 | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_2)
        | (~ fsm_output))) & mux_15_nl ) begin
      weight_mem_banks_read_1_read_data_7_lpi_1_dfm_1 <= weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_0_1_itm_2_cse
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(PECore_RunFSM_switch_lp_equal_tmp_1_2 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3))
        & while_stage_0_5 ) begin
      reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_0_1_itm_2_cse
          <= PECore_PushOutput_PECore_PushOutput_if_and_svs_st_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(PECore_UpdateFSM_switch_lp_equal_tmp_2_3 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3))
        & while_stage_0_5 ) begin
      reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse
          <= PECore_RunMac_PECore_RunMac_if_and_svs_st_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_2_1_itm_2_cse
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(ProductSum_for_asn_16_itm_3 & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3))
        & while_stage_0_5 ) begin
      reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_2_1_itm_2_cse
          <= PECore_RunScale_PECore_RunScale_if_and_1_svs_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_3_1_itm_2_cse
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ mux_16_nl) & while_stage_0_5 ) begin
      reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_3_1_itm_2_cse
          <= PECore_RunScale_PECore_RunScale_if_and_1_svs_st_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_2
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ ProductSum_for_asn_42_itm_3) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
        & while_stage_0_5 ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_2
          <= weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_2
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ ProductSum_for_asn_51_itm_3) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
        & while_stage_0_5 ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_2
          <= weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_0_14_4_lpi_1_dfm_1_4 <= 11'b00000000000;
    end
    else if ( weight_read_addrs_and_7_enex5 ) begin
      weight_read_addrs_0_14_4_lpi_1_dfm_1_4 <= weight_read_addrs_0_14_4_lpi_1_dfm_1_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_2
          <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_69 & (~ ProductSum_for_asn_64_itm_3) ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_2
          <= weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_slc_weight_read_addrs_0_3_0_3_23_itm_1 <= 1'b0;
    end
    else if ( PECoreRun_wen & weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_1
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
        & while_stage_0_5 & (~ ProductSum_for_asn_73_itm_3) ) begin
      weight_read_addrs_slc_weight_read_addrs_0_3_0_3_23_itm_1 <= weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_2
          <= 1'b0;
    end
    else if ( PECoreRun_wen & and_dcpl_69 & (~ ProductSum_for_asn_73_itm_3) ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_2
          <= weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_11_1
          <= 11'b00000000000;
    end
    else if ( weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_11_1
          <= MUX_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
          (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
          (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
          (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
          {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_2 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_1
          , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_0});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_0
          <= 1'b0;
    end
    else if ( weight_mem_read_arbxbar_xbar_1_for_3_and_8_cse ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_6_itm_1_0
          <= MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, (weight_read_addrs_1_lpi_1_dfm_1[3]),
          (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]), (weight_read_addrs_3_lpi_1_dfm_1[3]),
          (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]), (weight_read_addrs_5_lpi_1_dfm_1[3]),
          (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]), (weight_read_addrs_7_lpi_1_dfm_1[3]),
          {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_2 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_1
          , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_30_0});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_11_1
          <= 11'b00000000000;
    end
    else if ( weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_11_1
          <= MUX_v_11_8_2(weight_read_addrs_0_14_4_lpi_1_dfm_1_3, (weight_read_addrs_1_lpi_1_dfm_1[14:4]),
          (weight_read_addrs_2_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_3_lpi_1_dfm_1[14:4]),
          (weight_read_addrs_4_14_2_lpi_1_dfm_1[12:2]), (weight_read_addrs_5_lpi_1_dfm_1[14:4]),
          (weight_read_addrs_6_14_1_lpi_1_dfm_1[13:3]), (weight_read_addrs_7_lpi_1_dfm_1[14:4]),
          {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_2 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_1
          , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_0});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_0
          <= 1'b0;
    end
    else if ( weight_mem_read_arbxbar_xbar_1_for_3_and_10_cse ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_weight_mem_read_arbxbar_xbar_1_for_3_and_7_itm_1_0
          <= MUX_s_1_8_2(weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, (weight_read_addrs_1_lpi_1_dfm_1[3]),
          (weight_read_addrs_2_14_1_lpi_1_dfm_1[2]), (weight_read_addrs_3_lpi_1_dfm_1[3]),
          (weight_read_addrs_4_14_2_lpi_1_dfm_1[1]), (weight_read_addrs_5_lpi_1_dfm_1[3]),
          (weight_read_addrs_6_14_1_lpi_1_dfm_1[2]), (weight_read_addrs_7_lpi_1_dfm_1[3]),
          {weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_2 , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_1
          , weight_mem_read_arbxbar_xbar_1_for_3_if_1_conc_32_0});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
          <= 1'b0;
      weight_mem_run_3_for_land_4_lpi_1_dfm_1 <= 1'b0;
      weight_mem_run_3_for_land_2_lpi_1_dfm_1 <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_run_3_for_land_3_lpi_1_dfm_1 <= 1'b0;
      weight_mem_run_3_for_land_5_lpi_1_dfm_1 <= 1'b0;
      weight_mem_run_3_for_land_7_lpi_1_dfm_1 <= 1'b0;
      weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= 1'b0;
      weight_mem_run_3_for_land_1_lpi_1_dfm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2 <= 1'b0;
      rva_in_reg_rw_sva_4 <= 1'b0;
    end
    else if ( while_if_and_10_cse ) begin
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3;
      weight_mem_run_3_for_land_4_lpi_1_dfm_1 <= weight_mem_run_3_for_land_4_lpi_1_dfm_1_1;
      weight_mem_run_3_for_land_2_lpi_1_dfm_1 <= weight_mem_run_3_for_land_2_lpi_1_dfm_1_1;
      weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp;
      weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp;
      weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp;
      weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp;
      weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp;
      weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp;
      weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp;
      weight_mem_run_3_for_land_3_lpi_1_dfm_1 <= PECore_RunFSM_switch_lp_equal_tmp_1_2
          & or_196_cse;
      weight_mem_run_3_for_land_5_lpi_1_dfm_1 <= PECore_RunFSM_switch_lp_equal_tmp_1_2
          & or_162_cse;
      weight_mem_run_3_for_land_7_lpi_1_dfm_1 <= PECore_RunFSM_switch_lp_equal_tmp_1_2
          & or_186_cse;
      weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
          <= weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp;
      weight_mem_run_3_for_land_1_lpi_1_dfm_2 <= weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1;
      rva_in_reg_rw_sva_4 <= rva_in_reg_rw_sva_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_7_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_7_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_7_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_7_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_7_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_7_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_50_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_7_1_sva <= weight_mem_read_arbxbar_arbiters_next_7_1_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_7_2_sva <= weight_mem_read_arbxbar_arbiters_next_7_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_7_3_sva <= weight_mem_read_arbxbar_arbiters_next_7_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_7_4_sva <= weight_mem_read_arbxbar_arbiters_next_7_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_7_5_sva <= weight_mem_read_arbxbar_arbiters_next_7_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_7_6_sva <= weight_mem_read_arbxbar_arbiters_next_7_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_6_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_6_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_6_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_6_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_6_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_6_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_56_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_6_1_sva <= weight_mem_read_arbxbar_arbiters_next_6_1_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_6_2_sva <= weight_mem_read_arbxbar_arbiters_next_6_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_6_3_sva <= weight_mem_read_arbxbar_arbiters_next_6_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_6_4_sva <= weight_mem_read_arbxbar_arbiters_next_6_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_6_5_sva <= weight_mem_read_arbxbar_arbiters_next_6_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_6_6_sva <= weight_mem_read_arbxbar_arbiters_next_6_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_5_1_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_cse & (and_dcpl_69 | Arbiter_8U_Roundrobin_pick_and_1_cse)
        & or_dcpl_16 ) begin
      weight_mem_read_arbxbar_arbiters_next_5_1_sva <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_41_mx1w0,
          Arbiter_8U_Roundrobin_pick_1_mux_396_itm_1, Arbiter_8U_Roundrobin_pick_and_1_cse);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_5_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_5_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_5_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_5_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_5_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_62_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_5_2_sva <= weight_mem_read_arbxbar_arbiters_next_5_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_5_3_sva <= weight_mem_read_arbxbar_arbiters_next_5_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_5_4_sva <= weight_mem_read_arbxbar_arbiters_next_5_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_5_5_sva <= weight_mem_read_arbxbar_arbiters_next_5_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_5_6_sva <= weight_mem_read_arbxbar_arbiters_next_5_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_4_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_4_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_4_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_4_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_4_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_4_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_67_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_4_1_sva <= weight_mem_read_arbxbar_arbiters_next_4_1_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_4_2_sva <= weight_mem_read_arbxbar_arbiters_next_4_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_4_3_sva <= weight_mem_read_arbxbar_arbiters_next_4_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_4_4_sva <= weight_mem_read_arbxbar_arbiters_next_4_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_4_5_sva <= weight_mem_read_arbxbar_arbiters_next_4_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_4_6_sva <= weight_mem_read_arbxbar_arbiters_next_4_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_3_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_3_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_3_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_3_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_3_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_3_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_73_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_3_1_sva <= weight_mem_read_arbxbar_arbiters_next_3_1_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_3_2_sva <= weight_mem_read_arbxbar_arbiters_next_3_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_3_3_sva <= weight_mem_read_arbxbar_arbiters_next_3_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_3_4_sva <= weight_mem_read_arbxbar_arbiters_next_3_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_3_5_sva <= weight_mem_read_arbxbar_arbiters_next_3_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_3_6_sva <= weight_mem_read_arbxbar_arbiters_next_3_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_2_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_2_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_2_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_2_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_2_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_2_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_79_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_2_1_sva <= weight_mem_read_arbxbar_arbiters_next_2_1_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_2_2_sva <= weight_mem_read_arbxbar_arbiters_next_2_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_2_3_sva <= weight_mem_read_arbxbar_arbiters_next_2_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_2_4_sva <= weight_mem_read_arbxbar_arbiters_next_2_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_2_5_sva <= weight_mem_read_arbxbar_arbiters_next_2_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_2_6_sva <= weight_mem_read_arbxbar_arbiters_next_2_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_1_1_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_1_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_1_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_1_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_1_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_1_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_85_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_1_1_sva <= weight_mem_read_arbxbar_arbiters_next_1_1_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_1_2_sva <= weight_mem_read_arbxbar_arbiters_next_1_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_1_3_sva <= weight_mem_read_arbxbar_arbiters_next_1_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_1_4_sva <= weight_mem_read_arbxbar_arbiters_next_1_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_1_5_sva <= weight_mem_read_arbxbar_arbiters_next_1_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_1_6_sva <= weight_mem_read_arbxbar_arbiters_next_1_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_0_1_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_cse & (and_dcpl_69 | Arbiter_8U_Roundrobin_pick_and_13_cse)
        & or_dcpl_21 ) begin
      weight_mem_read_arbxbar_arbiters_next_0_1_sva <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_6_mx1w0,
          Arbiter_8U_Roundrobin_pick_1_mux_31_itm_1, Arbiter_8U_Roundrobin_pick_and_13_cse);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_arbiters_next_0_2_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_0_3_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_0_4_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_0_5_sva <= 1'b1;
      weight_mem_read_arbxbar_arbiters_next_0_6_sva <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_arbiters_next_and_91_cse ) begin
      weight_mem_read_arbxbar_arbiters_next_0_2_sva <= weight_mem_read_arbxbar_arbiters_next_0_2_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_0_3_sva <= weight_mem_read_arbxbar_arbiters_next_0_3_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_0_4_sva <= weight_mem_read_arbxbar_arbiters_next_0_4_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_0_5_sva <= weight_mem_read_arbxbar_arbiters_next_0_5_sva_mx1;
      weight_mem_read_arbxbar_arbiters_next_0_6_sva <= weight_mem_read_arbxbar_arbiters_next_0_6_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_base_weight_sva <= 15'b000000000000000;
    end
    else if ( (~ mux_514_nl) & fsm_output & while_stage_0_5 & PECoreRun_wen ) begin
      pe_manager_base_weight_sva <= pe_manager_base_weight_sva_mx2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_0_14_4_lpi_1_dfm_1_3 <= 11'b00000000000;
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3 <= 1'b0;
    end
    else if ( weight_read_addrs_and_9_cse ) begin
      weight_read_addrs_0_14_4_lpi_1_dfm_1_3 <= MUX_v_11_2_2(PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_6_nl,
          weight_read_addrs_0_14_4_lpi_1_dfm_1_2, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
      weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3 <= MUX_s_1_2_2((weight_read_addrs_0_3_0_lpi_1_dfm_4[3]),
          (weight_read_addrs_0_3_0_lpi_1_dfm_1_2[3]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_1
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4]))
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
        & while_stage_0_4 ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_4_1_itm_1
          <= weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[4];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_1
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5]))
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
        & while_stage_0_4 ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_5_1_itm_1
          <= weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[5];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_7_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_24_enex5 ) begin
      weight_write_data_data_0_7_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_7_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_6_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_25_enex5 ) begin
      weight_write_data_data_0_6_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_6_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_5_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_26_enex5 ) begin
      weight_write_data_data_0_5_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_5_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_4_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_27_enex5 ) begin
      weight_write_data_data_0_4_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_4_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_3_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_28_enex5 ) begin
      weight_write_data_data_0_3_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_3_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_2_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_29_enex5 ) begin
      weight_write_data_data_0_2_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_2_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_1_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_30_enex5 ) begin
      weight_write_data_data_0_1_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_1_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_0_lpi_1_dfm_1_3_2 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_31_enex5 ) begin
      weight_write_data_data_0_0_lpi_1_dfm_1_3_2 <= weight_write_data_data_0_0_lpi_1_dfm_1_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_addrs_lpi_1_dfm_1_3_14_3 <= 12'b000000000000;
    end
    else if ( weight_write_addrs_and_enex5 ) begin
      weight_write_addrs_lpi_1_dfm_1_3_14_3 <= weight_write_addrs_lpi_1_dfm_1_2[14:3];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_1
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6]))
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
        & while_stage_0_4 ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_1
          <= weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[6];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_1
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7]))
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
        & while_stage_0_4 ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_7_1_itm_1
          <= weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[7];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_3
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_4
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_5
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_6
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_0
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_1
          <= 1'b0;
      weight_read_addrs_1_lpi_1_dfm_1 <= 15'b000000000000000;
      weight_read_addrs_2_14_1_lpi_1_dfm_1 <= 14'b00000000000000;
      weight_read_addrs_3_lpi_1_dfm_1 <= 15'b000000000000000;
      weight_read_addrs_4_14_2_lpi_1_dfm_1 <= 13'b0000000000000;
      weight_read_addrs_5_lpi_1_dfm_1 <= 15'b000000000000000;
      weight_read_addrs_6_14_1_lpi_1_dfm_1 <= 14'b00000000000000;
      weight_read_addrs_7_lpi_1_dfm_1 <= 15'b000000000000000;
      Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_0 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_5_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_2 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_3 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_0 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_5_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_2 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_3 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_0 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_5_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_1_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_2_cse <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_3_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_0 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_5_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_2 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_3 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_0 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_5_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_2 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_3 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_6_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_0 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_5_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_4_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_2 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_3 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_0_2_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_0 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_5_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_1 <= 1'b0;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_cse <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_2 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_3 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_1_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_6 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_0 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_5 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_4 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_2 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_3 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_576_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_496_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_423_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_350_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_277_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_204_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_131_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_57_itm_1 <= 1'b0;
      accum_vector_operator_1_for_asn_70_itm_2 <= 1'b0;
      accum_vector_operator_1_for_asn_61_itm_2 <= 1'b0;
      accum_vector_operator_1_for_asn_34_itm_2 <= 1'b0;
      accum_vector_operator_1_for_asn_25_itm_2 <= 1'b0;
      accum_vector_operator_1_for_asn_16_itm_2 <= 1'b0;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_cse
        ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_3
          <= MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1,
          nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3_mx1,
          and_149_cse);
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_4
          <= MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1,
          nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4_mx1,
          and_149_cse);
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_5
          <= MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1,
          nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5_mx1,
          and_149_cse);
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_6
          <= MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1,
          nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6_mx1,
          and_149_cse);
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_0
          <= MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_0_1,
          nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0_mx1,
          and_149_cse);
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_2
          <= MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1,
          nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2_mx1,
          and_149_cse);
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_1_1_1
          <= MUX_s_1_2_2(nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1,
          nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1_mx1,
          and_149_cse);
      weight_read_addrs_1_lpi_1_dfm_1 <= weight_read_addrs_1_lpi_1_dfm_1_1;
      weight_read_addrs_2_14_1_lpi_1_dfm_1 <= weight_read_addrs_2_14_1_lpi_1_dfm_1_1;
      weight_read_addrs_3_lpi_1_dfm_1 <= weight_read_addrs_3_lpi_1_dfm_1_1;
      weight_read_addrs_4_14_2_lpi_1_dfm_1 <= weight_read_addrs_4_14_2_lpi_1_dfm_1_1;
      weight_read_addrs_5_lpi_1_dfm_1 <= weight_read_addrs_5_lpi_1_dfm_1_1;
      weight_read_addrs_6_14_1_lpi_1_dfm_1 <= weight_read_addrs_6_14_1_lpi_1_dfm_1_1;
      weight_read_addrs_7_lpi_1_dfm_1 <= weight_read_addrs_7_lpi_1_dfm_1_1;
      Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_2;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1 <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_0_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_5_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_5_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_4_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_2 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_2_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_3 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_3_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
      Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_2;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_6_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1 <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_0_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_5_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_5_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_4_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_4_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_2 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_2_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_3 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_3_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_9;
      Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_2;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_6_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_5_1 <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_10;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_0_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_10;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_5_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_5_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_1_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_4_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_4_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_2_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_2_1;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_6_lpi_1_dfm_1_3_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_3_1;
      Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_2;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_6_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_4_1 <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_0_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_5_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_5_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_4_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_4_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_2 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_2_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_5_lpi_1_dfm_1_3 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_3_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_11;
      Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_2;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_6_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_3_1 <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_12;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_0_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_12;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_5_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_5_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_1_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_12;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_4_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_4_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_2 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_2_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_12;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_4_lpi_1_dfm_1_3 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_3_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_12;
      Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_2;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_6_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_2_1 <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_13;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_0_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_13;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_5_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_5_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_13;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_4_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_4_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_2 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_2_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_13;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_3_lpi_1_dfm_1_3 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_3_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_13;
      Arbiter_8U_Roundrobin_pick_return_1_0_2_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_return_1_0_2_lpi_1_dfm_2;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_6_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1_1 <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_14;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_0_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_14;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_5_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_5_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_14;
      reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_4_cse <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_4_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_2 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_2_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_14;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_2_lpi_1_dfm_1_3 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_3_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_14;
      Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_1_1 <= Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_2;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_6 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1;
      Arbiter_8U_Roundrobin_pick_1_unequal_tmp_1 <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_15;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_0 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_0_1
          & Arbiter_8U_Roundrobin_pick_1_unequal_tmp_15;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_5 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_4 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_2 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1;
      Arbiter_8U_Roundrobin_pick_return_1_7_1_1_lpi_1_dfm_1_3 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1;
      Arbiter_8U_Roundrobin_pick_1_mux_576_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_1_if_1_not_185,
          weight_mem_read_arbxbar_arbiters_next_7_7_sva_mx0, and_100_cse);
      Arbiter_8U_Roundrobin_pick_1_mux_496_itm_1 <= MUX_s_1_2_2((~ weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1),
          weight_mem_read_arbxbar_arbiters_next_6_7_sva_mx0, and_dcpl_533);
      Arbiter_8U_Roundrobin_pick_1_mux_423_itm_1 <= MUX_s_1_2_2((~ weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1),
          weight_mem_read_arbxbar_arbiters_next_5_7_sva_mx0, and_114_cse);
      Arbiter_8U_Roundrobin_pick_1_mux_350_itm_1 <= MUX_s_1_2_2((~ weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1),
          weight_mem_read_arbxbar_arbiters_next_4_7_sva_mx0, and_dcpl_547);
      Arbiter_8U_Roundrobin_pick_1_mux_277_itm_1 <= MUX_s_1_2_2((~ weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1),
          weight_mem_read_arbxbar_arbiters_next_3_7_sva_mx0, and_dcpl_554);
      Arbiter_8U_Roundrobin_pick_1_mux_204_itm_1 <= MUX_s_1_2_2((~ weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1),
          weight_mem_read_arbxbar_arbiters_next_2_7_sva_mx0, and_dcpl_561);
      Arbiter_8U_Roundrobin_pick_1_mux_131_itm_1 <= MUX_s_1_2_2((~ weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1),
          weight_mem_read_arbxbar_arbiters_next_1_7_sva_mx0, and_dcpl_568);
      Arbiter_8U_Roundrobin_pick_1_mux_57_itm_1 <= MUX_s_1_2_2((~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1),
          weight_mem_read_arbxbar_arbiters_next_0_7_sva_mx0, and_149_cse);
      accum_vector_operator_1_for_asn_70_itm_2 <= accum_vector_operator_1_for_asn_70_itm_1;
      accum_vector_operator_1_for_asn_61_itm_2 <= PECore_DecodeAxiWrite_switch_lp_equal_tmp_1_2;
      accum_vector_operator_1_for_asn_34_itm_2 <= PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_2;
      accum_vector_operator_1_for_asn_25_itm_2 <= PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_2;
      accum_vector_operator_1_for_asn_16_itm_2 <= PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunFSM_switch_lp_equal_tmp_1_2 <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
          <= 1'b0;
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_178_itm_1 <= 1'b0;
      weight_mem_run_3_for_land_1_lpi_1_dfm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1 <= 1'b0;
      rva_in_reg_rw_sva_3 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_3 <= 1'b0;
    end
    else if ( PECore_RunFSM_switch_lp_and_cse ) begin
      PECore_RunFSM_switch_lp_equal_tmp_1_2 <= MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2,
          (weight_mem_write_arbxbar_xbar_for_lshift_tmp[0]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2;
      pe_manager_base_weight_slc_pe_manager_base_weight_2_0_178_itm_1 <= MUX_s_1_2_2((pe_manager_base_weight_sva_mx1_3_0[1]),
          reg_rva_in_reg_rw_sva_2_cse, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
      weight_mem_run_3_for_land_1_lpi_1_dfm_1 <= weight_mem_run_3_for_land_1_lpi_1_dfm_1_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1_1;
      rva_in_reg_rw_sva_3 <= reg_rva_in_reg_rw_sva_2_cse;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_3 <= MUX_s_1_2_2(PECore_DecodeAxiRead_switch_lp_equal_tmp_1_1,
          (weight_mem_write_arbxbar_xbar_for_lshift_tmp[1]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0
          <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_396_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_395_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_394_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_393_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_392_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_391_itm_1 <= 1'b0;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_13_cse
        ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_0_1;
      Arbiter_8U_Roundrobin_pick_1_mux_396_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_395_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_394_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_393_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_392_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_6_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_391_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_6_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_6_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_3
          <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_323_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_322_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_321_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_320_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_319_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_318_itm_1 <= 1'b0;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_14_cse
        ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_0_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_2
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_2_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_3
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_3_1;
      Arbiter_8U_Roundrobin_pick_1_mux_323_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_1_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_322_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_321_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_320_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_319_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_5_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_318_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_6_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_5_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_3
          <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_250_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_249_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_248_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_247_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_246_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_245_itm_1 <= 1'b0;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_18_cse
        ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_0_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_1_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_2
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_2_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_3
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_3_1;
      Arbiter_8U_Roundrobin_pick_1_mux_250_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_1_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_249_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_248_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_247_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_246_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_4_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_245_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_6_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_4_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_3
          <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_177_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_176_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_175_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_174_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_173_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_172_itm_1 <= 1'b0;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_22_cse
        ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_0_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_2
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_2_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_3
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_3_1;
      Arbiter_8U_Roundrobin_pick_1_mux_177_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_1_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_176_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_175_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_174_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_173_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_3_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_172_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_6_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_3_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_0
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_3
          <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_104_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_103_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_102_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_101_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_100_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_99_itm_1 <= 1'b0;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_26_cse
        ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_0_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_2
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_2_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_3
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_3_1;
      Arbiter_8U_Roundrobin_pick_1_mux_104_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_1_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_103_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_102_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_101_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_100_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_2_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_99_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_6_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_2_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_mux_542_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_541_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_540_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_539_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_538_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_537_itm_1 <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_0
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_3
          <= 1'b0;
    end
    else if ( Arbiter_8U_Roundrobin_pick_1_and_15_cse ) begin
      Arbiter_8U_Roundrobin_pick_1_mux_542_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1
          | Arbiter_8U_Roundrobin_pick_1_if_1_not_185;
      Arbiter_8U_Roundrobin_pick_1_mux_541_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
          | Arbiter_8U_Roundrobin_pick_1_if_1_not_185;
      Arbiter_8U_Roundrobin_pick_1_mux_540_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
          | Arbiter_8U_Roundrobin_pick_1_if_1_not_185;
      Arbiter_8U_Roundrobin_pick_1_mux_539_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
          | Arbiter_8U_Roundrobin_pick_1_if_1_not_185;
      Arbiter_8U_Roundrobin_pick_1_mux_538_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_sva_1
          | Arbiter_8U_Roundrobin_pick_1_if_1_not_185;
      Arbiter_8U_Roundrobin_pick_1_mux_537_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_6_1
          | Arbiter_8U_Roundrobin_pick_1_if_1_not_185;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_0_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_2
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_2_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_3
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_3_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1 <= 8'b00000000;
      weight_mem_write_arbxbar_xbar_for_empty_sva_1 <= 8'b00000000;
      crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1 <= 3'b000;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_and_15_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_and_8_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_and_45_itm_1 <= 1'b0;
      rva_in_reg_rw_sva_st_3 <= 1'b0;
    end
    else if ( weight_mem_read_arbxbar_xbar_requests_transpose_and_14_cse ) begin
      weight_mem_read_arbxbar_xbar_requests_transpose_0_sva_1 <= weight_mem_read_arbxbar_xbar_for_1_lshift_tmp;
      weight_mem_write_arbxbar_xbar_for_empty_sva_1 <= weight_mem_write_arbxbar_xbar_for_lshift_tmp;
      crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_and_15_itm_1 <= (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1_1==3'b101)
          & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_and_8_itm_1 <= (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1_1==3'b110)
          & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_and_45_itm_1 <= (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1_1==3'b011)
          & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1_1;
      rva_in_reg_rw_sva_st_3 <= reg_rva_in_reg_rw_sva_2_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1 <= 1'b1;
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1 <= 1'b1;
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_itm_1 <= 1'b1;
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_itm_1 <= 1'b1;
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_itm_1 <= 1'b1;
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_itm_1 <= 1'b1;
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1 <= 1'b1;
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1 <= 1'b1;
    end
    else if ( Arbiter_8U_Roundrobin_pick_and_cse ) begin
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_576_itm_1, and_dcpl_525);
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_496_itm_1, and_dcpl_525);
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_423_itm_1, and_dcpl_525);
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_350_itm_1, and_dcpl_525);
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_277_itm_1, and_dcpl_525);
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_204_itm_1, and_dcpl_525);
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_131_itm_1, and_dcpl_525);
      Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_itm_1 <= MUX_s_1_2_2(Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_nl,
          Arbiter_8U_Roundrobin_pick_1_mux_57_itm_1, and_dcpl_525);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_mux_469_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_468_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_467_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_466_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_465_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_464_itm_1 <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_0
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3
          <= 1'b0;
    end
    else if ( Arbiter_8U_Roundrobin_pick_1_and_22_cse ) begin
      Arbiter_8U_Roundrobin_pick_1_mux_469_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_468_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_467_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_466_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_465_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_7_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_464_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_6_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_0_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_2
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_2_1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_3
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_3_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_mux_31_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_30_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_29_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_28_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_27_itm_1 <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_mux_26_itm_1 <= 1'b0;
    end
    else if ( Arbiter_8U_Roundrobin_pick_1_and_64_cse ) begin
      Arbiter_8U_Roundrobin_pick_1_mux_31_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
          | nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_30_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_29_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_28_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_27_itm_1 <= Arbiter_8U_Roundrobin_pick_1_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_1_if_1_if_for_or_1_cse_1_sva_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
      Arbiter_8U_Roundrobin_pick_1_mux_26_itm_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1
          | (~ weight_mem_read_arbxbar_xbar_1_for_3_1_operator_4_false_3_operator_4_false_3_nand_mdf_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_base_weight_sva_dfm_3_1 <= 15'b000000000000000;
    end
    else if ( PECore_RunFSM_switch_lp_and_cse & ((~ while_stage_0_5) | while_and_1126_itm_1)
        ) begin
      pe_manager_base_weight_sva_dfm_3_1 <= MUX_v_15_2_2(pe_manager_base_weight_sva_mx2,
          PEManager_15U_PEManagerWrite_slc_rva_in_reg_data_30_16_itm_1, while_and_1126_itm_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_7_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_32_enex5 ) begin
      weight_write_data_data_0_7_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_7_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_6_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_33_enex5 ) begin
      weight_write_data_data_0_6_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_6_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_5_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_34_enex5 ) begin
      weight_write_data_data_0_5_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_5_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_4_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_35_enex5 ) begin
      weight_write_data_data_0_4_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_4_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_3_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_36_enex5 ) begin
      weight_write_data_data_0_3_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_3_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_2_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_37_enex5 ) begin
      weight_write_data_data_0_2_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_2_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_1_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_38_enex5 ) begin
      weight_write_data_data_0_1_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_1_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_data_data_0_0_lpi_1_dfm_1_2_6 <= 8'b00000000;
    end
    else if ( weight_write_data_data_and_39_enex5 ) begin
      weight_write_data_data_0_0_lpi_1_dfm_1_2_6 <= weight_write_data_data_0_0_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_write_addrs_lpi_1_dfm_1_2 <= 15'b000000000000000;
    end
    else if ( weight_write_addrs_and_2_enex5 ) begin
      weight_write_addrs_lpi_1_dfm_1_2 <= pe_manager_base_input_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiWrite_switch_lp_equal_tmp_1_2 <= 1'b0;
      reg_rva_in_reg_rw_sva_2_cse <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2 <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
          <= 1'b0;
      while_and_1126_itm_1 <= 1'b0;
    end
    else if ( PECore_DecodeAxiWrite_switch_lp_and_2_cse ) begin
      PECore_DecodeAxiWrite_switch_lp_equal_tmp_1_2 <= MUX_s_1_2_2(accum_vector_data_6_sva_1_load_mx0w1,
          PECore_DecodeAxiWrite_switch_lp_equal_tmp_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
      reg_rva_in_reg_rw_sva_2_cse <= reg_rva_in_reg_rw_sva_st_1_1_cse;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2 <= MUX_s_1_2_2(PECore_RunFSM_switch_lp_equal_tmp_1_mx0w1,
          PECore_DecodeAxiRead_switch_lp_equal_tmp_2, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2
          <= while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
      while_and_1126_itm_1 <= PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_1_1
          & PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_nor_1_cse_1
          & reg_rva_in_reg_rw_sva_st_1_1_cse & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_0_3_0_lpi_1_dfm_1_2 <= 4'b0000;
    end
    else if ( weight_read_addrs_and_28_enex5 ) begin
      weight_read_addrs_0_3_0_lpi_1_dfm_1_2 <= weight_read_addrs_0_3_0_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PEManager_15U_GetWeightAddr_else_acc_3_1 <= 11'b00000000000;
    end
    else if ( PECoreRun_wen & and_dcpl_207 ) begin
      PEManager_15U_GetWeightAddr_else_acc_3_1 <= PEManager_15U_GetWeightAddr_else_acc_4_cmp_z;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      state_2_1_sva <= 2'b00;
      pe_config_is_zero_first_sva <= 1'b0;
    end
    else if ( state_and_cse ) begin
      state_2_1_sva <= state_mux_1_cse;
      pe_config_is_zero_first_sva <= pe_config_is_zero_first_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      state_0_sva <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ or_dcpl_616) ) begin
      state_0_sva <= PECore_UpdateFSM_next_state_0_lpi_1_dfm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_config_manager_counter_sva <= 4'b0000;
    end
    else if ( (((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7:2]==6'b000000) & nor_907_cse
        & nor_909_cse & nor_910_cse & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])
        & (~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19])))
        & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & rva_in_PopNB_mioi_return_rsc_z_mxwt
        & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17:16]==2'b00) & and_dcpl_211)
        | and_1065_cse) & PECoreRun_wen ) begin
      pe_config_manager_counter_sva <= MUX_v_4_2_2(pe_config_manager_counter_sva_dfm_3_1,
          PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_and_nl,
          and_601_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_config_num_manager_sva <= 4'b0001;
      pe_config_num_output_sva <= 8'b00000001;
    end
    else if ( pe_config_num_manager_and_cse ) begin
      pe_config_num_manager_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[35:32];
      pe_config_num_output_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[47:40];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_in_reg_rw_sva_st_1_1_cse <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
          <= 1'b0;
      PECore_DecodeAxiWrite_switch_lp_nor_tmp_1 <= 1'b0;
      state_2_1_sva_dfm_1 <= 2'b00;
      PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_1_1 <= 1'b0;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4
          <= 8'b00000000;
      input_write_req_valid_lpi_1_dfm_1_1 <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_6_cse ) begin
      reg_rva_in_reg_rw_sva_st_1_1_cse <= rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
          <= rva_in_PopNB_mioi_return_rsc_z_mxwt;
      PECore_DecodeAxiWrite_switch_lp_nor_tmp_1 <= PECore_DecodeAxiWrite_switch_lp_nor_tmp_1_1;
      state_2_1_sva_dfm_1 <= MUX_v_2_2_2(PECore_UpdateFSM_switch_lp_and_1_nl, state_mux_1_cse,
          rva_in_PopNB_mioi_return_rsc_z_mxwt);
      PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_1_1 <= and_321_cse;
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_1_11_4
          <= rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7:0];
      input_write_req_valid_lpi_1_dfm_1_1 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0
          & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_UpdateFSM_switch_lp_equal_tmp_5_1 <= 1'b0;
      PECore_UpdateFSM_switch_lp_and_7_itm_1 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_1 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_3_1 <= 1'b0;
      PECore_UpdateFSM_switch_lp_nor_7_itm_1 <= 1'b0;
      PECore_RunFSM_switch_lp_nor_tmp_1 <= 1'b0;
    end
    else if ( PECore_UpdateFSM_switch_lp_and_9_cse ) begin
      PECore_UpdateFSM_switch_lp_equal_tmp_5_1 <= PECore_PushOutput_PECore_PushOutput_if_and_svs_1;
      PECore_UpdateFSM_switch_lp_and_7_itm_1 <= PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_1_cse_1;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_1 <= PECore_UpdateFSM_switch_lp_equal_tmp_6;
      PECore_UpdateFSM_switch_lp_equal_tmp_3_1 <= PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_1_cse_1;
      PECore_UpdateFSM_switch_lp_nor_7_itm_1 <= ~(PECore_RunScale_PECore_RunScale_if_and_1_svs_1
          | PECore_UpdateFSM_switch_lp_nor_tmp_1);
      PECore_RunFSM_switch_lp_nor_tmp_1 <= ~(PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_1_cse_1
          | PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_1_cse_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva
          <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(or_dcpl_632 | or_dcpl_616)) ) begin
      PECore_RunFSM_case_0_Connections_InBlocking_spec_StreamType_Connections_SYN_PORT_PopNB_return_sva
          <= input_port_PopNB_mioi_return_rsc_z_mxwt;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_config_input_counter_sva <= 8'b00000000;
    end
    else if ( or_1491_cse & mux_515_nl & weight_mem_read_arbxbar_arbiters_next_and_cse
        & while_stage_0_3 ) begin
      pe_config_input_counter_sva <= pe_config_input_counter_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_config_output_counter_sva <= 8'b00000000;
    end
    else if ( or_1491_cse & mux_516_nl & and_dcpl_759 & PECoreRun_wen ) begin
      pe_config_output_counter_sva <= pe_config_output_counter_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      operator_8_false_acc_sdt_sva_1 <= 9'b000000000;
    end
    else if ( pe_config_UpdateManagerCounter_if_if_and_enex5 ) begin
      operator_8_false_acc_sdt_sva_1 <= nl_operator_8_false_acc_sdt_sva_1[8:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiWrite_switch_lp_equal_tmp_2 <= 1'b0;
      PECore_DecodeAxiWrite_switch_lp_equal_tmp_1 <= 1'b0;
    end
    else if ( PECore_DecodeAxiWrite_switch_lp_and_cse ) begin
      PECore_DecodeAxiWrite_switch_lp_equal_tmp_2 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0;
      PECore_DecodeAxiWrite_switch_lp_equal_tmp_1 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_reg_data_19_0_sva <= 20'b00000000000000000000;
      act_port_reg_data_51_32_sva <= 20'b00000000000000000000;
      act_port_reg_data_83_64_sva <= 20'b00000000000000000000;
      act_port_reg_data_115_96_sva <= 20'b00000000000000000000;
      act_port_reg_data_147_128_sva <= 20'b00000000000000000000;
      act_port_reg_data_179_160_sva <= 20'b00000000000000000000;
      act_port_reg_data_211_192_sva <= 20'b00000000000000000000;
      act_port_reg_data_243_224_sva <= 20'b00000000000000000000;
    end
    else if ( and_1098_cse ) begin
      act_port_reg_data_19_0_sva <= act_port_reg_data_19_0_sva_mx1;
      act_port_reg_data_51_32_sva <= act_port_reg_data_51_32_sva_mx1;
      act_port_reg_data_83_64_sva <= act_port_reg_data_83_64_sva_mx1;
      act_port_reg_data_115_96_sva <= act_port_reg_data_115_96_sva_mx1;
      act_port_reg_data_147_128_sva <= act_port_reg_data_147_128_sva_mx1;
      act_port_reg_data_179_160_sva <= act_port_reg_data_179_160_sva_mx1;
      act_port_reg_data_211_192_sva <= act_port_reg_data_211_192_sva_mx1;
      act_port_reg_data_243_224_sva <= act_port_reg_data_243_224_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_7_sva <= 23'b00000000000000000000000;
      accum_vector_data_0_sva <= 23'b00000000000000000000000;
      accum_vector_data_6_sva <= 23'b00000000000000000000000;
      accum_vector_data_1_sva <= 23'b00000000000000000000000;
      accum_vector_data_5_sva <= 23'b00000000000000000000000;
      accum_vector_data_2_sva <= 23'b00000000000000000000000;
      accum_vector_data_4_sva <= 23'b00000000000000000000000;
      accum_vector_data_3_sva <= 23'b00000000000000000000000;
    end
    else if ( accum_vector_data_and_40_cse ) begin
      accum_vector_data_7_sva <= nl_accum_vector_data_7_sva[22:0];
      accum_vector_data_0_sva <= nl_accum_vector_data_0_sva[22:0];
      accum_vector_data_6_sva <= nl_accum_vector_data_6_sva[22:0];
      accum_vector_data_1_sva <= nl_accum_vector_data_1_sva[22:0];
      accum_vector_data_5_sva <= nl_accum_vector_data_5_sva[22:0];
      accum_vector_data_2_sva <= nl_accum_vector_data_2_sva[22:0];
      accum_vector_data_4_sva <= nl_accum_vector_data_4_sva[22:0];
      accum_vector_data_3_sva <= nl_accum_vector_data_3_sva[22:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_8 <= 1'b0;
      accum_vector_operator_1_for_asn_64_itm_7 <= 1'b0;
      accum_vector_operator_1_for_asn_55_itm_7 <= 1'b0;
      accum_vector_operator_1_for_asn_46_itm_7 <= 1'b0;
      accum_vector_operator_1_for_asn_37_itm_7 <= 1'b0;
      accum_vector_operator_1_for_asn_28_itm_7 <= 1'b0;
      accum_vector_operator_1_for_asn_22_itm_7 <= 1'b0;
      accum_vector_operator_1_for_asn_10_itm_7 <= 1'b0;
      accum_vector_operator_1_for_asn_1_itm_7 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_8 <= 1'b0;
    end
    else if ( PECore_RunScale_if_and_cse ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_8 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_7;
      accum_vector_operator_1_for_asn_64_itm_7 <= accum_vector_operator_1_for_asn_70_itm_6;
      accum_vector_operator_1_for_asn_55_itm_7 <= accum_vector_operator_1_for_asn_61_itm_6;
      accum_vector_operator_1_for_asn_46_itm_7 <= accum_vector_operator_1_for_asn_52_itm_6;
      accum_vector_operator_1_for_asn_37_itm_7 <= accum_vector_operator_1_for_asn_43_itm_6;
      accum_vector_operator_1_for_asn_28_itm_7 <= accum_vector_operator_1_for_asn_34_itm_6;
      accum_vector_operator_1_for_asn_22_itm_7 <= accum_vector_operator_1_for_asn_25_itm_6;
      accum_vector_operator_1_for_asn_10_itm_7 <= accum_vector_operator_1_for_asn_16_itm_6;
      accum_vector_operator_1_for_asn_1_itm_7 <= accum_vector_operator_1_for_asn_7_itm_6;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_8 <= PECore_UpdateFSM_switch_lp_equal_tmp_2_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_25_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_31_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_27_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_26_itm_1
          <= 8'b00000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_cse ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_25_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[15:8]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_122_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_31_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[63:56]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_125_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_27_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[31:24]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_128_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_26_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[23:16]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_76_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_41_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_47_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_45_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_43_itm_1
          <= 8'b00000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_1_cse ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_41_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[15:8]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_108_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_47_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[63:56]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_111_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_45_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[47:40]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_112_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_43_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[31:24]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_114_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_4_itm_1
          <= 8'b00000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_2_cse ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[7:0]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_130_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_4_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[39:32]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_134_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_7_sva_dfm_1_1 <= 8'b00000000;
    end
    else if ( (and_1129_cse | or_dcpl_718 | weight_mem_run_3_for_5_and_156_itm_2)
        & while_stage_0_7 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & PECoreRun_wen ) begin
      weight_port_read_out_data_7_7_sva_dfm_1_1 <= weight_port_read_out_data_7_7_sva_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_6_sva_dfm_1_1 <= 8'b00000000;
    end
    else if ( (and_1129_cse | or_dcpl_751 | weight_mem_run_3_for_5_and_156_itm_2)
        & while_stage_0_7 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & PECoreRun_wen ) begin
      weight_port_read_out_data_7_6_sva_dfm_1_1 <= weight_port_read_out_data_7_6_sva_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_5_sva_dfm_1_1 <= 8'b00000000;
      weight_port_read_out_data_7_3_sva_dfm_1_1 <= 8'b00000000;
    end
    else if ( and_1138_cse ) begin
      weight_port_read_out_data_7_5_sva_dfm_1_1 <= weight_port_read_out_data_7_5_sva_dfm_2;
      weight_port_read_out_data_7_3_sva_dfm_1_1 <= weight_port_read_out_data_7_3_sva_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_4_sva_dfm_1_1 <= 8'b00000000;
    end
    else if ( (and_1129_cse | or_dcpl_751 | weight_mem_run_3_for_5_and_108_itm_1)
        & while_stage_0_7 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & PECoreRun_wen ) begin
      weight_port_read_out_data_7_4_sva_dfm_1_1 <= weight_port_read_out_data_7_4_sva_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_7_2_sva_dfm_1_1 <= 8'b00000000;
    end
    else if ( (and_1044_cse | or_dcpl_751 | or_dcpl_717) & while_stage_0_7 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & PECoreRun_wen ) begin
      weight_port_read_out_data_7_2_sva_dfm_1_1 <= weight_port_read_out_data_7_2_sva_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_5_7_sva_dfm_1_1 <= 8'b00000000;
    end
    else if ( (and_1048_cse | weight_mem_run_3_for_5_and_39_itm_2 | weight_mem_run_3_for_5_and_38_itm_1
        | or_dcpl_727) & while_stage_0_7 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & PECoreRun_wen ) begin
      weight_port_read_out_data_5_7_sva_dfm_1_1 <= weight_port_read_out_data_5_7_sva_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_5_6_sva_dfm_1_1 <= 8'b00000000;
    end
    else if ( (((xor_7_cse | weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_10_itm_1)
        & weight_mem_run_3_for_land_6_lpi_1_dfm_2) | or_dcpl_779 | weight_mem_run_3_for_5_and_84_itm_1)
        & while_stage_0_7 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & PECoreRun_wen ) begin
      weight_port_read_out_data_5_6_sva_dfm_1_1 <= weight_port_read_out_data_5_6_sva_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_5_5_sva_dfm_1_1 <= 8'b00000000;
      weight_port_read_out_data_5_3_sva_dfm_1_1 <= 8'b00000000;
    end
    else if ( and_1162_cse ) begin
      weight_port_read_out_data_5_5_sva_dfm_1_1 <= weight_port_read_out_data_5_5_sva_dfm_2;
      weight_port_read_out_data_5_3_sva_dfm_1_1 <= weight_port_read_out_data_5_3_sva_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_5_4_sva_dfm_1_1 <= 8'b00000000;
      weight_port_read_out_data_5_2_sva_dfm_1_1 <= 8'b00000000;
    end
    else if ( and_1166_cse ) begin
      weight_port_read_out_data_5_4_sva_dfm_1_1 <= weight_port_read_out_data_5_4_sva_dfm_2;
      weight_port_read_out_data_5_2_sva_dfm_1_1 <= weight_port_read_out_data_5_2_sva_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_3_7_sva_dfm_1_1 <= 8'b00000000;
    end
    else if ( (and_1177_cse | or_dcpl_801 | weight_mem_run_3_for_5_and_28_itm_1)
        & while_stage_0_7 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & PECoreRun_wen ) begin
      weight_port_read_out_data_3_7_sva_dfm_1_1 <= weight_port_read_out_data_3_7_sva_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_3_6_sva_dfm_1_1 <= 8'b00000000;
    end
    else if ( (and_1177_cse | weight_mem_run_3_for_5_and_23_itm_1 | weight_mem_run_3_for_5_and_22_itm_1
        | weight_mem_run_3_for_5_and_20_itm_2) & while_stage_0_7 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & PECoreRun_wen ) begin
      weight_port_read_out_data_3_6_sva_dfm_1_1 <= weight_port_read_out_data_3_6_sva_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_3_5_sva_dfm_1_1 <= 8'b00000000;
    end
    else if ( (((xor_13_cse | reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_2_cse)
        & weight_mem_run_3_for_land_4_lpi_1_dfm_2) | or_dcpl_801 | weight_mem_run_3_for_5_and_20_itm_2)
        & while_stage_0_7 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & PECoreRun_wen ) begin
      weight_port_read_out_data_3_5_sva_dfm_1_1 <= weight_port_read_out_data_3_5_sva_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_3_4_sva_dfm_1_1 <= 8'b00000000;
    end
    else if ( ((((((weight_read_addrs_3_lpi_1_dfm_3_2_0[2:1]!=2'b00)) ^ (weight_read_addrs_3_lpi_1_dfm_3_2_0[0]))
        | reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_2_cse) & weight_mem_run_3_for_land_4_lpi_1_dfm_2)
        | weight_mem_run_3_for_5_and_30_itm_2 | weight_mem_run_3_for_5_and_20_itm_2
        | weight_mem_run_3_for_5_and_8_itm_1) & while_stage_0_7 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5)
        & PECoreRun_wen ) begin
      weight_port_read_out_data_3_4_sva_dfm_1_1 <= weight_port_read_out_data_3_4_sva_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_7_lpi_1_dfm_2_2_0 <= 3'b000;
      weight_mem_run_3_for_land_lpi_1_dfm_1 <= 1'b0;
      weight_read_addrs_5_lpi_1_dfm_2_2_0 <= 3'b000;
      weight_mem_run_3_for_land_6_lpi_1_dfm_1 <= 1'b0;
      weight_read_addrs_3_lpi_1_dfm_2_2_0 <= 3'b000;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_13_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_103_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_102_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_46_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_44_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_5_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_39_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_168_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_167_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_166_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_165_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_164_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_163_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_162_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_20_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_156_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_31_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_30_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_and_20_itm_1 <= 1'b0;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_1 <= 1'b0;
      accum_vector_operator_1_for_asn_70_itm_3 <= 1'b0;
      accum_vector_operator_1_for_asn_61_itm_3 <= 1'b0;
      accum_vector_operator_1_for_asn_52_itm_3 <= 1'b0;
      accum_vector_operator_1_for_asn_43_itm_3 <= 1'b0;
      accum_vector_operator_1_for_asn_34_itm_3 <= 1'b0;
      accum_vector_operator_1_for_asn_25_itm_3 <= 1'b0;
      accum_vector_operator_1_for_asn_16_itm_3 <= 1'b0;
      accum_vector_operator_1_for_asn_7_itm_3 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_4 <= 1'b0;
    end
    else if ( weight_read_addrs_and_19_cse ) begin
      weight_read_addrs_7_lpi_1_dfm_2_2_0 <= weight_read_addrs_7_lpi_1_dfm_1[2:0];
      weight_mem_run_3_for_land_lpi_1_dfm_1 <= weight_mem_run_3_for_land_lpi_1_dfm_1_1;
      weight_read_addrs_5_lpi_1_dfm_2_2_0 <= weight_read_addrs_5_lpi_1_dfm_1[2:0];
      weight_mem_run_3_for_land_6_lpi_1_dfm_1 <= weight_mem_run_3_for_land_6_lpi_1_dfm_1_1;
      weight_read_addrs_3_lpi_1_dfm_2_2_0 <= weight_read_addrs_3_lpi_1_dfm_1[2:0];
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_13_itm_1 <= ~((weight_read_addrs_7_lpi_1_dfm_1[2:0]!=3'b000));
      weight_mem_run_3_for_5_and_103_itm_1 <= (weight_read_addrs_7_lpi_1_dfm_1[2:0]==3'b110)
          & weight_mem_run_3_for_land_lpi_1_dfm_1_1;
      weight_mem_run_3_for_5_and_102_itm_1 <= (weight_read_addrs_7_lpi_1_dfm_1[2:0]==3'b101)
          & weight_mem_run_3_for_land_lpi_1_dfm_1_1;
      weight_mem_run_3_for_5_and_46_itm_1 <= (weight_read_addrs_5_lpi_1_dfm_1[2:0]==3'b101)
          & weight_mem_run_3_for_land_6_lpi_1_dfm_1_1;
      weight_mem_run_3_for_5_and_44_itm_1 <= (weight_read_addrs_5_lpi_1_dfm_1[2:0]==3'b011)
          & weight_mem_run_3_for_land_6_lpi_1_dfm_1_1;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_5_itm_1 <= ~((weight_read_addrs_5_lpi_1_dfm_1[2:0]!=3'b000));
      weight_mem_run_3_for_5_and_39_itm_1 <= (weight_read_addrs_5_lpi_1_dfm_1[2:0]==3'b110)
          & weight_mem_run_3_for_land_6_lpi_1_dfm_1_1;
      weight_mem_run_3_for_5_and_168_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_1;
      weight_mem_run_3_for_5_and_167_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_1;
      weight_mem_run_3_for_5_and_166_itm_1 <= (pe_manager_base_weight_sva[2:0]==3'b101)
          & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      weight_mem_run_3_for_5_and_165_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_9_itm_1;
      weight_mem_run_3_for_5_and_164_itm_1 <= pe_manager_base_weight_slc_pe_manager_base_weight_2_0_178_itm_1
          & (pe_manager_base_weight_sva[0]) & (~ (pe_manager_base_weight_sva[2]))
          & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      weight_mem_run_3_for_5_and_163_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_7_itm_1;
      weight_mem_run_3_for_5_and_162_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_6_itm_1;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_20_itm_1 <= ~((pe_manager_base_weight_sva[2:0]!=3'b000));
      weight_mem_run_3_for_5_and_156_itm_1 <= (weight_read_addrs_7_lpi_1_dfm_1[2:0]==3'b011)
          & weight_mem_run_3_for_land_lpi_1_dfm_1_1;
      weight_mem_run_3_for_5_and_31_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_95_itm_mx0w0;
      weight_mem_run_3_for_5_and_30_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_mx0w0;
      weight_mem_run_3_for_5_and_20_itm_1 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_1_1;
      weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_1_itm_1 <= ~((weight_read_addrs_3_lpi_1_dfm_1[2:0]!=3'b000));
      accum_vector_operator_1_for_asn_70_itm_3 <= accum_vector_operator_1_for_asn_70_itm_2;
      accum_vector_operator_1_for_asn_61_itm_3 <= accum_vector_operator_1_for_asn_61_itm_2;
      accum_vector_operator_1_for_asn_52_itm_3 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_3;
      accum_vector_operator_1_for_asn_43_itm_3 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_3;
      accum_vector_operator_1_for_asn_34_itm_3 <= accum_vector_operator_1_for_asn_34_itm_2;
      accum_vector_operator_1_for_asn_25_itm_3 <= accum_vector_operator_1_for_asn_25_itm_2;
      accum_vector_operator_1_for_asn_16_itm_3 <= accum_vector_operator_1_for_asn_16_itm_2;
      accum_vector_operator_1_for_asn_7_itm_3 <= input_read_req_valid_lpi_1_dfm_1_3;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_4 <= PECore_UpdateFSM_switch_lp_equal_tmp_2_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
        & while_stage_0_6 & fsm_output & ((~ weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp)
        | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
        | (~ while_stage_0_5)) ) begin
      weight_mem_banks_read_1_read_data_6_lpi_1_dfm_1_1 <= weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
        & while_stage_0_6 & fsm_output & ((~ weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp)
        | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
        | (~ while_stage_0_5)) ) begin
      weight_mem_banks_read_1_read_data_5_lpi_1_dfm_1_1 <= weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
        & while_stage_0_6 & fsm_output & ((~ weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp)
        | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
        | (~ while_stage_0_5)) ) begin
      weight_mem_banks_read_1_read_data_4_lpi_1_dfm_1_1 <= weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
        & while_stage_0_6 & fsm_output & ((~ weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp)
        | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
        | (~ while_stage_0_5)) ) begin
      weight_mem_banks_read_1_read_data_3_lpi_1_dfm_1_1 <= weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
        & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
        & while_stage_0_6 & fsm_output & ((~ weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp)
        | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
        | (~ while_stage_0_5)) ) begin
      weight_mem_banks_read_1_read_data_2_lpi_1_dfm_1_1 <= weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_read_1_read_data_1_lpi_1_dfm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( PECoreRun_wen & (~(or_tmp_382 | (~ while_stage_0_6) | (~ fsm_output)))
        & ((~ weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp)
        | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
        | (~ while_stage_0_5)) ) begin
      weight_mem_banks_read_1_read_data_1_lpi_1_dfm_1 <= weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2
          <= 1'b0;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3
          <= 1'b0;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_30_cse
        ) begin
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_6_mx1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_0_mx1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_5_mx1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_1_mx1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_4_mx1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_2_mx1;
      nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_lpi_1_dfm_16_3_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_0_14_4_lpi_1_dfm_1_2 <= 11'b00000000000;
    end
    else if ( weight_read_addrs_and_29_enex5 ) begin
      weight_read_addrs_0_14_4_lpi_1_dfm_1_2 <= weight_read_addrs_0_14_4_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs
          <= 1'b0;
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112 <= 1'b0;
    end
    else if ( operator_15_false_1_and_cse ) begin
      weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs
          <= Arbiter_8U_Roundrobin_pick_1_unequal_tmp_8;
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_112_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(and_149_cse | or_dcpl_13)) ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_7_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(and_dcpl_568 | or_dcpl_13)) ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_22_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(and_dcpl_561 | or_dcpl_13)) ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_37_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(and_dcpl_554 | or_dcpl_13)) ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_52_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(and_dcpl_547 | or_dcpl_13)) ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_67_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(and_114_cse | or_dcpl_13)) ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_82_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(and_dcpl_533 | or_dcpl_13)) ) begin
      Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97 <= Arbiter_8U_Roundrobin_pick_1_if_1_and_tmp_97_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PEManager_15U_PEManagerWrite_slc_rva_in_reg_data_30_16_itm_1 <= 15'b000000000000000;
    end
    else if ( PEManager_15U_PEManagerWrite_and_enex5 ) begin
      PEManager_15U_PEManagerWrite_slc_rva_in_reg_data_30_16_itm_1 <= rva_in_reg_data_sva_1[30:16];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_num_input_sva <= 8'b00000001;
      pe_manager_base_bias_sva <= 15'b000000000000000;
    end
    else if ( pe_manager_num_input_and_cse ) begin
      pe_manager_num_input_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[15:8];
      pe_manager_base_bias_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[46:32];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_config_is_valid_sva <= 1'b0;
      pe_config_is_cluster_sva <= 1'b0;
      pe_config_is_bias_sva <= 1'b0;
    end
    else if ( pe_config_is_valid_and_cse ) begin
      pe_config_is_valid_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[0];
      pe_config_is_cluster_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[16];
      pe_config_is_bias_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[24];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_zero_active_sva <= 1'b0;
    end
    else if ( PECoreRun_wen & and_321_cse & (~ PECore_DecodeAxiWrite_switch_lp_or_5_cse_1)
        & (~ or_dcpl_627) ) begin
      pe_manager_zero_active_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_config_output_counter_sva_dfm_1 <= 8'b00000000;
    end
    else if ( (((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5:2]==4'b0000) & nor_922_cse
        & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[13:8]==6'b000000) & nor_910_cse
        & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1:0]==2'b01)) | PECore_DecodeAxiWrite_switch_lp_equal_tmp_1
        | PECore_DecodeAxiWrite_switch_lp_equal_tmp_2 | PECore_DecodeAxiWrite_switch_lp_nor_tmp_1
        | (~(reg_rva_in_reg_rw_sva_st_1_1_cse & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1
        & while_stage_0_3))) & rva_in_PopNB_mioi_return_rsc_z_mxwt & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:16]==4'b0100)
        & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt & rva_in_reg_rw_and_6_cse ) begin
      pe_config_output_counter_sva_dfm_1 <= MUX_v_8_2_2(8'b00000000, pe_config_output_counter_sva_mx1,
          PECore_DecodeAxiWrite_case_4_switch_lp_or_cse_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_config_input_counter_sva_dfm_1 <= 8'b00000000;
    end
    else if ( and_1217_tmp ) begin
      pe_config_input_counter_sva_dfm_1 <= MUX_v_8_2_2(PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_20_nl,
          PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_and_1_nl,
          rva_in_PopNB_mioi_data_rw_rsc_z_mxwt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_if_mux_19_itm_1 <= 1'b0;
      weight_read_addrs_0_3_0_lpi_1_dfm_1_1 <= 4'b0000;
      weight_write_data_data_0_7_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_write_data_data_0_6_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_write_data_data_0_5_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_write_data_data_0_4_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_write_data_data_0_3_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_write_data_data_0_2_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_write_data_data_0_1_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_write_data_data_0_0_lpi_1_dfm_1_1 <= 8'b00000000;
      weight_read_addrs_0_14_4_lpi_1_dfm_1_1 <= 11'b00000000000;
    end
    else if ( while_if_and_14_cse ) begin
      while_if_mux_19_itm_1 <= MUX_s_1_2_2(pe_config_is_zero_first_sva_mx1, PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_mux_19_nl,
          rva_in_PopNB_mioi_data_rw_rsc_z_mxwt);
      weight_read_addrs_0_3_0_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3:0])
          & ({{3{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & (signext_4_1(~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt));
      weight_write_data_data_0_7_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[63:56])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_6_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[55:48])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_5_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[47:40])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_4_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[39:32])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_3_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[31:24])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_2_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[23:16])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_1_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[15:8])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_write_data_data_0_0_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[7:0])
          & ({{7{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & ({{7{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
      weight_read_addrs_0_14_4_lpi_1_dfm_1_1 <= (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[14:4])
          & ({{10{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
          & (signext_11_1(~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_7 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_6
        | PECore_RunMac_PECore_RunMac_if_and_svs_st_6)) & while_stage_0_8 ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_7 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_st_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_st_1_4 <= 1'b0;
      rva_in_reg_rw_sva_st_4 <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_7_cse ) begin
      rva_in_reg_rw_sva_st_1_4 <= pe_manager_base_weight_slc_pe_manager_base_weight_2_0_178_itm_1;
      rva_in_reg_rw_sva_st_4 <= rva_in_reg_rw_sva_st_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_rw_sva_st_1_6 <= 1'b0;
      rva_in_reg_rw_sva_st_6 <= 1'b0;
    end
    else if ( rva_in_reg_rw_and_8_cse ) begin
      rva_in_reg_rw_sva_st_1_6 <= rva_in_reg_rw_sva_st_1_5;
      rva_in_reg_rw_sva_st_6 <= rva_in_reg_rw_sva_st_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1
          <= 4'b0000;
    end
    else if ( PECoreRun_wen & and_dcpl_242 ) begin
      while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1
          <= rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:16];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ProductSum_for_asn_16_itm_4 <= 1'b0;
      ProductSum_for_asn_25_itm_4 <= 1'b0;
      ProductSum_for_asn_42_itm_4 <= 1'b0;
      ProductSum_for_asn_51_itm_4 <= 1'b0;
      ProductSum_for_asn_64_itm_4 <= 1'b0;
      ProductSum_for_asn_73_itm_4 <= 1'b0;
      ProductSum_for_asn_82_itm_4 <= 1'b0;
      ProductSum_for_asn_98_itm_4 <= 1'b0;
    end
    else if ( ProductSum_for_and_16_cse ) begin
      ProductSum_for_asn_16_itm_4 <= ProductSum_for_asn_16_itm_3;
      ProductSum_for_asn_25_itm_4 <= ProductSum_for_asn_25_itm_3;
      ProductSum_for_asn_42_itm_4 <= ProductSum_for_asn_42_itm_3;
      ProductSum_for_asn_51_itm_4 <= ProductSum_for_asn_51_itm_3;
      ProductSum_for_asn_64_itm_4 <= ProductSum_for_asn_64_itm_3;
      ProductSum_for_asn_73_itm_4 <= ProductSum_for_asn_73_itm_3;
      ProductSum_for_asn_82_itm_4 <= ProductSum_for_asn_82_itm_3;
      ProductSum_for_asn_98_itm_4 <= ProductSum_for_asn_98_itm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_base_weight_slc_pe_manager_base_weight_1_0_1_itm_1 <= 2'b00;
    end
    else if ( PECoreRun_wen & or_162_cse & and_dcpl_248 ) begin
      pe_manager_base_weight_slc_pe_manager_base_weight_1_0_1_itm_1 <= pe_manager_base_weight_sva[1:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_95_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_86_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_78_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_76_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_1 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_122_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_95_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_95_itm_mx0w0,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_86_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_mx0w0,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_1_nl,
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_78_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_mx0w0,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_and_8_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_76_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_1_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_and_7_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_70_itm_mx0w0,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_and_45_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_1_1,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_and_9_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2 <= 3'b000;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_46_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_44_itm_1 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_124_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_7_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_and_16_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2 <= MUX_v_3_2_2((weight_read_addrs_1_lpi_1_dfm_1[2:0]),
          crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_46_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_14_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_and_15_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_44_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_4_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_and_5_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_6_itm_1
          <= 1'b0;
    end
    else if ( PECoreRun_wen & weight_mem_read_arbxbar_xbar_1_for_3_8_for_2_or_cse
        & and_dcpl_248 ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_6_itm_1
          <= ~((weight_read_addrs_1_lpi_1_dfm_1[2:0]!=3'b000));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_56_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_2_itm_1
          <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_2 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_2
          <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_72_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_56_itm_1 <= (pe_manager_base_weight_sva[2:0]==3'b011)
          & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_2_itm_1
          <= ~(pe_manager_base_weight_slc_pe_manager_base_weight_2_0_95_itm_1 | (pe_manager_base_weight_sva[1:0]!=2'b00));
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_2 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_18_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_2
          <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_54_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_44_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_35_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_34_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_20_itm_1 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_19_itm_1 <= 1'b0;
    end
    else if ( crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_73_cse ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_54_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_6_itm_1,
          ProductSum_for_asn_73_itm_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_44_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_28_nl,
          ProductSum_for_asn_64_itm_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_35_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_35_nl,
          ProductSum_for_asn_51_itm_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_34_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_34_nl,
          ProductSum_for_asn_42_itm_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_nl,
          ProductSum_for_asn_25_itm_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_nl,
          ProductSum_for_asn_16_itm_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_20_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_12_itm_1,
          PECore_UpdateFSM_switch_lp_equal_tmp_2_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_19_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_11_itm_1,
          PECore_RunFSM_switch_lp_equal_tmp_1_2, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_1 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_1 <=
          1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_1
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_1
          <= 1'b0;
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_1
          <= 1'b0;
    end
    else if ( input_mem_banks_read_read_data_and_9_cse ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_0_itm_1 <=
          input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0[0];
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_8_itm_1 <=
          input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0[8];
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_16_itm_1
          <= input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0[16];
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_31_itm_1
          <= input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0[31];
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_24_itm_1
          <= input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0[24];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_1
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_26_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_1
          <= input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0[7:1];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_1
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_27_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_1
          <= input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0[15:9];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_1
          <= 7'b0000000;
    end
    else if ( input_mem_banks_read_read_data_and_28_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_1
          <= input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0[23:17];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_1
          <= 6'b000000;
    end
    else if ( input_mem_banks_read_read_data_and_29_enex5 ) begin
      input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_1
          <= input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0[30:25];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_8
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_8
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_6
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_6
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_4_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_8
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_7;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_8
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_7;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_6
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_5;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_6
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_3 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_1_read_data_and_3_enex5 ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_3 <= input_mem_banks_read_1_read_data_lpi_1_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_6_14_1_lpi_1_dfm_2_1_0 <= 2'b00;
    end
    else if ( PECoreRun_wen & or_186_cse & and_dcpl_248 ) begin
      weight_read_addrs_6_14_1_lpi_1_dfm_2_1_0 <= weight_read_addrs_6_14_1_lpi_1_dfm_1[1:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_4_14_2_lpi_1_dfm_2_0 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ mux_31_nl) & while_stage_0_5 ) begin
      weight_read_addrs_4_14_2_lpi_1_dfm_2_0 <= MUX_s_1_2_2((weight_read_addrs_4_14_2_lpi_1_dfm_1[0]),
          weight_read_addrs_0_3_0_lpi_1_dfm_1_3_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_read_addrs_2_14_1_lpi_1_dfm_2_1_0 <= 2'b00;
    end
    else if ( PECoreRun_wen & or_196_cse & and_dcpl_248 ) begin
      weight_read_addrs_2_14_1_lpi_1_dfm_2_1_0 <= weight_read_addrs_2_14_1_lpi_1_dfm_1[1:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_read_req_valid_lpi_1_dfm_1_8 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6 <= 1'b0;
      rva_out_reg_data_39_36_sva_dfm_4_3_rsp_0 <= 1'b0;
      rva_out_reg_data_39_36_sva_dfm_4_3_rsp_1 <= 1'b0;
      rva_out_reg_data_39_36_sva_dfm_4_3_rsp_2 <= 2'b00;
      rva_out_reg_data_46_40_sva_dfm_4_3_rsp_0 <= 3'b000;
    end
    else if ( input_read_req_valid_and_1_cse ) begin
      input_read_req_valid_lpi_1_dfm_1_8 <= input_read_req_valid_lpi_1_dfm_1_7;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_6 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5;
      rva_out_reg_data_39_36_sva_dfm_4_3_rsp_0 <= rva_out_reg_data_39_36_sva_dfm_4_2_3;
      rva_out_reg_data_39_36_sva_dfm_4_3_rsp_1 <= rva_out_reg_data_39_36_sva_dfm_4_2_2;
      rva_out_reg_data_39_36_sva_dfm_4_3_rsp_2 <= rva_out_reg_data_39_36_sva_dfm_4_2_1_0;
      rva_out_reg_data_46_40_sva_dfm_4_3_rsp_0 <= rva_out_reg_data_46_40_sva_dfm_4_2_6_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_8 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_8 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_7 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_8 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_7_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_8 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_7;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_8 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_7;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_7 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_1_6;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_8 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_6 <= 6'b000000;
    end
    else if ( rva_out_reg_data_and_86_enex5 ) begin
      rva_out_reg_data_30_25_sva_dfm_6 <= rva_out_reg_data_30_25_sva_dfm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_23_17_sva_dfm_6 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_87_enex5 ) begin
      rva_out_reg_data_23_17_sva_dfm_6 <= rva_out_reg_data_23_17_sva_dfm_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_8 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_88_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_8 <= rva_out_reg_data_15_9_sva_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_4_3 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_89_enex5 ) begin
      rva_out_reg_data_35_32_sva_dfm_4_3 <= rva_out_reg_data_35_32_sva_dfm_4_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_56_sva_dfm_4_3 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_90_enex5 ) begin
      rva_out_reg_data_62_56_sva_dfm_4_3 <= rva_out_reg_data_62_56_sva_dfm_4_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_7_sva_5 <= 23'b00000000000000000000000;
    end
    else if ( mux_538_nl & and_dcpl_885 & PECoreRun_wen & or_dcpl_824 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8)
        ) begin
      accum_vector_data_7_sva_5 <= accum_vector_data_7_sva_5_mx1w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_7_sva_4 <= 23'b00000000000000000000000;
    end
    else if ( or_dcpl_824 & while_stage_0_10 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8)
        & PECoreRun_wen ) begin
      accum_vector_data_7_sva_4 <= accum_vector_data_7_sva_4_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_6_sva_5 <= 23'b00000000000000000000000;
    end
    else if ( mux_546_nl & and_dcpl_885 & PECoreRun_wen & or_dcpl_826 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8)
        ) begin
      accum_vector_data_6_sva_5 <= accum_vector_data_6_sva_5_mx1w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_6_sva_4 <= 23'b00000000000000000000000;
    end
    else if ( or_dcpl_826 & while_stage_0_10 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8)
        & PECoreRun_wen ) begin
      accum_vector_data_6_sva_4 <= accum_vector_data_6_sva_4_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_5_sva_5 <= 23'b00000000000000000000000;
    end
    else if ( or_dcpl_828 & while_stage_0_10 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8)
        & PECoreRun_wen ) begin
      accum_vector_data_5_sva_5 <= accum_vector_data_5_sva_5_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_5_sva_4 <= 23'b00000000000000000000000;
    end
    else if ( mux_554_nl & and_dcpl_885 & PECoreRun_wen & or_dcpl_828 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8)
        ) begin
      accum_vector_data_5_sva_4 <= accum_vector_data_5_sva_4_mx1w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_4_sva_5 <= 23'b00000000000000000000000;
      accum_vector_data_4_sva_4 <= 23'b00000000000000000000000;
    end
    else if ( and_1250_cse ) begin
      accum_vector_data_4_sva_5 <= accum_vector_data_4_sva_5_mx1w0;
      accum_vector_data_4_sva_4 <= accum_vector_data_4_sva_4_mx1w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_3_sva_5 <= 23'b00000000000000000000000;
      accum_vector_data_3_sva_4 <= 23'b00000000000000000000000;
    end
    else if ( and_1262_cse ) begin
      accum_vector_data_3_sva_5 <= accum_vector_data_3_sva_5_mx1w0;
      accum_vector_data_3_sva_4 <= accum_vector_data_3_sva_4_mx1w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_2_sva_6 <= 23'b00000000000000000000000;
      accum_vector_data_2_sva_5 <= 23'b00000000000000000000000;
      accum_vector_data_2_sva_4 <= 23'b00000000000000000000000;
    end
    else if ( and_1274_cse ) begin
      accum_vector_data_2_sva_6 <= accum_vector_data_2_sva_6_mx1w0;
      accum_vector_data_2_sva_5 <= accum_vector_data_2_sva_5_mx1w0;
      accum_vector_data_2_sva_4 <= accum_vector_data_2_sva_4_mx1w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_1_sva_5 <= 23'b00000000000000000000000;
      accum_vector_data_1_sva_4 <= 23'b00000000000000000000000;
    end
    else if ( and_1292_cse ) begin
      accum_vector_data_1_sva_5 <= accum_vector_data_1_sva_5_mx1w0;
      accum_vector_data_1_sva_4 <= accum_vector_data_1_sva_4_mx1w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_0_sva_5 <= 23'b00000000000000000000000;
      accum_vector_data_0_sva_4 <= 23'b00000000000000000000000;
    end
    else if ( and_1304_cse ) begin
      accum_vector_data_0_sva_5 <= accum_vector_data_0_sva_5_mx1w0;
      accum_vector_data_0_sva_4 <= accum_vector_data_0_sva_4_mx1w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_2_sva_7 <= 23'b00000000000000000000000;
    end
    else if ( and_dcpl_964 & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7)
        & or_tmp_864 & PECoreRun_wen ) begin
      accum_vector_data_2_sva_7 <= MUX_v_23_2_2(23'b00000000000000000000000, PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_z,
          accum_vector_operator_1_for_not_13_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0 <= 32'b00000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_read_data_and_18_enex5 ) begin
      input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0 <= input_mem_banks_read_read_data_lpi_1_dfm_1_5_31_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_6_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_22_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_30_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_38_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_46_itm_1
          <= 8'b00000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_3_cse ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_6_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[55:48]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_131_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_22_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[55:48]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_117_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_30_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[55:48]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_124_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_38_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[55:48]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_96_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_46_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[55:48]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_110_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1_7_4
          <= 4'b0000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1_3_0
          <= 4'b0000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_4_ssc ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1_7_4
          <= weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm[7:4];
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1_3_0
          <= MUX_v_4_2_2(rva_out_reg_data_39_36_sva_dfm_1_4, (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm[3:0]),
          crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_7_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_5_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_3_itm_1
          <= 8'b00000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_9_cse ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_7_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[63:56]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_132_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_5_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[47:40]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_133_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_3_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[31:24]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_135_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1_7
          <= 1'b0;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1_6_0
          <= 7'b0000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1_7_4
          <= 4'b0000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1_3_0
          <= 4'b0000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_10_ssc ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1_7
          <= weight_mem_banks_load_store_for_else_mux1h_11_nl & (~ or_dcpl_679);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1_6_0
          <= MUX_v_7_2_2(7'b0000000, weight_mem_banks_load_store_for_else_mux1h_38_nl,
          not_2441_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1_7_4
          <= MUX_v_4_2_2(4'b0000, weight_mem_banks_load_store_for_else_mux1h_18_nl,
          not_2442_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1_3_0
          <= MUX_v_4_2_2(4'b0000, weight_mem_banks_load_store_for_else_mux1h_39_nl,
          not_2443_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_23_itm_1
          <= 8'b00000000;
    end
    else if ( PECoreRun_wen & mux_110_nl & and_dcpl_228 & while_stage_0_6 ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_23_itm_1
          <= MUX_v_8_2_2(8'b00000000, mux1h_2_nl, not_2450_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_21_itm_1
          <= 8'b00000000;
    end
    else if ( PECoreRun_wen & (~ mux_117_nl) & while_stage_0_6 ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_21_itm_1
          <= MUX_v_8_2_2(8'b00000000, mux_489_nl, nor_522_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_29_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_28_itm_1
          <= 8'b00000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_17_cse ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_29_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[47:40]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_126_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_28_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[39:32]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_127_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_itm_1_7_6
          <= 2'b00;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_itm_1_5_0
          <= 6'b000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1_7
          <= 1'b0;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1_6_0
          <= 7'b0000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_itm_1_7
          <= 1'b0;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_itm_1_6_0
          <= 7'b0000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_20_ssc ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_itm_1_7_6
          <= MUX_v_2_2_2(2'b00, weight_mem_banks_load_store_for_else_mux1h_25_nl,
          not_2444_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_12_itm_1_5_0
          <= MUX_v_6_2_2(6'b000000, weight_mem_banks_load_store_for_else_mux1h_40_nl,
          not_2445_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1_7
          <= weight_mem_banks_load_store_for_else_mux1h_30_nl & (~ or_dcpl_679);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_11_itm_1_6_0
          <= MUX_v_7_2_2(7'b0000000, weight_mem_banks_load_store_for_else_mux1h_41_nl,
          not_2447_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_itm_1_7
          <= weight_mem_banks_load_store_for_else_mux1h_35_nl & (~ or_dcpl_679);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_10_itm_1_6_0
          <= MUX_v_7_2_2(7'b0000000, weight_mem_banks_load_store_for_else_mux1h_42_nl,
          not_2449_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_44_itm_1
          <= 8'b00000000;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_42_itm_1
          <= 8'b00000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_22_cse ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_44_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[39:32]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_113_nl);
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_42_itm_1
          <= MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[23:16]),
          weight_mem_write_arbxbar_xbar_for_1_for_not_72_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1_7
          <= 1'b0;
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1_6_0
          <= 7'b0000000;
      rva_out_reg_data_55_48_sva_dfm_1_5 <= 8'b00000000;
    end
    else if ( weight_mem_banks_load_store_for_else_and_27_ssc ) begin
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1_7
          <= weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm[7];
      weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1_6_0
          <= MUX_v_7_2_2(rva_out_reg_data_62_56_sva_dfm_1_4, (weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm[6:0]),
          crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
      rva_out_reg_data_55_48_sva_dfm_1_5 <= MUX_v_8_2_2(rva_out_reg_data_55_48_sva_dfm_1_4,
          weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_1_nl,
          crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_mem_write_arbxbar_xbar_for_empty_sva_2 <= 8'b00000000;
    end
    else if ( weight_mem_write_arbxbar_xbar_for_empty_and_enex5 ) begin
      weight_mem_write_arbxbar_xbar_for_empty_sva_2 <= weight_mem_write_arbxbar_xbar_for_empty_sva_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_reg_data_sva_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( rva_in_reg_data_and_tmp ) begin
      rva_in_reg_data_sva_1 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_6 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
        | PECore_RunMac_PECore_RunMac_if_and_svs_st_5)) & while_stage_0_7 ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_6 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_st_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_3 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~((weight_mem_write_arbxbar_xbar_for_lshift_tmp[1])
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2))
        & while_stage_0_4 ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_3 <= MUX_s_1_2_2(PECore_RunMac_PECore_RunMac_if_and_svs_st_2,
          (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[1]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ProductSum_for_asn_16_itm_3 <= 1'b0;
      ProductSum_for_asn_25_itm_3 <= 1'b0;
      ProductSum_for_asn_42_itm_3 <= 1'b0;
      ProductSum_for_asn_51_itm_3 <= 1'b0;
      ProductSum_for_asn_64_itm_3 <= 1'b0;
      ProductSum_for_asn_73_itm_3 <= 1'b0;
    end
    else if ( ProductSum_for_and_24_cse ) begin
      ProductSum_for_asn_16_itm_3 <= MUX_s_1_2_2(ProductSum_for_asn_16_itm_2, (weight_mem_write_arbxbar_xbar_for_lshift_tmp[2]),
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
      ProductSum_for_asn_25_itm_3 <= MUX_s_1_2_2(ProductSum_for_asn_25_itm_2, (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3]),
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
      ProductSum_for_asn_42_itm_3 <= MUX_s_1_2_2(ProductSum_for_asn_42_itm_2, (weight_mem_write_arbxbar_xbar_for_lshift_tmp[4]),
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
      ProductSum_for_asn_51_itm_3 <= MUX_s_1_2_2(ProductSum_for_asn_51_itm_2, (weight_mem_write_arbxbar_xbar_for_lshift_tmp[5]),
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
      ProductSum_for_asn_64_itm_3 <= MUX_s_1_2_2(ProductSum_for_asn_64_itm_2, (weight_mem_write_arbxbar_xbar_for_lshift_tmp[6]),
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
      ProductSum_for_asn_73_itm_3 <= MUX_s_1_2_2(ProductSum_for_asn_73_itm_2, (weight_mem_write_arbxbar_xbar_for_lshift_tmp[7]),
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ProductSum_for_asn_82_itm_3 <= 1'b0;
      ProductSum_for_asn_98_itm_3 <= 1'b0;
    end
    else if ( ProductSum_for_and_30_cse ) begin
      ProductSum_for_asn_82_itm_3 <= ProductSum_for_asn_82_itm_2;
      ProductSum_for_asn_98_itm_3 <= ProductSum_for_asn_98_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_17_itm_1 <= 1'b0;
    end
    else if ( PECoreRun_wen & mux_122_nl & while_stage_0_5 ) begin
      crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_17_itm_1 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_9_itm_1,
          input_read_req_valid_lpi_1_dfm_1_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_7
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_7
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_5
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_5
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_8_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_7
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_6;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_7
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_6;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_5
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_4;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_5
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_1_read_data_and_4_enex5 ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_2 <= input_mem_banks_read_1_read_data_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_read_req_valid_lpi_1_dfm_1_7 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5 <= 1'b0;
      rva_out_reg_data_39_36_sva_dfm_4_2_3 <= 1'b0;
      rva_out_reg_data_39_36_sva_dfm_4_2_2 <= 1'b0;
      rva_out_reg_data_39_36_sva_dfm_4_2_1_0 <= 2'b00;
      rva_out_reg_data_46_40_sva_dfm_4_2_6_4 <= 3'b000;
    end
    else if ( input_read_req_valid_and_2_cse ) begin
      input_read_req_valid_lpi_1_dfm_1_7 <= input_read_req_valid_lpi_1_dfm_1_6;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_5 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_4;
      rva_out_reg_data_39_36_sva_dfm_4_2_3 <= rva_out_reg_data_39_36_sva_dfm_4_1_3;
      rva_out_reg_data_39_36_sva_dfm_4_2_2 <= rva_out_reg_data_39_36_sva_dfm_4_1_2;
      rva_out_reg_data_39_36_sva_dfm_4_2_1_0 <= rva_out_reg_data_39_36_sva_dfm_4_1_1_0;
      rva_out_reg_data_46_40_sva_dfm_4_2_6_4 <= rva_out_reg_data_46_40_sva_dfm_4_1_6_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_7 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_7 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_6 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_7 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_11_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_7 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_6;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_7 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_6;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_6 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_1_5;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_7 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_5 <= 6'b000000;
    end
    else if ( rva_out_reg_data_and_91_enex5 ) begin
      rva_out_reg_data_30_25_sva_dfm_5 <= weight_mem_run_3_for_5_mux_12_itm_1_5_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_23_17_sva_dfm_5 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_92_enex5 ) begin
      rva_out_reg_data_23_17_sva_dfm_5 <= weight_mem_run_3_for_5_mux_11_itm_1_6_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_7 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_93_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_7 <= weight_mem_run_3_for_5_mux_10_itm_1_6_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_4_2 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_94_enex5 ) begin
      rva_out_reg_data_35_32_sva_dfm_4_2 <= rva_out_reg_data_35_32_sva_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_56_sva_dfm_4_2 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_95_enex5 ) begin
      rva_out_reg_data_62_56_sva_dfm_4_2 <= rva_out_reg_data_62_56_sva_dfm_4_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_7 <= 1'b0;
      accum_vector_operator_1_for_asn_70_itm_6 <= 1'b0;
      accum_vector_operator_1_for_asn_61_itm_6 <= 1'b0;
      accum_vector_operator_1_for_asn_52_itm_6 <= 1'b0;
      accum_vector_operator_1_for_asn_43_itm_6 <= 1'b0;
      accum_vector_operator_1_for_asn_34_itm_6 <= 1'b0;
      accum_vector_operator_1_for_asn_25_itm_6 <= 1'b0;
      accum_vector_operator_1_for_asn_16_itm_6 <= 1'b0;
      accum_vector_operator_1_for_asn_7_itm_6 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_7 <= 1'b0;
    end
    else if ( PECore_RunScale_if_and_3_cse ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_7 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_6;
      accum_vector_operator_1_for_asn_70_itm_6 <= accum_vector_operator_1_for_asn_70_itm_5;
      accum_vector_operator_1_for_asn_61_itm_6 <= accum_vector_operator_1_for_asn_61_itm_5;
      accum_vector_operator_1_for_asn_52_itm_6 <= accum_vector_operator_1_for_asn_52_itm_5;
      accum_vector_operator_1_for_asn_43_itm_6 <= accum_vector_operator_1_for_asn_43_itm_5;
      accum_vector_operator_1_for_asn_34_itm_6 <= accum_vector_operator_1_for_asn_34_itm_5;
      accum_vector_operator_1_for_asn_25_itm_6 <= accum_vector_operator_1_for_asn_25_itm_5;
      accum_vector_operator_1_for_asn_16_itm_6 <= accum_vector_operator_1_for_asn_16_itm_5;
      accum_vector_operator_1_for_asn_7_itm_6 <= accum_vector_operator_1_for_asn_7_itm_5;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_7 <= PECore_UpdateFSM_switch_lp_equal_tmp_2_6;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_7_sva_7 <= 23'b00000000000000000000000;
      accum_vector_data_7_sva_6 <= 23'b00000000000000000000000;
    end
    else if ( and_1320_cse ) begin
      accum_vector_data_7_sva_7 <= accum_vector_data_7_sva_7_mx1w0;
      accum_vector_data_7_sva_6 <= accum_vector_data_7_sva_6_mx1w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_6_sva_7 <= 23'b00000000000000000000000;
      accum_vector_data_6_sva_6 <= 23'b00000000000000000000000;
    end
    else if ( and_1332_cse ) begin
      accum_vector_data_6_sva_7 <= accum_vector_data_6_sva_7_mx1w0;
      accum_vector_data_6_sva_6 <= accum_vector_data_6_sva_6_mx1w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_5_sva_7 <= 23'b00000000000000000000000;
      accum_vector_data_5_sva_6 <= 23'b00000000000000000000000;
    end
    else if ( and_1344_cse ) begin
      accum_vector_data_5_sva_7 <= accum_vector_data_5_sva_7_mx1w0;
      accum_vector_data_5_sva_6 <= accum_vector_data_5_sva_6_mx1w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_4_sva_7 <= 23'b00000000000000000000000;
      accum_vector_data_4_sva_6 <= 23'b00000000000000000000000;
    end
    else if ( and_1356_cse ) begin
      accum_vector_data_4_sva_7 <= accum_vector_data_4_sva_7_mx1w0;
      accum_vector_data_4_sva_6 <= accum_vector_data_4_sva_6_mx1w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_3_sva_7 <= 23'b00000000000000000000000;
      accum_vector_data_3_sva_6 <= 23'b00000000000000000000000;
    end
    else if ( and_1368_cse ) begin
      accum_vector_data_3_sva_7 <= accum_vector_data_3_sva_7_mx1w0;
      accum_vector_data_3_sva_6 <= accum_vector_data_3_sva_6_mx1w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_1_sva_7 <= 23'b00000000000000000000000;
      accum_vector_data_1_sva_6 <= 23'b00000000000000000000000;
    end
    else if ( and_1380_cse ) begin
      accum_vector_data_1_sva_7 <= accum_vector_data_1_sva_7_mx1w0;
      accum_vector_data_1_sva_6 <= accum_vector_data_1_sva_6_mx1w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_0_sva_7 <= 23'b00000000000000000000000;
      accum_vector_data_0_sva_6 <= 23'b00000000000000000000000;
    end
    else if ( and_1392_cse ) begin
      accum_vector_data_0_sva_7 <= accum_vector_data_0_sva_7_mx1w0;
      accum_vector_data_0_sva_6 <= accum_vector_data_0_sva_6_mx1w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_5 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_1_1_itm_2_cse
        | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4))
        & while_stage_0_6 ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_5 <= reg_weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_3_1_itm_2_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_2 <= 1'b0;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_2 <= 1'b0;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_2 <= 1'b0;
      accum_vector_operator_1_for_asn_70_itm_1 <= 1'b0;
    end
    else if ( PECore_RunMac_if_and_5_cse ) begin
      PECore_RunMac_PECore_RunMac_if_and_svs_st_2 <= PECore_UpdateFSM_switch_lp_equal_tmp_3_1;
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_2 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_1_1;
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_2 <= PECore_UpdateFSM_switch_lp_equal_tmp_5_1;
      accum_vector_operator_1_for_asn_70_itm_1 <= accum_vector_data_7_sva_1_load_mx0w1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ProductSum_for_asn_16_itm_2 <= 1'b0;
      ProductSum_for_asn_25_itm_2 <= 1'b0;
      ProductSum_for_asn_42_itm_2 <= 1'b0;
      ProductSum_for_asn_51_itm_2 <= 1'b0;
      ProductSum_for_asn_64_itm_2 <= 1'b0;
      ProductSum_for_asn_73_itm_2 <= 1'b0;
      ProductSum_for_asn_82_itm_2 <= 1'b0;
      ProductSum_for_asn_98_itm_2 <= 1'b0;
    end
    else if ( ProductSum_for_and_32_cse ) begin
      ProductSum_for_asn_16_itm_2 <= PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_1;
      ProductSum_for_asn_25_itm_2 <= PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1;
      ProductSum_for_asn_42_itm_2 <= PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1;
      ProductSum_for_asn_51_itm_2 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_1;
      ProductSum_for_asn_64_itm_2 <= ProductSum_for_asn_64_itm_1;
      ProductSum_for_asn_73_itm_2 <= ProductSum_for_asn_73_itm_1;
      ProductSum_for_asn_82_itm_2 <= ProductSum_for_asn_82_itm_1;
      ProductSum_for_asn_98_itm_2 <= ProductSum_for_asn_98_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_6
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_6
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_4
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_4
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_12_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_6
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_5;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_6
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_5;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_4
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_3;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_4
          <= reg_pe_manager_base_weight_slc_pe_manager_base_weight_0_2_itm_2_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      input_mem_banks_read_1_read_data_lpi_1_dfm_1_1 <= MUX_v_64_2_2(input_mem_banks_read_1_for_mux_4_nl,
          input_mem_banks_read_read_data_sva_1, and_629_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_lpi_1_dfm_1_5_31_0 <= 32'b00000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_read_data_and_19_enex5 ) begin
      input_mem_banks_read_read_data_lpi_1_dfm_1_5_31_0 <= input_mem_banks_read_read_data_lpi_1_dfm_1_4[31:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_read_req_valid_lpi_1_dfm_1_6 <= 1'b0;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( input_read_req_valid_and_3_cse ) begin
      input_read_req_valid_lpi_1_dfm_1_6 <= crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_nor_11_itm_1;
      crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_4 <= crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_6 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_6 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_5 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_6 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_15_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_6 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_5;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_6 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_5;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_5 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_6 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_4_1 <= 4'b0000;
      rva_out_reg_data_62_56_sva_dfm_4_1 <= 7'b0000000;
      rva_out_reg_data_46_40_sva_dfm_4_1_3_0 <= 4'b0000;
      rva_out_reg_data_55_48_sva_dfm_4_1_7_4 <= 4'b0000;
      rva_out_reg_data_55_48_sva_dfm_4_1_3_0 <= 4'b0000;
    end
    else if ( and_1402_cse ) begin
      rva_out_reg_data_35_32_sva_dfm_4_1 <= MUX1HOT_v_4_4_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_13_itm_1_3_0,
          rva_out_reg_data_35_32_sva_dfm_6_mx1, (input_mem_banks_read_read_data_lpi_1_dfm_1_4[35:32]),
          (weight_port_read_out_data_0_4_sva_dfm_3_5_0[3:0]), {PECore_PushAxiRsp_if_asn_61
          , PECore_PushAxiRsp_if_asn_63 , PECore_PushAxiRsp_if_asn_65 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
      rva_out_reg_data_62_56_sva_dfm_4_1 <= MUX1HOT_v_7_4_2(weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_2_itm_1_6_0,
          rva_out_reg_data_62_56_sva_dfm_6_mx1, (input_mem_banks_read_read_data_lpi_1_dfm_1_4[62:56]),
          weight_port_read_out_data_0_7_sva_dfm_3_6_0, {PECore_PushAxiRsp_if_asn_61
          , PECore_PushAxiRsp_if_asn_63 , PECore_PushAxiRsp_if_asn_65 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
      rva_out_reg_data_46_40_sva_dfm_4_1_3_0 <= MUX1HOT_v_4_4_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1_6_0[3:0]),
          rva_out_reg_data_46_40_sva_dfm_6_mx1_3_0, (input_mem_banks_read_read_data_lpi_1_dfm_1_4[43:40]),
          weight_port_read_out_data_0_5_sva_dfm_3_3_0, {PECore_PushAxiRsp_if_asn_61
          , PECore_PushAxiRsp_if_asn_63 , PECore_PushAxiRsp_if_asn_65 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
      rva_out_reg_data_55_48_sva_dfm_4_1_7_4 <= MUX1HOT_v_4_4_2((rva_out_reg_data_55_48_sva_dfm_1_5[7:4]),
          rva_out_reg_data_55_48_sva_dfm_6_mx1_7_4, (input_mem_banks_read_read_data_lpi_1_dfm_1_4[55:52]),
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_8_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_64_63_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_2_0_8_7_0_sdt_47_40_sva_1_7_4,
          {PECore_PushAxiRsp_if_asn_61 , PECore_PushAxiRsp_if_asn_63 , PECore_PushAxiRsp_if_asn_65
          , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
      rva_out_reg_data_55_48_sva_dfm_4_1_3_0 <= MUX1HOT_v_4_4_2((rva_out_reg_data_55_48_sva_dfm_1_5[3:0]),
          rva_out_reg_data_55_48_sva_dfm_6_mx1_3_0, (input_mem_banks_read_read_data_lpi_1_dfm_1_4[51:48]),
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_8_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_64_63_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_2_0_8_7_0_sdt_47_40_sva_1_3_0,
          {PECore_PushAxiRsp_if_asn_61 , PECore_PushAxiRsp_if_asn_63 , PECore_PushAxiRsp_if_asn_65
          , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_6 <= 1'b0;
      accum_vector_operator_1_for_asn_70_itm_5 <= 1'b0;
      accum_vector_operator_1_for_asn_61_itm_5 <= 1'b0;
      accum_vector_operator_1_for_asn_52_itm_5 <= 1'b0;
      accum_vector_operator_1_for_asn_43_itm_5 <= 1'b0;
      accum_vector_operator_1_for_asn_34_itm_5 <= 1'b0;
      accum_vector_operator_1_for_asn_25_itm_5 <= 1'b0;
      accum_vector_operator_1_for_asn_16_itm_5 <= 1'b0;
      accum_vector_operator_1_for_asn_7_itm_5 <= 1'b0;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_6 <= 1'b0;
    end
    else if ( PECore_RunScale_if_and_5_cse ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_6 <= PECore_RunScale_PECore_RunScale_if_and_1_svs_5;
      accum_vector_operator_1_for_asn_70_itm_5 <= accum_vector_operator_1_for_asn_70_itm_4;
      accum_vector_operator_1_for_asn_61_itm_5 <= accum_vector_operator_1_for_asn_61_itm_4;
      accum_vector_operator_1_for_asn_52_itm_5 <= accum_vector_operator_1_for_asn_52_itm_4;
      accum_vector_operator_1_for_asn_43_itm_5 <= accum_vector_operator_1_for_asn_43_itm_4;
      accum_vector_operator_1_for_asn_34_itm_5 <= accum_vector_operator_1_for_asn_34_itm_4;
      accum_vector_operator_1_for_asn_25_itm_5 <= accum_vector_operator_1_for_asn_25_itm_4;
      accum_vector_operator_1_for_asn_16_itm_5 <= accum_vector_operator_1_for_asn_16_itm_4;
      accum_vector_operator_1_for_asn_7_itm_5 <= accum_vector_operator_1_for_asn_7_itm_4;
      PECore_UpdateFSM_switch_lp_equal_tmp_2_6 <= PECore_UpdateFSM_switch_lp_equal_tmp_2_5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_56_sva_dfm_6 <= 7'b0000000;
      rva_out_reg_data_35_32_sva_dfm_6 <= 4'b0000;
      rva_out_reg_data_55_48_sva_dfm_6_rsp_0 <= 4'b0000;
      rva_out_reg_data_55_48_sva_dfm_6_rsp_1 <= 4'b0000;
      rva_out_reg_data_46_40_sva_dfm_6_rsp_1 <= 4'b0000;
    end
    else if ( and_1411_cse ) begin
      rva_out_reg_data_62_56_sva_dfm_6 <= rva_out_reg_data_62_56_sva_dfm_6_mx1;
      rva_out_reg_data_35_32_sva_dfm_6 <= rva_out_reg_data_35_32_sva_dfm_6_mx1;
      rva_out_reg_data_55_48_sva_dfm_6_rsp_0 <= rva_out_reg_data_55_48_sva_dfm_6_mx1_7_4;
      rva_out_reg_data_55_48_sva_dfm_6_rsp_1 <= rva_out_reg_data_55_48_sva_dfm_6_mx1_3_0;
      rva_out_reg_data_46_40_sva_dfm_6_rsp_1 <= rva_out_reg_data_46_40_sva_dfm_6_mx1_3_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_PushAxiRsp_mux_13_itm_1 <= 1'b0;
    end
    else if ( PECoreRun_wen & ((and_dcpl_241 & rva_in_reg_rw_sva_5) | PECore_PushAxiRsp_mux_13_itm_1_mx0c1)
        ) begin
      PECore_PushAxiRsp_mux_13_itm_1 <= MUX_s_1_2_2(rva_out_reg_data_63_sva_dfm_7,
          weight_port_read_out_data_mux_20_nl, PECore_PushAxiRsp_mux_13_itm_1_mx0c1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_PushAxiRsp_mux_10_itm_1 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(nand_27_cse | rva_in_reg_rw_sva_5)) ) begin
      PECore_PushAxiRsp_mux_10_itm_1 <= MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_10_mx0w2,
          (weight_port_read_out_data_0_5_sva_dfm_3_7_4[3]), crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_lpi_1_dfm_1_4 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_read_data_and_20_tmp ) begin
      input_mem_banks_read_read_data_lpi_1_dfm_1_4 <= MUX1HOT_v_64_3_2(input_mem_banks_read_1_read_data_lpi_1_dfm_1_3,
          weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d, weight_mem_banks_read_1_read_data_1_lpi_1_dfm_1,
          {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
          , (~ or_tmp_382) , nor_469_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_0_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1419_tmp ) begin
      input_mem_banks_bank_a_0_sva_dfm_2 <= input_mem_banks_bank_a_0_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_1_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1422_tmp ) begin
      input_mem_banks_bank_a_1_sva_dfm_2 <= input_mem_banks_bank_a_1_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_2_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1425_tmp ) begin
      input_mem_banks_bank_a_2_sva_dfm_2 <= input_mem_banks_bank_a_2_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_3_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1428_tmp ) begin
      input_mem_banks_bank_a_3_sva_dfm_2 <= input_mem_banks_bank_a_3_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_4_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1431_tmp ) begin
      input_mem_banks_bank_a_4_sva_dfm_2 <= input_mem_banks_bank_a_4_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_5_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1434_tmp ) begin
      input_mem_banks_bank_a_5_sva_dfm_2 <= input_mem_banks_bank_a_5_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_6_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1437_tmp ) begin
      input_mem_banks_bank_a_6_sva_dfm_2 <= input_mem_banks_bank_a_6_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_7_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1440_tmp ) begin
      input_mem_banks_bank_a_7_sva_dfm_2 <= input_mem_banks_bank_a_7_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_8_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1443_tmp ) begin
      input_mem_banks_bank_a_8_sva_dfm_2 <= input_mem_banks_bank_a_8_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_9_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1446_tmp ) begin
      input_mem_banks_bank_a_9_sva_dfm_2 <= input_mem_banks_bank_a_9_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_10_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1449_tmp ) begin
      input_mem_banks_bank_a_10_sva_dfm_2 <= input_mem_banks_bank_a_10_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_11_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1452_tmp ) begin
      input_mem_banks_bank_a_11_sva_dfm_2 <= input_mem_banks_bank_a_11_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_12_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1455_tmp ) begin
      input_mem_banks_bank_a_12_sva_dfm_2 <= input_mem_banks_bank_a_12_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_13_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1458_tmp ) begin
      input_mem_banks_bank_a_13_sva_dfm_2 <= input_mem_banks_bank_a_13_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_14_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1461_tmp ) begin
      input_mem_banks_bank_a_14_sva_dfm_2 <= input_mem_banks_bank_a_14_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_15_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1464_tmp ) begin
      input_mem_banks_bank_a_15_sva_dfm_2 <= input_mem_banks_bank_a_15_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_16_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1467_tmp ) begin
      input_mem_banks_bank_a_16_sva_dfm_2 <= input_mem_banks_bank_a_16_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_17_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1470_tmp ) begin
      input_mem_banks_bank_a_17_sva_dfm_2 <= input_mem_banks_bank_a_17_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_18_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1473_tmp ) begin
      input_mem_banks_bank_a_18_sva_dfm_2 <= input_mem_banks_bank_a_18_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_19_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1476_tmp ) begin
      input_mem_banks_bank_a_19_sva_dfm_2 <= input_mem_banks_bank_a_19_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_20_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1479_tmp ) begin
      input_mem_banks_bank_a_20_sva_dfm_2 <= input_mem_banks_bank_a_20_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_21_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1482_tmp ) begin
      input_mem_banks_bank_a_21_sva_dfm_2 <= input_mem_banks_bank_a_21_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_22_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1485_tmp ) begin
      input_mem_banks_bank_a_22_sva_dfm_2 <= input_mem_banks_bank_a_22_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_23_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1488_tmp ) begin
      input_mem_banks_bank_a_23_sva_dfm_2 <= input_mem_banks_bank_a_23_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_24_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1491_tmp ) begin
      input_mem_banks_bank_a_24_sva_dfm_2 <= input_mem_banks_bank_a_24_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_25_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1494_tmp ) begin
      input_mem_banks_bank_a_25_sva_dfm_2 <= input_mem_banks_bank_a_25_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_26_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1497_tmp ) begin
      input_mem_banks_bank_a_26_sva_dfm_2 <= input_mem_banks_bank_a_26_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_27_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1500_tmp ) begin
      input_mem_banks_bank_a_27_sva_dfm_2 <= input_mem_banks_bank_a_27_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_28_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1503_tmp ) begin
      input_mem_banks_bank_a_28_sva_dfm_2 <= input_mem_banks_bank_a_28_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_29_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1506_tmp ) begin
      input_mem_banks_bank_a_29_sva_dfm_2 <= input_mem_banks_bank_a_29_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_30_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1509_tmp ) begin
      input_mem_banks_bank_a_30_sva_dfm_2 <= input_mem_banks_bank_a_30_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_31_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1512_tmp ) begin
      input_mem_banks_bank_a_31_sva_dfm_2 <= input_mem_banks_bank_a_31_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_32_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1515_tmp ) begin
      input_mem_banks_bank_a_32_sva_dfm_2 <= input_mem_banks_bank_a_32_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_33_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1518_tmp ) begin
      input_mem_banks_bank_a_33_sva_dfm_2 <= input_mem_banks_bank_a_33_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_34_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1521_tmp ) begin
      input_mem_banks_bank_a_34_sva_dfm_2 <= input_mem_banks_bank_a_34_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_35_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1524_tmp ) begin
      input_mem_banks_bank_a_35_sva_dfm_2 <= input_mem_banks_bank_a_35_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_36_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1527_tmp ) begin
      input_mem_banks_bank_a_36_sva_dfm_2 <= input_mem_banks_bank_a_36_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_37_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1530_tmp ) begin
      input_mem_banks_bank_a_37_sva_dfm_2 <= input_mem_banks_bank_a_37_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_38_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1533_tmp ) begin
      input_mem_banks_bank_a_38_sva_dfm_2 <= input_mem_banks_bank_a_38_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_39_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1536_tmp ) begin
      input_mem_banks_bank_a_39_sva_dfm_2 <= input_mem_banks_bank_a_39_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_40_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1539_tmp ) begin
      input_mem_banks_bank_a_40_sva_dfm_2 <= input_mem_banks_bank_a_40_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_41_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1542_tmp ) begin
      input_mem_banks_bank_a_41_sva_dfm_2 <= input_mem_banks_bank_a_41_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_42_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1545_tmp ) begin
      input_mem_banks_bank_a_42_sva_dfm_2 <= input_mem_banks_bank_a_42_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_43_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1548_tmp ) begin
      input_mem_banks_bank_a_43_sva_dfm_2 <= input_mem_banks_bank_a_43_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_44_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1551_tmp ) begin
      input_mem_banks_bank_a_44_sva_dfm_2 <= input_mem_banks_bank_a_44_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_45_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1554_tmp ) begin
      input_mem_banks_bank_a_45_sva_dfm_2 <= input_mem_banks_bank_a_45_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_46_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1557_tmp ) begin
      input_mem_banks_bank_a_46_sva_dfm_2 <= input_mem_banks_bank_a_46_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_47_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1560_tmp ) begin
      input_mem_banks_bank_a_47_sva_dfm_2 <= input_mem_banks_bank_a_47_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_48_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1563_tmp ) begin
      input_mem_banks_bank_a_48_sva_dfm_2 <= input_mem_banks_bank_a_48_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_49_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1566_tmp ) begin
      input_mem_banks_bank_a_49_sva_dfm_2 <= input_mem_banks_bank_a_49_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_50_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1569_tmp ) begin
      input_mem_banks_bank_a_50_sva_dfm_2 <= input_mem_banks_bank_a_50_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_51_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1572_tmp ) begin
      input_mem_banks_bank_a_51_sva_dfm_2 <= input_mem_banks_bank_a_51_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_52_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1575_tmp ) begin
      input_mem_banks_bank_a_52_sva_dfm_2 <= input_mem_banks_bank_a_52_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_53_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1578_tmp ) begin
      input_mem_banks_bank_a_53_sva_dfm_2 <= input_mem_banks_bank_a_53_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_54_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1581_tmp ) begin
      input_mem_banks_bank_a_54_sva_dfm_2 <= input_mem_banks_bank_a_54_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_55_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1584_tmp ) begin
      input_mem_banks_bank_a_55_sva_dfm_2 <= input_mem_banks_bank_a_55_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_56_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1587_tmp ) begin
      input_mem_banks_bank_a_56_sva_dfm_2 <= input_mem_banks_bank_a_56_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_57_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1590_tmp ) begin
      input_mem_banks_bank_a_57_sva_dfm_2 <= input_mem_banks_bank_a_57_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_58_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1593_tmp ) begin
      input_mem_banks_bank_a_58_sva_dfm_2 <= input_mem_banks_bank_a_58_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_59_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1596_tmp ) begin
      input_mem_banks_bank_a_59_sva_dfm_2 <= input_mem_banks_bank_a_59_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_60_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1599_tmp ) begin
      input_mem_banks_bank_a_60_sva_dfm_2 <= input_mem_banks_bank_a_60_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_61_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1602_tmp ) begin
      input_mem_banks_bank_a_61_sva_dfm_2 <= input_mem_banks_bank_a_61_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_62_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1605_tmp ) begin
      input_mem_banks_bank_a_62_sva_dfm_2 <= input_mem_banks_bank_a_62_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_63_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1608_tmp ) begin
      input_mem_banks_bank_a_63_sva_dfm_2 <= input_mem_banks_bank_a_63_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_64_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1611_tmp ) begin
      input_mem_banks_bank_a_64_sva_dfm_2 <= input_mem_banks_bank_a_64_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_65_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1614_tmp ) begin
      input_mem_banks_bank_a_65_sva_dfm_2 <= input_mem_banks_bank_a_65_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_66_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1617_tmp ) begin
      input_mem_banks_bank_a_66_sva_dfm_2 <= input_mem_banks_bank_a_66_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_67_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1620_tmp ) begin
      input_mem_banks_bank_a_67_sva_dfm_2 <= input_mem_banks_bank_a_67_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_68_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1623_tmp ) begin
      input_mem_banks_bank_a_68_sva_dfm_2 <= input_mem_banks_bank_a_68_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_69_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1626_tmp ) begin
      input_mem_banks_bank_a_69_sva_dfm_2 <= input_mem_banks_bank_a_69_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_70_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1629_tmp ) begin
      input_mem_banks_bank_a_70_sva_dfm_2 <= input_mem_banks_bank_a_70_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_71_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1632_tmp ) begin
      input_mem_banks_bank_a_71_sva_dfm_2 <= input_mem_banks_bank_a_71_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_72_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1635_tmp ) begin
      input_mem_banks_bank_a_72_sva_dfm_2 <= input_mem_banks_bank_a_72_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_73_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1638_tmp ) begin
      input_mem_banks_bank_a_73_sva_dfm_2 <= input_mem_banks_bank_a_73_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_74_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1641_tmp ) begin
      input_mem_banks_bank_a_74_sva_dfm_2 <= input_mem_banks_bank_a_74_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_75_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1644_tmp ) begin
      input_mem_banks_bank_a_75_sva_dfm_2 <= input_mem_banks_bank_a_75_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_76_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1647_tmp ) begin
      input_mem_banks_bank_a_76_sva_dfm_2 <= input_mem_banks_bank_a_76_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_77_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1650_tmp ) begin
      input_mem_banks_bank_a_77_sva_dfm_2 <= input_mem_banks_bank_a_77_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_78_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1653_tmp ) begin
      input_mem_banks_bank_a_78_sva_dfm_2 <= input_mem_banks_bank_a_78_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_79_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1656_tmp ) begin
      input_mem_banks_bank_a_79_sva_dfm_2 <= input_mem_banks_bank_a_79_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_80_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1659_tmp ) begin
      input_mem_banks_bank_a_80_sva_dfm_2 <= input_mem_banks_bank_a_80_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_81_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1662_tmp ) begin
      input_mem_banks_bank_a_81_sva_dfm_2 <= input_mem_banks_bank_a_81_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_82_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1665_tmp ) begin
      input_mem_banks_bank_a_82_sva_dfm_2 <= input_mem_banks_bank_a_82_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_83_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1668_tmp ) begin
      input_mem_banks_bank_a_83_sva_dfm_2 <= input_mem_banks_bank_a_83_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_84_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1671_tmp ) begin
      input_mem_banks_bank_a_84_sva_dfm_2 <= input_mem_banks_bank_a_84_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_85_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1674_tmp ) begin
      input_mem_banks_bank_a_85_sva_dfm_2 <= input_mem_banks_bank_a_85_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_86_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1677_tmp ) begin
      input_mem_banks_bank_a_86_sva_dfm_2 <= input_mem_banks_bank_a_86_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_87_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1680_tmp ) begin
      input_mem_banks_bank_a_87_sva_dfm_2 <= input_mem_banks_bank_a_87_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_88_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1683_tmp ) begin
      input_mem_banks_bank_a_88_sva_dfm_2 <= input_mem_banks_bank_a_88_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_89_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1686_tmp ) begin
      input_mem_banks_bank_a_89_sva_dfm_2 <= input_mem_banks_bank_a_89_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_90_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1689_tmp ) begin
      input_mem_banks_bank_a_90_sva_dfm_2 <= input_mem_banks_bank_a_90_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_91_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1692_tmp ) begin
      input_mem_banks_bank_a_91_sva_dfm_2 <= input_mem_banks_bank_a_91_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_92_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1695_tmp ) begin
      input_mem_banks_bank_a_92_sva_dfm_2 <= input_mem_banks_bank_a_92_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_93_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1698_tmp ) begin
      input_mem_banks_bank_a_93_sva_dfm_2 <= input_mem_banks_bank_a_93_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_94_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1701_tmp ) begin
      input_mem_banks_bank_a_94_sva_dfm_2 <= input_mem_banks_bank_a_94_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_95_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1704_tmp ) begin
      input_mem_banks_bank_a_95_sva_dfm_2 <= input_mem_banks_bank_a_95_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_96_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1707_tmp ) begin
      input_mem_banks_bank_a_96_sva_dfm_2 <= input_mem_banks_bank_a_96_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_97_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1710_tmp ) begin
      input_mem_banks_bank_a_97_sva_dfm_2 <= input_mem_banks_bank_a_97_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_98_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1713_tmp ) begin
      input_mem_banks_bank_a_98_sva_dfm_2 <= input_mem_banks_bank_a_98_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_99_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1716_tmp ) begin
      input_mem_banks_bank_a_99_sva_dfm_2 <= input_mem_banks_bank_a_99_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_100_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1719_tmp ) begin
      input_mem_banks_bank_a_100_sva_dfm_2 <= input_mem_banks_bank_a_100_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_101_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1722_tmp ) begin
      input_mem_banks_bank_a_101_sva_dfm_2 <= input_mem_banks_bank_a_101_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_102_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1725_tmp ) begin
      input_mem_banks_bank_a_102_sva_dfm_2 <= input_mem_banks_bank_a_102_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_103_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1728_tmp ) begin
      input_mem_banks_bank_a_103_sva_dfm_2 <= input_mem_banks_bank_a_103_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_104_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1731_tmp ) begin
      input_mem_banks_bank_a_104_sva_dfm_2 <= input_mem_banks_bank_a_104_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_105_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1734_tmp ) begin
      input_mem_banks_bank_a_105_sva_dfm_2 <= input_mem_banks_bank_a_105_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_106_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1737_tmp ) begin
      input_mem_banks_bank_a_106_sva_dfm_2 <= input_mem_banks_bank_a_106_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_107_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1740_tmp ) begin
      input_mem_banks_bank_a_107_sva_dfm_2 <= input_mem_banks_bank_a_107_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_108_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1743_tmp ) begin
      input_mem_banks_bank_a_108_sva_dfm_2 <= input_mem_banks_bank_a_108_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_109_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1746_tmp ) begin
      input_mem_banks_bank_a_109_sva_dfm_2 <= input_mem_banks_bank_a_109_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_110_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1749_tmp ) begin
      input_mem_banks_bank_a_110_sva_dfm_2 <= input_mem_banks_bank_a_110_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_111_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1752_tmp ) begin
      input_mem_banks_bank_a_111_sva_dfm_2 <= input_mem_banks_bank_a_111_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_112_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1755_tmp ) begin
      input_mem_banks_bank_a_112_sva_dfm_2 <= input_mem_banks_bank_a_112_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_113_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1758_tmp ) begin
      input_mem_banks_bank_a_113_sva_dfm_2 <= input_mem_banks_bank_a_113_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_114_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1761_tmp ) begin
      input_mem_banks_bank_a_114_sva_dfm_2 <= input_mem_banks_bank_a_114_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_115_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1764_tmp ) begin
      input_mem_banks_bank_a_115_sva_dfm_2 <= input_mem_banks_bank_a_115_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_116_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1767_tmp ) begin
      input_mem_banks_bank_a_116_sva_dfm_2 <= input_mem_banks_bank_a_116_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_117_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1770_tmp ) begin
      input_mem_banks_bank_a_117_sva_dfm_2 <= input_mem_banks_bank_a_117_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_118_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1773_tmp ) begin
      input_mem_banks_bank_a_118_sva_dfm_2 <= input_mem_banks_bank_a_118_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_119_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1776_tmp ) begin
      input_mem_banks_bank_a_119_sva_dfm_2 <= input_mem_banks_bank_a_119_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_120_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1779_tmp ) begin
      input_mem_banks_bank_a_120_sva_dfm_2 <= input_mem_banks_bank_a_120_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_121_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1782_tmp ) begin
      input_mem_banks_bank_a_121_sva_dfm_2 <= input_mem_banks_bank_a_121_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_122_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1785_tmp ) begin
      input_mem_banks_bank_a_122_sva_dfm_2 <= input_mem_banks_bank_a_122_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_123_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1788_tmp ) begin
      input_mem_banks_bank_a_123_sva_dfm_2 <= input_mem_banks_bank_a_123_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_124_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1791_tmp ) begin
      input_mem_banks_bank_a_124_sva_dfm_2 <= input_mem_banks_bank_a_124_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_125_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1794_tmp ) begin
      input_mem_banks_bank_a_125_sva_dfm_2 <= input_mem_banks_bank_a_125_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_126_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1797_tmp ) begin
      input_mem_banks_bank_a_126_sva_dfm_2 <= input_mem_banks_bank_a_126_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_127_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1800_tmp ) begin
      input_mem_banks_bank_a_127_sva_dfm_2 <= input_mem_banks_bank_a_127_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_128_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1803_tmp ) begin
      input_mem_banks_bank_a_128_sva_dfm_2 <= input_mem_banks_bank_a_128_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_129_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1806_tmp ) begin
      input_mem_banks_bank_a_129_sva_dfm_2 <= input_mem_banks_bank_a_129_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_130_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1809_tmp ) begin
      input_mem_banks_bank_a_130_sva_dfm_2 <= input_mem_banks_bank_a_130_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_131_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1812_tmp ) begin
      input_mem_banks_bank_a_131_sva_dfm_2 <= input_mem_banks_bank_a_131_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_132_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1815_tmp ) begin
      input_mem_banks_bank_a_132_sva_dfm_2 <= input_mem_banks_bank_a_132_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_133_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1818_tmp ) begin
      input_mem_banks_bank_a_133_sva_dfm_2 <= input_mem_banks_bank_a_133_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_134_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1821_tmp ) begin
      input_mem_banks_bank_a_134_sva_dfm_2 <= input_mem_banks_bank_a_134_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_135_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1824_tmp ) begin
      input_mem_banks_bank_a_135_sva_dfm_2 <= input_mem_banks_bank_a_135_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_136_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1827_tmp ) begin
      input_mem_banks_bank_a_136_sva_dfm_2 <= input_mem_banks_bank_a_136_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_137_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1830_tmp ) begin
      input_mem_banks_bank_a_137_sva_dfm_2 <= input_mem_banks_bank_a_137_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_138_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1833_tmp ) begin
      input_mem_banks_bank_a_138_sva_dfm_2 <= input_mem_banks_bank_a_138_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_139_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1836_tmp ) begin
      input_mem_banks_bank_a_139_sva_dfm_2 <= input_mem_banks_bank_a_139_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_140_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1839_tmp ) begin
      input_mem_banks_bank_a_140_sva_dfm_2 <= input_mem_banks_bank_a_140_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_141_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1842_tmp ) begin
      input_mem_banks_bank_a_141_sva_dfm_2 <= input_mem_banks_bank_a_141_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_142_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1845_tmp ) begin
      input_mem_banks_bank_a_142_sva_dfm_2 <= input_mem_banks_bank_a_142_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_143_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1848_tmp ) begin
      input_mem_banks_bank_a_143_sva_dfm_2 <= input_mem_banks_bank_a_143_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_144_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1851_tmp ) begin
      input_mem_banks_bank_a_144_sva_dfm_2 <= input_mem_banks_bank_a_144_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_145_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1854_tmp ) begin
      input_mem_banks_bank_a_145_sva_dfm_2 <= input_mem_banks_bank_a_145_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_146_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1857_tmp ) begin
      input_mem_banks_bank_a_146_sva_dfm_2 <= input_mem_banks_bank_a_146_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_147_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1860_tmp ) begin
      input_mem_banks_bank_a_147_sva_dfm_2 <= input_mem_banks_bank_a_147_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_148_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1863_tmp ) begin
      input_mem_banks_bank_a_148_sva_dfm_2 <= input_mem_banks_bank_a_148_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_149_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1866_tmp ) begin
      input_mem_banks_bank_a_149_sva_dfm_2 <= input_mem_banks_bank_a_149_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_150_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1869_tmp ) begin
      input_mem_banks_bank_a_150_sva_dfm_2 <= input_mem_banks_bank_a_150_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_151_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1872_tmp ) begin
      input_mem_banks_bank_a_151_sva_dfm_2 <= input_mem_banks_bank_a_151_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_152_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1875_tmp ) begin
      input_mem_banks_bank_a_152_sva_dfm_2 <= input_mem_banks_bank_a_152_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_153_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1878_tmp ) begin
      input_mem_banks_bank_a_153_sva_dfm_2 <= input_mem_banks_bank_a_153_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_154_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1881_tmp ) begin
      input_mem_banks_bank_a_154_sva_dfm_2 <= input_mem_banks_bank_a_154_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_155_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1884_tmp ) begin
      input_mem_banks_bank_a_155_sva_dfm_2 <= input_mem_banks_bank_a_155_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_156_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1887_tmp ) begin
      input_mem_banks_bank_a_156_sva_dfm_2 <= input_mem_banks_bank_a_156_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_157_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1890_tmp ) begin
      input_mem_banks_bank_a_157_sva_dfm_2 <= input_mem_banks_bank_a_157_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_158_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1893_tmp ) begin
      input_mem_banks_bank_a_158_sva_dfm_2 <= input_mem_banks_bank_a_158_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_159_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1896_tmp ) begin
      input_mem_banks_bank_a_159_sva_dfm_2 <= input_mem_banks_bank_a_159_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_160_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1899_tmp ) begin
      input_mem_banks_bank_a_160_sva_dfm_2 <= input_mem_banks_bank_a_160_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_161_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1902_tmp ) begin
      input_mem_banks_bank_a_161_sva_dfm_2 <= input_mem_banks_bank_a_161_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_162_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1905_tmp ) begin
      input_mem_banks_bank_a_162_sva_dfm_2 <= input_mem_banks_bank_a_162_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_163_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1908_tmp ) begin
      input_mem_banks_bank_a_163_sva_dfm_2 <= input_mem_banks_bank_a_163_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_164_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1911_tmp ) begin
      input_mem_banks_bank_a_164_sva_dfm_2 <= input_mem_banks_bank_a_164_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_165_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1914_tmp ) begin
      input_mem_banks_bank_a_165_sva_dfm_2 <= input_mem_banks_bank_a_165_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_166_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1917_tmp ) begin
      input_mem_banks_bank_a_166_sva_dfm_2 <= input_mem_banks_bank_a_166_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_167_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1920_tmp ) begin
      input_mem_banks_bank_a_167_sva_dfm_2 <= input_mem_banks_bank_a_167_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_168_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1923_tmp ) begin
      input_mem_banks_bank_a_168_sva_dfm_2 <= input_mem_banks_bank_a_168_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_169_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1926_tmp ) begin
      input_mem_banks_bank_a_169_sva_dfm_2 <= input_mem_banks_bank_a_169_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_170_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1929_tmp ) begin
      input_mem_banks_bank_a_170_sva_dfm_2 <= input_mem_banks_bank_a_170_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_171_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1932_tmp ) begin
      input_mem_banks_bank_a_171_sva_dfm_2 <= input_mem_banks_bank_a_171_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_172_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1935_tmp ) begin
      input_mem_banks_bank_a_172_sva_dfm_2 <= input_mem_banks_bank_a_172_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_173_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1938_tmp ) begin
      input_mem_banks_bank_a_173_sva_dfm_2 <= input_mem_banks_bank_a_173_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_174_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1941_tmp ) begin
      input_mem_banks_bank_a_174_sva_dfm_2 <= input_mem_banks_bank_a_174_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_175_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1944_tmp ) begin
      input_mem_banks_bank_a_175_sva_dfm_2 <= input_mem_banks_bank_a_175_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_176_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1947_tmp ) begin
      input_mem_banks_bank_a_176_sva_dfm_2 <= input_mem_banks_bank_a_176_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_177_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1950_tmp ) begin
      input_mem_banks_bank_a_177_sva_dfm_2 <= input_mem_banks_bank_a_177_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_178_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1953_tmp ) begin
      input_mem_banks_bank_a_178_sva_dfm_2 <= input_mem_banks_bank_a_178_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_179_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1956_tmp ) begin
      input_mem_banks_bank_a_179_sva_dfm_2 <= input_mem_banks_bank_a_179_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_180_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1959_tmp ) begin
      input_mem_banks_bank_a_180_sva_dfm_2 <= input_mem_banks_bank_a_180_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_181_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1962_tmp ) begin
      input_mem_banks_bank_a_181_sva_dfm_2 <= input_mem_banks_bank_a_181_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_182_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1965_tmp ) begin
      input_mem_banks_bank_a_182_sva_dfm_2 <= input_mem_banks_bank_a_182_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_183_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1968_tmp ) begin
      input_mem_banks_bank_a_183_sva_dfm_2 <= input_mem_banks_bank_a_183_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_184_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1971_tmp ) begin
      input_mem_banks_bank_a_184_sva_dfm_2 <= input_mem_banks_bank_a_184_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_185_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1974_tmp ) begin
      input_mem_banks_bank_a_185_sva_dfm_2 <= input_mem_banks_bank_a_185_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_186_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1977_tmp ) begin
      input_mem_banks_bank_a_186_sva_dfm_2 <= input_mem_banks_bank_a_186_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_187_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1980_tmp ) begin
      input_mem_banks_bank_a_187_sva_dfm_2 <= input_mem_banks_bank_a_187_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_188_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1983_tmp ) begin
      input_mem_banks_bank_a_188_sva_dfm_2 <= input_mem_banks_bank_a_188_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_189_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1986_tmp ) begin
      input_mem_banks_bank_a_189_sva_dfm_2 <= input_mem_banks_bank_a_189_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_190_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1989_tmp ) begin
      input_mem_banks_bank_a_190_sva_dfm_2 <= input_mem_banks_bank_a_190_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_191_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1992_tmp ) begin
      input_mem_banks_bank_a_191_sva_dfm_2 <= input_mem_banks_bank_a_191_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_192_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1995_tmp ) begin
      input_mem_banks_bank_a_192_sva_dfm_2 <= input_mem_banks_bank_a_192_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_193_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_1998_tmp ) begin
      input_mem_banks_bank_a_193_sva_dfm_2 <= input_mem_banks_bank_a_193_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_194_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2001_tmp ) begin
      input_mem_banks_bank_a_194_sva_dfm_2 <= input_mem_banks_bank_a_194_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_195_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2004_tmp ) begin
      input_mem_banks_bank_a_195_sva_dfm_2 <= input_mem_banks_bank_a_195_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_196_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2007_tmp ) begin
      input_mem_banks_bank_a_196_sva_dfm_2 <= input_mem_banks_bank_a_196_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_197_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2010_tmp ) begin
      input_mem_banks_bank_a_197_sva_dfm_2 <= input_mem_banks_bank_a_197_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_198_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2013_tmp ) begin
      input_mem_banks_bank_a_198_sva_dfm_2 <= input_mem_banks_bank_a_198_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_199_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2016_tmp ) begin
      input_mem_banks_bank_a_199_sva_dfm_2 <= input_mem_banks_bank_a_199_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_200_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2019_tmp ) begin
      input_mem_banks_bank_a_200_sva_dfm_2 <= input_mem_banks_bank_a_200_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_201_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2022_tmp ) begin
      input_mem_banks_bank_a_201_sva_dfm_2 <= input_mem_banks_bank_a_201_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_202_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2025_tmp ) begin
      input_mem_banks_bank_a_202_sva_dfm_2 <= input_mem_banks_bank_a_202_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_203_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2028_tmp ) begin
      input_mem_banks_bank_a_203_sva_dfm_2 <= input_mem_banks_bank_a_203_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_204_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2031_tmp ) begin
      input_mem_banks_bank_a_204_sva_dfm_2 <= input_mem_banks_bank_a_204_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_205_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2034_tmp ) begin
      input_mem_banks_bank_a_205_sva_dfm_2 <= input_mem_banks_bank_a_205_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_206_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2037_tmp ) begin
      input_mem_banks_bank_a_206_sva_dfm_2 <= input_mem_banks_bank_a_206_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_207_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2040_tmp ) begin
      input_mem_banks_bank_a_207_sva_dfm_2 <= input_mem_banks_bank_a_207_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_208_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2043_tmp ) begin
      input_mem_banks_bank_a_208_sva_dfm_2 <= input_mem_banks_bank_a_208_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_209_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2046_tmp ) begin
      input_mem_banks_bank_a_209_sva_dfm_2 <= input_mem_banks_bank_a_209_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_210_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2049_tmp ) begin
      input_mem_banks_bank_a_210_sva_dfm_2 <= input_mem_banks_bank_a_210_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_211_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2052_tmp ) begin
      input_mem_banks_bank_a_211_sva_dfm_2 <= input_mem_banks_bank_a_211_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_212_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2055_tmp ) begin
      input_mem_banks_bank_a_212_sva_dfm_2 <= input_mem_banks_bank_a_212_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_213_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2058_tmp ) begin
      input_mem_banks_bank_a_213_sva_dfm_2 <= input_mem_banks_bank_a_213_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_214_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2061_tmp ) begin
      input_mem_banks_bank_a_214_sva_dfm_2 <= input_mem_banks_bank_a_214_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_215_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2064_tmp ) begin
      input_mem_banks_bank_a_215_sva_dfm_2 <= input_mem_banks_bank_a_215_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_216_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2067_tmp ) begin
      input_mem_banks_bank_a_216_sva_dfm_2 <= input_mem_banks_bank_a_216_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_217_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2070_tmp ) begin
      input_mem_banks_bank_a_217_sva_dfm_2 <= input_mem_banks_bank_a_217_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_218_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2073_tmp ) begin
      input_mem_banks_bank_a_218_sva_dfm_2 <= input_mem_banks_bank_a_218_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_219_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2076_tmp ) begin
      input_mem_banks_bank_a_219_sva_dfm_2 <= input_mem_banks_bank_a_219_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_220_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2079_tmp ) begin
      input_mem_banks_bank_a_220_sva_dfm_2 <= input_mem_banks_bank_a_220_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_221_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2082_tmp ) begin
      input_mem_banks_bank_a_221_sva_dfm_2 <= input_mem_banks_bank_a_221_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_222_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2085_tmp ) begin
      input_mem_banks_bank_a_222_sva_dfm_2 <= input_mem_banks_bank_a_222_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_223_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2088_tmp ) begin
      input_mem_banks_bank_a_223_sva_dfm_2 <= input_mem_banks_bank_a_223_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_224_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2091_tmp ) begin
      input_mem_banks_bank_a_224_sva_dfm_2 <= input_mem_banks_bank_a_224_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_225_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2094_tmp ) begin
      input_mem_banks_bank_a_225_sva_dfm_2 <= input_mem_banks_bank_a_225_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_226_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2097_tmp ) begin
      input_mem_banks_bank_a_226_sva_dfm_2 <= input_mem_banks_bank_a_226_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_227_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2100_tmp ) begin
      input_mem_banks_bank_a_227_sva_dfm_2 <= input_mem_banks_bank_a_227_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_228_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2103_tmp ) begin
      input_mem_banks_bank_a_228_sva_dfm_2 <= input_mem_banks_bank_a_228_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_229_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2106_tmp ) begin
      input_mem_banks_bank_a_229_sva_dfm_2 <= input_mem_banks_bank_a_229_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_230_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2109_tmp ) begin
      input_mem_banks_bank_a_230_sva_dfm_2 <= input_mem_banks_bank_a_230_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_231_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2112_tmp ) begin
      input_mem_banks_bank_a_231_sva_dfm_2 <= input_mem_banks_bank_a_231_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_232_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2115_tmp ) begin
      input_mem_banks_bank_a_232_sva_dfm_2 <= input_mem_banks_bank_a_232_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_233_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2118_tmp ) begin
      input_mem_banks_bank_a_233_sva_dfm_2 <= input_mem_banks_bank_a_233_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_234_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2121_tmp ) begin
      input_mem_banks_bank_a_234_sva_dfm_2 <= input_mem_banks_bank_a_234_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_235_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2124_tmp ) begin
      input_mem_banks_bank_a_235_sva_dfm_2 <= input_mem_banks_bank_a_235_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_236_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2127_tmp ) begin
      input_mem_banks_bank_a_236_sva_dfm_2 <= input_mem_banks_bank_a_236_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_237_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2130_tmp ) begin
      input_mem_banks_bank_a_237_sva_dfm_2 <= input_mem_banks_bank_a_237_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_238_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2133_tmp ) begin
      input_mem_banks_bank_a_238_sva_dfm_2 <= input_mem_banks_bank_a_238_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_239_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2136_tmp ) begin
      input_mem_banks_bank_a_239_sva_dfm_2 <= input_mem_banks_bank_a_239_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_240_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2139_tmp ) begin
      input_mem_banks_bank_a_240_sva_dfm_2 <= input_mem_banks_bank_a_240_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_241_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2142_tmp ) begin
      input_mem_banks_bank_a_241_sva_dfm_2 <= input_mem_banks_bank_a_241_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_242_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2145_tmp ) begin
      input_mem_banks_bank_a_242_sva_dfm_2 <= input_mem_banks_bank_a_242_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_243_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2148_tmp ) begin
      input_mem_banks_bank_a_243_sva_dfm_2 <= input_mem_banks_bank_a_243_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_244_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2151_tmp ) begin
      input_mem_banks_bank_a_244_sva_dfm_2 <= input_mem_banks_bank_a_244_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_245_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2154_tmp ) begin
      input_mem_banks_bank_a_245_sva_dfm_2 <= input_mem_banks_bank_a_245_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_246_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2157_tmp ) begin
      input_mem_banks_bank_a_246_sva_dfm_2 <= input_mem_banks_bank_a_246_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_247_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2160_tmp ) begin
      input_mem_banks_bank_a_247_sva_dfm_2 <= input_mem_banks_bank_a_247_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_248_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2163_tmp ) begin
      input_mem_banks_bank_a_248_sva_dfm_2 <= input_mem_banks_bank_a_248_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_249_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2166_tmp ) begin
      input_mem_banks_bank_a_249_sva_dfm_2 <= input_mem_banks_bank_a_249_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_250_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2169_tmp ) begin
      input_mem_banks_bank_a_250_sva_dfm_2 <= input_mem_banks_bank_a_250_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_251_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2172_tmp ) begin
      input_mem_banks_bank_a_251_sva_dfm_2 <= input_mem_banks_bank_a_251_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_252_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2175_tmp ) begin
      input_mem_banks_bank_a_252_sva_dfm_2 <= input_mem_banks_bank_a_252_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_253_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2178_tmp ) begin
      input_mem_banks_bank_a_253_sva_dfm_2 <= input_mem_banks_bank_a_253_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_254_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2181_tmp ) begin
      input_mem_banks_bank_a_254_sva_dfm_2 <= input_mem_banks_bank_a_254_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_bank_a_255_sva_dfm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_2184_tmp ) begin
      input_mem_banks_bank_a_255_sva_dfm_2 <= input_mem_banks_bank_a_255_sva_dfm_2_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_5
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_5
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_3
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_16_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_5
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_4;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_5
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_4;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_3
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_5 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_5 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_5 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_19_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_5 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_84_itm_mx0w0,
          PECore_DecodeAxiRead_switch_lp_equal_tmp_3_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_5 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_72_itm_1_1,
          PECore_DecodeAxiRead_switch_lp_equal_tmp_2_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_4 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_71_itm_1_1,
          PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
      PECore_DecodeAxiRead_switch_lp_nor_tmp_5 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_94_itm_1,
          PECore_DecodeAxiRead_switch_lp_nor_tmp_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_base_input_sva <= 15'b000000000000000;
    end
    else if ( pe_manager_base_input_and_tmp ) begin
      pe_manager_base_input_sva <= MUX_v_15_2_2(pe_manager_base_input_sva_dfm_3_1,
          while_if_while_if_and_2_nl, and_692_cse);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_data_7_sva_1_load <= 1'b1;
      accum_vector_data_6_sva_1_load <= 1'b1;
      accum_vector_data_5_sva_1_load <= 1'b1;
      accum_vector_data_4_sva_1_load <= 1'b1;
      accum_vector_data_3_sva_1_load <= 1'b1;
      accum_vector_data_2_sva_1_load <= 1'b1;
      accum_vector_data_1_sva_1_load <= 1'b1;
      accum_vector_data_0_sva_1_load <= 1'b1;
    end
    else if ( and_680_cse ) begin
      accum_vector_data_7_sva_1_load <= accum_vector_data_7_sva_1_load_mx0w1 & (~
          and_dcpl_616);
      accum_vector_data_6_sva_1_load <= accum_vector_data_6_sva_1_load_mx0w1 & (~
          and_dcpl_616);
      accum_vector_data_5_sva_1_load <= accum_vector_data_5_sva_1_load_mx0w1 & (~
          and_dcpl_616);
      accum_vector_data_4_sva_1_load <= accum_vector_data_4_sva_1_load_mx0w1 & (~
          and_dcpl_616);
      accum_vector_data_3_sva_1_load <= accum_vector_data_3_sva_1_load_mx0w0 & (~
          and_dcpl_616);
      accum_vector_data_2_sva_1_load <= accum_vector_data_2_sva_1_load_mx0w0 & (~
          and_dcpl_616);
      accum_vector_data_1_sva_1_load <= accum_vector_data_1_sva_1_load_mx0w0 & (~
          and_dcpl_616);
      accum_vector_data_0_sva_1_load <= accum_vector_data_0_sva_1_load_mx0w0 & (~
          and_dcpl_616);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      pe_manager_base_input_sva_dfm_3_1 <= 15'b000000000000000;
    end
    else if ( (~((~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19:18]==2'b01) & rva_in_PopNB_mioi_return_rsc_z_mxwt
        & (~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])
        | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2]))) & (~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5:3]!=3'b000)))
        & nor_922_cse & nor_907_cse & nor_909_cse & nor_910_cse & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
        & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])) & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt))
        & while_stage_0_3)) & rva_in_reg_rw_and_6_cse ) begin
      pe_manager_base_input_sva_dfm_3_1 <= MUX_v_15_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[62:48]),
          pe_manager_base_input_sva_mx2, or_1096_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_3 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~ mux_177_nl) & while_stage_0_4 ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_st_3 <= MUX_s_1_2_2(PECore_RunScale_PECore_RunScale_if_and_1_svs_st_2,
          (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[3]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_4
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_4
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_2
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_19_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_4
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_3;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_4
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_3;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_2
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_4
          <= 1'b0;
    end
    else if ( PECoreRun_wen & mux_180_nl & while_stage_0_5 ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_4
          <= MUX_s_1_2_2((pe_manager_base_weight_sva[0]), PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_3,
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_2
          <= 1'b0;
    end
    else if ( PECoreRun_wen & mux_184_nl & while_stage_0_5 ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_2
          <= MUX_s_1_2_2((pe_manager_base_weight_sva[0]), PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_1,
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_4 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_4 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_4 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_23_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_4 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_7_itm_1,
          PECore_DecodeAxiRead_switch_lp_equal_tmp_3_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_4 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_6_itm_1,
          PECore_DecodeAxiRead_switch_lp_equal_tmp_2_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_nl,
          PECore_DecodeAxiRead_switch_lp_equal_tmp_1_2, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
      PECore_DecodeAxiRead_switch_lp_nor_tmp_4 <= MUX_s_1_2_2(crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_nl,
          PECore_DecodeAxiRead_switch_lp_nor_tmp_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_2 <= 6'b000000;
    end
    else if ( rva_out_reg_data_and_96_enex5 ) begin
      rva_out_reg_data_30_25_sva_dfm_2 <= rva_out_reg_data_30_25_sva_dfm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_23_17_sva_dfm_2 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_97_enex5 ) begin
      rva_out_reg_data_23_17_sva_dfm_2 <= rva_out_reg_data_23_17_sva_dfm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_4 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_98_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_4 <= rva_out_reg_data_15_9_sva_dfm_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_1_4 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_99_enex5 ) begin
      rva_out_reg_data_35_32_sva_dfm_1_4 <= rva_out_reg_data_35_32_sva_dfm_1_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_39_36_sva_dfm_1_4 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_100_enex5 ) begin
      rva_out_reg_data_39_36_sva_dfm_1_4 <= rva_out_reg_data_39_36_sva_dfm_1_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_46_40_sva_dfm_1_4 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_101_enex5 ) begin
      rva_out_reg_data_46_40_sva_dfm_1_4 <= rva_out_reg_data_46_40_sva_dfm_1_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_56_sva_dfm_1_4 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_102_enex5 ) begin
      rva_out_reg_data_62_56_sva_dfm_1_4 <= rva_out_reg_data_62_56_sva_dfm_1_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_1_4 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_103_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_1_4 <= rva_out_reg_data_55_48_sva_dfm_1_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_3 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~((weight_mem_write_arbxbar_xbar_for_lshift_tmp[0])
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2))
        & while_stage_0_4 ) begin
      PECore_PushOutput_PECore_PushOutput_if_and_svs_st_3 <= MUX_s_1_2_2(PECore_PushOutput_PECore_PushOutput_if_and_svs_st_2,
          (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[0]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_3
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_3
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_1
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_1
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_24_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_3
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_2;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_3
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_2;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_6_itm_1
          <= PECore_DecodeAxiRead_case_4_switch_lp_mux_2_nl & (~ PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_2);
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_4_itm_1
          <= PECore_DecodeAxiRead_case_4_switch_lp_mux_3_nl & (~ PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_3
          <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_3 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_2 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_25_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_3
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_2;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_3 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_2 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_read_req_valid_lpi_1_dfm_1_3 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~(reg_rva_in_reg_rw_sva_2_cse & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2))
        & while_stage_0_4 ) begin
      input_read_req_valid_lpi_1_dfm_1_3 <= accum_vector_operator_1_for_asn_7_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_3 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_3 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_27_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_3 <= PECore_DecodeAxiRead_switch_lp_equal_tmp_3_2;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_3 <= PECore_DecodeAxiRead_switch_lp_nor_tmp_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_30_25_sva_dfm_1 <= 6'b000000;
      rva_out_reg_data_23_17_sva_dfm_1 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_59_cse ) begin
      rva_out_reg_data_30_25_sva_dfm_1 <= MUX_v_6_2_2(6'b000000, (pe_manager_base_weight_sva_mx2[14:9]),
          PECore_DecodeAxiRead_case_4_switch_lp_nor_5_cse_1);
      rva_out_reg_data_23_17_sva_dfm_1 <= MUX_v_7_2_2(7'b0000000, (pe_manager_base_weight_sva_mx2[7:1]),
          PECore_DecodeAxiRead_case_4_switch_lp_nor_5_cse_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_3 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_104_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_3 <= rva_out_reg_data_15_9_sva_dfm_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_1_3 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_105_enex5 ) begin
      rva_out_reg_data_35_32_sva_dfm_1_3 <= rva_out_reg_data_35_32_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_39_36_sva_dfm_1_3 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_106_enex5 ) begin
      rva_out_reg_data_39_36_sva_dfm_1_3 <= rva_out_reg_data_39_36_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_46_40_sva_dfm_1_3 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_107_enex5 ) begin
      rva_out_reg_data_46_40_sva_dfm_1_3 <= rva_out_reg_data_46_40_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_56_sva_dfm_1_3 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_108_enex5 ) begin
      rva_out_reg_data_62_56_sva_dfm_1_3 <= rva_out_reg_data_62_56_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_1_3 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_109_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_1_3 <= rva_out_reg_data_55_48_sva_dfm_1_2;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_3 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~((weight_mem_write_arbxbar_xbar_for_lshift_tmp[2])
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2))
        & while_stage_0_4 ) begin
      PECore_RunScale_PECore_RunScale_if_and_1_svs_3 <= MUX_s_1_2_2(PECore_RunScale_PECore_RunScale_if_and_1_svs_st_2,
          (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[2]), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_2
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_2
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_29_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_2
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_1;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_2
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_2
          <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_30_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_2
          <= PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_2 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_1 <= 1'b0;
      PECore_DecodeAxiRead_switch_lp_nor_tmp_2 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_switch_lp_and_31_cse ) begin
      PECore_DecodeAxiRead_switch_lp_equal_tmp_3_2 <= MUX_s_1_2_2(accum_vector_data_4_sva_1_load_mx0w1,
          PECore_DecodeAxiRead_switch_lp_equal_tmp_3, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
      PECore_DecodeAxiRead_switch_lp_equal_tmp_1_1 <= MUX_s_1_2_2(PECore_UpdateFSM_switch_lp_equal_tmp_2_1,
          PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_1_nl,
          while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
      PECore_DecodeAxiRead_switch_lp_nor_tmp_2 <= MUX_s_1_2_2(accum_vector_data_5_sva_1_load_mx0w1,
          PECore_DecodeAxiRead_switch_lp_nor_tmp_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_15_9_sva_dfm_2 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_67_enex5 ) begin
      rva_out_reg_data_15_9_sva_dfm_2 <= rva_out_reg_data_15_9_sva_dfm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_35_32_sva_dfm_1_2 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_110_enex5 ) begin
      rva_out_reg_data_35_32_sva_dfm_1_2 <= rva_out_reg_data_35_32_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_39_36_sva_dfm_1_2 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_111_enex5 ) begin
      rva_out_reg_data_39_36_sva_dfm_1_2 <= rva_out_reg_data_39_36_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_46_40_sva_dfm_1_2 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_112_enex5 ) begin
      rva_out_reg_data_46_40_sva_dfm_1_2 <= rva_out_reg_data_46_40_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_62_56_sva_dfm_1_2 <= 7'b0000000;
    end
    else if ( rva_out_reg_data_and_113_enex5 ) begin
      rva_out_reg_data_62_56_sva_dfm_1_2 <= rva_out_reg_data_62_56_sva_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_1_2 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_114_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_1_2 <= pe_config_input_counter_sva_dfm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_2 <= 1'b0;
    end
    else if ( PECoreRun_wen & (~((~(and_dcpl_431 & (while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1[2])
        & (~(PECore_DecodeAxiRead_switch_lp_nor_tmp_1 | PECore_DecodeAxiRead_switch_lp_equal_tmp_3))
        & (~ PECore_DecodeAxiRead_switch_lp_equal_tmp_2) & PECore_DecodeAxiRead_switch_lp_nor_2_cse))
        & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1))
        & while_stage_0_3 ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_2 <= MUX_s_1_2_2(accum_vector_data_2_sva_1_load_mx0w0,
          PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_2 <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_2 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_33_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_2 <= MUX_s_1_2_2(accum_vector_data_3_sva_1_load_mx0w0,
          PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
      PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_2 <= MUX_s_1_2_2(accum_vector_data_1_sva_1_load_mx0w0,
          PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_2 <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_asn_1_itm_2 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_34_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_2 <= PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_1;
      PECore_DecodeAxiRead_case_4_switch_lp_asn_1_itm_2 <= PECore_DecodeAxiRead_case_4_switch_lp_asn_1_itm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_1
          <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_1
          <= 1'b0;
      rva_out_reg_data_15_9_sva_dfm_1 <= 7'b0000000;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_37_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_9_itm_1
          <= PECore_DecodeAxiRead_case_4_switch_lp_mux_7_nl & (~ PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_mx0w0);
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_8_itm_1
          <= PECore_DecodeAxiRead_case_4_switch_lp_mux_8_nl & (~ PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_mx0w0);
      rva_out_reg_data_15_9_sva_dfm_1 <= MUX_v_7_2_2(7'b0000000, (pe_manager_num_input_sva[7:1]),
          and_321_cse);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_1 <= 1'b0;
      PECore_DecodeAxiRead_case_4_switch_lp_asn_1_itm_1 <= 1'b0;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_39_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_1 <= pe_config_is_cluster_sva;
      PECore_DecodeAxiRead_case_4_switch_lp_asn_1_itm_1 <= pe_config_is_bias_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      input_mem_banks_read_read_data_sva_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( input_mem_banks_read_read_data_and_21_tmp ) begin
      input_mem_banks_read_read_data_sva_1 <= MUX_v_64_256_2(input_mem_banks_bank_a_0_sva_dfm_2_mx1,
          input_mem_banks_bank_a_1_sva_dfm_2_mx1, input_mem_banks_bank_a_2_sva_dfm_2_mx1,
          input_mem_banks_bank_a_3_sva_dfm_2_mx1, input_mem_banks_bank_a_4_sva_dfm_2_mx1,
          input_mem_banks_bank_a_5_sva_dfm_2_mx1, input_mem_banks_bank_a_6_sva_dfm_2_mx1,
          input_mem_banks_bank_a_7_sva_dfm_2_mx1, input_mem_banks_bank_a_8_sva_dfm_2_mx1,
          input_mem_banks_bank_a_9_sva_dfm_2_mx1, input_mem_banks_bank_a_10_sva_dfm_2_mx1,
          input_mem_banks_bank_a_11_sva_dfm_2_mx1, input_mem_banks_bank_a_12_sva_dfm_2_mx1,
          input_mem_banks_bank_a_13_sva_dfm_2_mx1, input_mem_banks_bank_a_14_sva_dfm_2_mx1,
          input_mem_banks_bank_a_15_sva_dfm_2_mx1, input_mem_banks_bank_a_16_sva_dfm_2_mx1,
          input_mem_banks_bank_a_17_sva_dfm_2_mx1, input_mem_banks_bank_a_18_sva_dfm_2_mx1,
          input_mem_banks_bank_a_19_sva_dfm_2_mx1, input_mem_banks_bank_a_20_sva_dfm_2_mx1,
          input_mem_banks_bank_a_21_sva_dfm_2_mx1, input_mem_banks_bank_a_22_sva_dfm_2_mx1,
          input_mem_banks_bank_a_23_sva_dfm_2_mx1, input_mem_banks_bank_a_24_sva_dfm_2_mx1,
          input_mem_banks_bank_a_25_sva_dfm_2_mx1, input_mem_banks_bank_a_26_sva_dfm_2_mx1,
          input_mem_banks_bank_a_27_sva_dfm_2_mx1, input_mem_banks_bank_a_28_sva_dfm_2_mx1,
          input_mem_banks_bank_a_29_sva_dfm_2_mx1, input_mem_banks_bank_a_30_sva_dfm_2_mx1,
          input_mem_banks_bank_a_31_sva_dfm_2_mx1, input_mem_banks_bank_a_32_sva_dfm_2_mx1,
          input_mem_banks_bank_a_33_sva_dfm_2_mx1, input_mem_banks_bank_a_34_sva_dfm_2_mx1,
          input_mem_banks_bank_a_35_sva_dfm_2_mx1, input_mem_banks_bank_a_36_sva_dfm_2_mx1,
          input_mem_banks_bank_a_37_sva_dfm_2_mx1, input_mem_banks_bank_a_38_sva_dfm_2_mx1,
          input_mem_banks_bank_a_39_sva_dfm_2_mx1, input_mem_banks_bank_a_40_sva_dfm_2_mx1,
          input_mem_banks_bank_a_41_sva_dfm_2_mx1, input_mem_banks_bank_a_42_sva_dfm_2_mx1,
          input_mem_banks_bank_a_43_sva_dfm_2_mx1, input_mem_banks_bank_a_44_sva_dfm_2_mx1,
          input_mem_banks_bank_a_45_sva_dfm_2_mx1, input_mem_banks_bank_a_46_sva_dfm_2_mx1,
          input_mem_banks_bank_a_47_sva_dfm_2_mx1, input_mem_banks_bank_a_48_sva_dfm_2_mx1,
          input_mem_banks_bank_a_49_sva_dfm_2_mx1, input_mem_banks_bank_a_50_sva_dfm_2_mx1,
          input_mem_banks_bank_a_51_sva_dfm_2_mx1, input_mem_banks_bank_a_52_sva_dfm_2_mx1,
          input_mem_banks_bank_a_53_sva_dfm_2_mx1, input_mem_banks_bank_a_54_sva_dfm_2_mx1,
          input_mem_banks_bank_a_55_sva_dfm_2_mx1, input_mem_banks_bank_a_56_sva_dfm_2_mx1,
          input_mem_banks_bank_a_57_sva_dfm_2_mx1, input_mem_banks_bank_a_58_sva_dfm_2_mx1,
          input_mem_banks_bank_a_59_sva_dfm_2_mx1, input_mem_banks_bank_a_60_sva_dfm_2_mx1,
          input_mem_banks_bank_a_61_sva_dfm_2_mx1, input_mem_banks_bank_a_62_sva_dfm_2_mx1,
          input_mem_banks_bank_a_63_sva_dfm_2_mx1, input_mem_banks_bank_a_64_sva_dfm_2_mx1,
          input_mem_banks_bank_a_65_sva_dfm_2_mx1, input_mem_banks_bank_a_66_sva_dfm_2_mx1,
          input_mem_banks_bank_a_67_sva_dfm_2_mx1, input_mem_banks_bank_a_68_sva_dfm_2_mx1,
          input_mem_banks_bank_a_69_sva_dfm_2_mx1, input_mem_banks_bank_a_70_sva_dfm_2_mx1,
          input_mem_banks_bank_a_71_sva_dfm_2_mx1, input_mem_banks_bank_a_72_sva_dfm_2_mx1,
          input_mem_banks_bank_a_73_sva_dfm_2_mx1, input_mem_banks_bank_a_74_sva_dfm_2_mx1,
          input_mem_banks_bank_a_75_sva_dfm_2_mx1, input_mem_banks_bank_a_76_sva_dfm_2_mx1,
          input_mem_banks_bank_a_77_sva_dfm_2_mx1, input_mem_banks_bank_a_78_sva_dfm_2_mx1,
          input_mem_banks_bank_a_79_sva_dfm_2_mx1, input_mem_banks_bank_a_80_sva_dfm_2_mx1,
          input_mem_banks_bank_a_81_sva_dfm_2_mx1, input_mem_banks_bank_a_82_sva_dfm_2_mx1,
          input_mem_banks_bank_a_83_sva_dfm_2_mx1, input_mem_banks_bank_a_84_sva_dfm_2_mx1,
          input_mem_banks_bank_a_85_sva_dfm_2_mx1, input_mem_banks_bank_a_86_sva_dfm_2_mx1,
          input_mem_banks_bank_a_87_sva_dfm_2_mx1, input_mem_banks_bank_a_88_sva_dfm_2_mx1,
          input_mem_banks_bank_a_89_sva_dfm_2_mx1, input_mem_banks_bank_a_90_sva_dfm_2_mx1,
          input_mem_banks_bank_a_91_sva_dfm_2_mx1, input_mem_banks_bank_a_92_sva_dfm_2_mx1,
          input_mem_banks_bank_a_93_sva_dfm_2_mx1, input_mem_banks_bank_a_94_sva_dfm_2_mx1,
          input_mem_banks_bank_a_95_sva_dfm_2_mx1, input_mem_banks_bank_a_96_sva_dfm_2_mx1,
          input_mem_banks_bank_a_97_sva_dfm_2_mx1, input_mem_banks_bank_a_98_sva_dfm_2_mx1,
          input_mem_banks_bank_a_99_sva_dfm_2_mx1, input_mem_banks_bank_a_100_sva_dfm_2_mx1,
          input_mem_banks_bank_a_101_sva_dfm_2_mx1, input_mem_banks_bank_a_102_sva_dfm_2_mx1,
          input_mem_banks_bank_a_103_sva_dfm_2_mx1, input_mem_banks_bank_a_104_sva_dfm_2_mx1,
          input_mem_banks_bank_a_105_sva_dfm_2_mx1, input_mem_banks_bank_a_106_sva_dfm_2_mx1,
          input_mem_banks_bank_a_107_sva_dfm_2_mx1, input_mem_banks_bank_a_108_sva_dfm_2_mx1,
          input_mem_banks_bank_a_109_sva_dfm_2_mx1, input_mem_banks_bank_a_110_sva_dfm_2_mx1,
          input_mem_banks_bank_a_111_sva_dfm_2_mx1, input_mem_banks_bank_a_112_sva_dfm_2_mx1,
          input_mem_banks_bank_a_113_sva_dfm_2_mx1, input_mem_banks_bank_a_114_sva_dfm_2_mx1,
          input_mem_banks_bank_a_115_sva_dfm_2_mx1, input_mem_banks_bank_a_116_sva_dfm_2_mx1,
          input_mem_banks_bank_a_117_sva_dfm_2_mx1, input_mem_banks_bank_a_118_sva_dfm_2_mx1,
          input_mem_banks_bank_a_119_sva_dfm_2_mx1, input_mem_banks_bank_a_120_sva_dfm_2_mx1,
          input_mem_banks_bank_a_121_sva_dfm_2_mx1, input_mem_banks_bank_a_122_sva_dfm_2_mx1,
          input_mem_banks_bank_a_123_sva_dfm_2_mx1, input_mem_banks_bank_a_124_sva_dfm_2_mx1,
          input_mem_banks_bank_a_125_sva_dfm_2_mx1, input_mem_banks_bank_a_126_sva_dfm_2_mx1,
          input_mem_banks_bank_a_127_sva_dfm_2_mx1, input_mem_banks_bank_a_128_sva_dfm_2_mx1,
          input_mem_banks_bank_a_129_sva_dfm_2_mx1, input_mem_banks_bank_a_130_sva_dfm_2_mx1,
          input_mem_banks_bank_a_131_sva_dfm_2_mx1, input_mem_banks_bank_a_132_sva_dfm_2_mx1,
          input_mem_banks_bank_a_133_sva_dfm_2_mx1, input_mem_banks_bank_a_134_sva_dfm_2_mx1,
          input_mem_banks_bank_a_135_sva_dfm_2_mx1, input_mem_banks_bank_a_136_sva_dfm_2_mx1,
          input_mem_banks_bank_a_137_sva_dfm_2_mx1, input_mem_banks_bank_a_138_sva_dfm_2_mx1,
          input_mem_banks_bank_a_139_sva_dfm_2_mx1, input_mem_banks_bank_a_140_sva_dfm_2_mx1,
          input_mem_banks_bank_a_141_sva_dfm_2_mx1, input_mem_banks_bank_a_142_sva_dfm_2_mx1,
          input_mem_banks_bank_a_143_sva_dfm_2_mx1, input_mem_banks_bank_a_144_sva_dfm_2_mx1,
          input_mem_banks_bank_a_145_sva_dfm_2_mx1, input_mem_banks_bank_a_146_sva_dfm_2_mx1,
          input_mem_banks_bank_a_147_sva_dfm_2_mx1, input_mem_banks_bank_a_148_sva_dfm_2_mx1,
          input_mem_banks_bank_a_149_sva_dfm_2_mx1, input_mem_banks_bank_a_150_sva_dfm_2_mx1,
          input_mem_banks_bank_a_151_sva_dfm_2_mx1, input_mem_banks_bank_a_152_sva_dfm_2_mx1,
          input_mem_banks_bank_a_153_sva_dfm_2_mx1, input_mem_banks_bank_a_154_sva_dfm_2_mx1,
          input_mem_banks_bank_a_155_sva_dfm_2_mx1, input_mem_banks_bank_a_156_sva_dfm_2_mx1,
          input_mem_banks_bank_a_157_sva_dfm_2_mx1, input_mem_banks_bank_a_158_sva_dfm_2_mx1,
          input_mem_banks_bank_a_159_sva_dfm_2_mx1, input_mem_banks_bank_a_160_sva_dfm_2_mx1,
          input_mem_banks_bank_a_161_sva_dfm_2_mx1, input_mem_banks_bank_a_162_sva_dfm_2_mx1,
          input_mem_banks_bank_a_163_sva_dfm_2_mx1, input_mem_banks_bank_a_164_sva_dfm_2_mx1,
          input_mem_banks_bank_a_165_sva_dfm_2_mx1, input_mem_banks_bank_a_166_sva_dfm_2_mx1,
          input_mem_banks_bank_a_167_sva_dfm_2_mx1, input_mem_banks_bank_a_168_sva_dfm_2_mx1,
          input_mem_banks_bank_a_169_sva_dfm_2_mx1, input_mem_banks_bank_a_170_sva_dfm_2_mx1,
          input_mem_banks_bank_a_171_sva_dfm_2_mx1, input_mem_banks_bank_a_172_sva_dfm_2_mx1,
          input_mem_banks_bank_a_173_sva_dfm_2_mx1, input_mem_banks_bank_a_174_sva_dfm_2_mx1,
          input_mem_banks_bank_a_175_sva_dfm_2_mx1, input_mem_banks_bank_a_176_sva_dfm_2_mx1,
          input_mem_banks_bank_a_177_sva_dfm_2_mx1, input_mem_banks_bank_a_178_sva_dfm_2_mx1,
          input_mem_banks_bank_a_179_sva_dfm_2_mx1, input_mem_banks_bank_a_180_sva_dfm_2_mx1,
          input_mem_banks_bank_a_181_sva_dfm_2_mx1, input_mem_banks_bank_a_182_sva_dfm_2_mx1,
          input_mem_banks_bank_a_183_sva_dfm_2_mx1, input_mem_banks_bank_a_184_sva_dfm_2_mx1,
          input_mem_banks_bank_a_185_sva_dfm_2_mx1, input_mem_banks_bank_a_186_sva_dfm_2_mx1,
          input_mem_banks_bank_a_187_sva_dfm_2_mx1, input_mem_banks_bank_a_188_sva_dfm_2_mx1,
          input_mem_banks_bank_a_189_sva_dfm_2_mx1, input_mem_banks_bank_a_190_sva_dfm_2_mx1,
          input_mem_banks_bank_a_191_sva_dfm_2_mx1, input_mem_banks_bank_a_192_sva_dfm_2_mx1,
          input_mem_banks_bank_a_193_sva_dfm_2_mx1, input_mem_banks_bank_a_194_sva_dfm_2_mx1,
          input_mem_banks_bank_a_195_sva_dfm_2_mx1, input_mem_banks_bank_a_196_sva_dfm_2_mx1,
          input_mem_banks_bank_a_197_sva_dfm_2_mx1, input_mem_banks_bank_a_198_sva_dfm_2_mx1,
          input_mem_banks_bank_a_199_sva_dfm_2_mx1, input_mem_banks_bank_a_200_sva_dfm_2_mx1,
          input_mem_banks_bank_a_201_sva_dfm_2_mx1, input_mem_banks_bank_a_202_sva_dfm_2_mx1,
          input_mem_banks_bank_a_203_sva_dfm_2_mx1, input_mem_banks_bank_a_204_sva_dfm_2_mx1,
          input_mem_banks_bank_a_205_sva_dfm_2_mx1, input_mem_banks_bank_a_206_sva_dfm_2_mx1,
          input_mem_banks_bank_a_207_sva_dfm_2_mx1, input_mem_banks_bank_a_208_sva_dfm_2_mx1,
          input_mem_banks_bank_a_209_sva_dfm_2_mx1, input_mem_banks_bank_a_210_sva_dfm_2_mx1,
          input_mem_banks_bank_a_211_sva_dfm_2_mx1, input_mem_banks_bank_a_212_sva_dfm_2_mx1,
          input_mem_banks_bank_a_213_sva_dfm_2_mx1, input_mem_banks_bank_a_214_sva_dfm_2_mx1,
          input_mem_banks_bank_a_215_sva_dfm_2_mx1, input_mem_banks_bank_a_216_sva_dfm_2_mx1,
          input_mem_banks_bank_a_217_sva_dfm_2_mx1, input_mem_banks_bank_a_218_sva_dfm_2_mx1,
          input_mem_banks_bank_a_219_sva_dfm_2_mx1, input_mem_banks_bank_a_220_sva_dfm_2_mx1,
          input_mem_banks_bank_a_221_sva_dfm_2_mx1, input_mem_banks_bank_a_222_sva_dfm_2_mx1,
          input_mem_banks_bank_a_223_sva_dfm_2_mx1, input_mem_banks_bank_a_224_sva_dfm_2_mx1,
          input_mem_banks_bank_a_225_sva_dfm_2_mx1, input_mem_banks_bank_a_226_sva_dfm_2_mx1,
          input_mem_banks_bank_a_227_sva_dfm_2_mx1, input_mem_banks_bank_a_228_sva_dfm_2_mx1,
          input_mem_banks_bank_a_229_sva_dfm_2_mx1, input_mem_banks_bank_a_230_sva_dfm_2_mx1,
          input_mem_banks_bank_a_231_sva_dfm_2_mx1, input_mem_banks_bank_a_232_sva_dfm_2_mx1,
          input_mem_banks_bank_a_233_sva_dfm_2_mx1, input_mem_banks_bank_a_234_sva_dfm_2_mx1,
          input_mem_banks_bank_a_235_sva_dfm_2_mx1, input_mem_banks_bank_a_236_sva_dfm_2_mx1,
          input_mem_banks_bank_a_237_sva_dfm_2_mx1, input_mem_banks_bank_a_238_sva_dfm_2_mx1,
          input_mem_banks_bank_a_239_sva_dfm_2_mx1, input_mem_banks_bank_a_240_sva_dfm_2_mx1,
          input_mem_banks_bank_a_241_sva_dfm_2_mx1, input_mem_banks_bank_a_242_sva_dfm_2_mx1,
          input_mem_banks_bank_a_243_sva_dfm_2_mx1, input_mem_banks_bank_a_244_sva_dfm_2_mx1,
          input_mem_banks_bank_a_245_sva_dfm_2_mx1, input_mem_banks_bank_a_246_sva_dfm_2_mx1,
          input_mem_banks_bank_a_247_sva_dfm_2_mx1, input_mem_banks_bank_a_248_sva_dfm_2_mx1,
          input_mem_banks_bank_a_249_sva_dfm_2_mx1, input_mem_banks_bank_a_250_sva_dfm_2_mx1,
          input_mem_banks_bank_a_251_sva_dfm_2_mx1, input_mem_banks_bank_a_252_sva_dfm_2_mx1,
          input_mem_banks_bank_a_253_sva_dfm_2_mx1, input_mem_banks_bank_a_254_sva_dfm_2_mx1,
          input_mem_banks_bank_a_255_sva_dfm_2_mx1, rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_vector_operator_1_for_asn_7_itm_1 <= 1'b0;
    end
    else if ( PECoreRun_wen & nand_372_cse & while_stage_0_3 ) begin
      accum_vector_operator_1_for_asn_7_itm_1 <= MUX_s_1_2_2(accum_vector_data_0_sva_1_load_mx0w0,
          ProductSum_for_asn_64_itm_1, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_1
          <= 1'b0;
      rva_out_reg_data_35_32_sva_dfm_1_1 <= 4'b0000;
      rva_out_reg_data_39_36_sva_dfm_1_1 <= 4'b0000;
      rva_out_reg_data_46_40_sva_dfm_1_1 <= 7'b0000000;
      rva_out_reg_data_62_56_sva_dfm_1_1 <= 7'b0000000;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_41_cse ) begin
      PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_PECore_DecodeAxiRead_case_4_switch_lp_and_itm_1
          <= (pe_config_num_output_sva[7]) & (~(and_321_cse | PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_mx0w0))
          & PECore_DecodeAxiRead_switch_lp_nor_13_cse_1;
      rva_out_reg_data_35_32_sva_dfm_1_1 <= PECore_DecodeAxiRead_case_4_switch_lp_mux_9_nl
          & (signext_4_1(~ PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_mx0w0))
          & ({{3{PECore_DecodeAxiRead_switch_lp_nor_13_cse_1}}, PECore_DecodeAxiRead_switch_lp_nor_13_cse_1});
      rva_out_reg_data_39_36_sva_dfm_1_1 <= (pe_manager_base_bias_sva[7:4]) & ({{3{and_321_cse}},
          and_321_cse}) & ({{3{PECore_DecodeAxiRead_switch_lp_nor_13_cse_1}}, PECore_DecodeAxiRead_switch_lp_nor_13_cse_1});
      rva_out_reg_data_46_40_sva_dfm_1_1 <= PECore_DecodeAxiRead_case_4_switch_lp_mux_10_nl
          & (signext_7_1(~ PECore_DecodeAxiRead_case_4_switch_lp_nor_tmp_mx0w0))
          & ({{6{PECore_DecodeAxiRead_switch_lp_nor_13_cse_1}}, PECore_DecodeAxiRead_switch_lp_nor_13_cse_1});
      rva_out_reg_data_62_56_sva_dfm_1_1 <= (pe_manager_base_input_sva_mx2[14:8])
          & ({{6{and_321_cse}}, and_321_cse}) & ({{6{PECore_DecodeAxiRead_switch_lp_nor_13_cse_1}},
          PECore_DecodeAxiRead_switch_lp_nor_13_cse_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_1_sva_dfm_2_7 <= 1'b0;
      weight_port_read_out_data_0_0_sva_dfm_2_7 <= 1'b0;
      weight_port_read_out_data_0_7_sva_dfm_2_7 <= 1'b0;
    end
    else if ( weight_port_read_out_data_and_14_cse ) begin
      weight_port_read_out_data_0_1_sva_dfm_2_7 <= MUX_s_1_2_2(weight_port_read_out_data_0_1_sva_dfm_mx0w0_7,
          PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_a_mx1_7, and_dcpl_32);
      weight_port_read_out_data_0_0_sva_dfm_2_7 <= MUX_s_1_2_2(weight_port_read_out_data_0_0_sva_dfm_mx0w0_7,
          weight_port_read_out_data_0_0_sva_dfm_3_7, and_dcpl_32);
      weight_port_read_out_data_0_7_sva_dfm_2_7 <= MUX_s_1_2_2(weight_port_read_out_data_0_7_sva_dfm_3_7,
          weight_port_read_out_data_0_7_sva_dfm_1_1_mx0_7, and_dcpl_32);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_1_sva_dfm_2_6_0 <= 7'b0000000;
    end
    else if ( mux_1256_nl & weight_mem_run_3_for_aelse_and_cse ) begin
      weight_port_read_out_data_0_1_sva_dfm_2_6_0 <= MUX_v_7_2_2(weight_port_read_out_data_0_1_sva_dfm_mx0w0_6_0,
          PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_a_mx1_6_0, and_dcpl_32);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_0_sva_dfm_2_6_0 <= 7'b0000000;
    end
    else if ( mux_1259_nl & weight_mem_run_3_for_aelse_and_cse ) begin
      weight_port_read_out_data_0_0_sva_dfm_2_6_0 <= MUX_v_7_2_2(weight_port_read_out_data_0_0_sva_dfm_mx0w0_6_0,
          weight_port_read_out_data_0_0_sva_dfm_3_6_0, and_dcpl_32);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_0_sva_dfm_3_rsp_0 <= 1'b0;
      weight_port_read_out_data_0_1_sva_dfm_3_rsp_0 <= 1'b0;
      weight_port_read_out_data_0_2_sva_dfm_3_rsp_0 <= 1'b0;
      weight_port_read_out_data_0_2_sva_dfm_3_rsp_1 <= 1'b0;
      weight_port_read_out_data_0_3_sva_dfm_3_rsp_0 <= 1'b0;
      weight_port_read_out_data_0_3_sva_dfm_3_rsp_1 <= 3'b000;
      weight_port_read_out_data_0_0_sva_dfm_3_rsp_1_6 <= 1'b0;
      weight_port_read_out_data_0_1_sva_dfm_3_rsp_1_6_4 <= 3'b000;
    end
    else if ( weight_port_read_out_data_and_92_cse ) begin
      weight_port_read_out_data_0_0_sva_dfm_3_rsp_0 <= weight_port_read_out_data_0_0_sva_dfm_2_7_1;
      weight_port_read_out_data_0_1_sva_dfm_3_rsp_0 <= weight_port_read_out_data_0_1_sva_dfm_2_7_1;
      weight_port_read_out_data_0_2_sva_dfm_3_rsp_0 <= weight_port_read_out_data_0_2_sva_dfm_2_7_1;
      weight_port_read_out_data_0_2_sva_dfm_3_rsp_1 <= weight_port_read_out_data_0_2_sva_dfm_2_6_1;
      weight_port_read_out_data_0_3_sva_dfm_3_rsp_0 <= weight_port_read_out_data_0_3_sva_dfm_2_7_1;
      weight_port_read_out_data_0_3_sva_dfm_3_rsp_1 <= weight_port_read_out_data_0_3_sva_dfm_2_6_4_1;
      weight_port_read_out_data_0_0_sva_dfm_3_rsp_1_6 <= reg_weight_port_read_out_data_0_0_sva_dfm_2_1_ftd;
      weight_port_read_out_data_0_1_sva_dfm_3_rsp_1_6_4 <= reg_weight_port_read_out_data_0_1_sva_dfm_2_1_ftd;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_2_sva_dfm_3_rsp_2 <= 6'b000000;
    end
    else if ( weight_port_read_out_data_and_106_enex5 ) begin
      weight_port_read_out_data_0_2_sva_dfm_3_rsp_2 <= weight_port_read_out_data_0_2_sva_dfm_2_5_0_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_6_sva_dfm_2_7_4 <= 4'b0000;
      weight_port_read_out_data_0_6_sva_dfm_2_3_0 <= 4'b0000;
    end
    else if ( weight_port_read_out_data_and_42_ssc ) begin
      weight_port_read_out_data_0_6_sva_dfm_2_7_4 <= MUX_v_4_2_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000000[7:4]),
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_8_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_64_63_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_2_0_8_7_0_sdt_47_40_sva_1_7_4,
          while_and_24_cse);
      weight_port_read_out_data_0_6_sva_dfm_2_3_0 <= MUX_v_4_2_2((crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000000[3:0]),
          crossbar_spec_PE_Weight_WordType_8U_8U_for_1_data_in_tmp_operator_for_8_slc_data_in_tmp_operator_for_slc_weight_mem_run_1_bank_read_out_data_64_63_0_data_in_tmp_operator_for_slc_data_in_tmp_operator_for_i_2_0_8_7_0_sdt_47_40_sva_1_3_0,
          while_and_24_cse);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_7_sva_dfm_2_6_0 <= 7'b0000000;
    end
    else if ( mux_1262_nl & weight_mem_run_3_for_aelse_and_cse ) begin
      weight_port_read_out_data_0_7_sva_dfm_2_6_0 <= MUX_v_7_2_2(weight_port_read_out_data_0_7_sva_dfm_3_6_0,
          weight_port_read_out_data_0_7_sva_dfm_1_1_mx0_6_0, and_dcpl_32);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_5_sva_dfm_2_7_4 <= 4'b0000;
      weight_port_read_out_data_0_5_sva_dfm_2_3_0 <= 4'b0000;
    end
    else if ( and_2218_cse ) begin
      weight_port_read_out_data_0_5_sva_dfm_2_7_4 <= MUX_v_4_2_2(weight_port_read_out_data_0_5_sva_dfm_3_7_4,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000001[7:4]),
          and_dcpl_32);
      weight_port_read_out_data_0_5_sva_dfm_2_3_0 <= MUX_v_4_2_2(weight_port_read_out_data_0_5_sva_dfm_3_3_0,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000001[3:0]),
          and_dcpl_32);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_4_sva_dfm_2_7 <= 1'b0;
      weight_port_read_out_data_0_4_sva_dfm_2_6 <= 1'b0;
      weight_port_read_out_data_0_3_sva_dfm_2_7 <= 1'b0;
      weight_port_read_out_data_0_3_sva_dfm_2_6_4 <= 3'b000;
      weight_port_read_out_data_0_2_sva_dfm_2_7 <= 1'b0;
      weight_port_read_out_data_0_2_sva_dfm_2_6 <= 1'b0;
    end
    else if ( weight_port_read_out_data_and_60_cse ) begin
      weight_port_read_out_data_0_4_sva_dfm_2_7 <= MUX_s_1_2_2(weight_port_read_out_data_0_4_sva_dfm_3_7,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000002[7]),
          and_dcpl_32);
      weight_port_read_out_data_0_4_sva_dfm_2_6 <= MUX_s_1_2_2(weight_port_read_out_data_0_4_sva_dfm_3_6,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000002[6]),
          and_dcpl_32);
      weight_port_read_out_data_0_3_sva_dfm_2_7 <= MUX_s_1_2_2(weight_port_read_out_data_0_3_sva_dfm_mx0w0_7,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000003[7]),
          and_dcpl_32);
      weight_port_read_out_data_0_3_sva_dfm_2_6_4 <= MUX_v_3_2_2(weight_port_read_out_data_0_3_sva_dfm_mx0w0_6_4,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000003[6:4]),
          and_dcpl_32);
      weight_port_read_out_data_0_2_sva_dfm_2_7 <= MUX_s_1_2_2(weight_port_read_out_data_0_2_sva_dfm_mx0w0_7,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000004[7]),
          and_dcpl_32);
      weight_port_read_out_data_0_2_sva_dfm_2_6 <= MUX_s_1_2_2(weight_port_read_out_data_0_2_sva_dfm_mx0w0_6,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000004[6]),
          and_dcpl_32);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_4_sva_dfm_2_5_0 <= 6'b000000;
    end
    else if ( mux_1283_nl & weight_mem_run_3_for_aelse_and_cse ) begin
      weight_port_read_out_data_0_4_sva_dfm_2_5_0 <= MUX_v_6_2_2(weight_port_read_out_data_0_4_sva_dfm_3_5_0,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000002[5:0]),
          and_dcpl_32);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_3_sva_dfm_2_3_0 <= 4'b0000;
    end
    else if ( mux_1290_nl & weight_mem_run_3_for_aelse_and_cse ) begin
      weight_port_read_out_data_0_3_sva_dfm_2_3_0 <= MUX_v_4_2_2(weight_port_read_out_data_0_3_sva_dfm_mx0w0_3_0,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000003[3:0]),
          and_dcpl_32);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_2_sva_dfm_2_5_0 <= 6'b000000;
    end
    else if ( mux_1297_nl & weight_mem_run_3_for_aelse_and_cse ) begin
      weight_port_read_out_data_0_2_sva_dfm_2_5_0 <= MUX_v_6_2_2(weight_port_read_out_data_0_2_sva_dfm_mx0w0_5_0,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000004[5:0]),
          and_dcpl_32);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_3_sva_dfm_3_rsp_2 <= 4'b0000;
    end
    else if ( weight_port_read_out_data_and_107_enex5 ) begin
      weight_port_read_out_data_0_3_sva_dfm_3_rsp_2 <= weight_port_read_out_data_0_3_sva_dfm_2_3_0_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_46_40_sva_dfm_4_3_rsp_1 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_115_enex5 ) begin
      rva_out_reg_data_46_40_sva_dfm_4_3_rsp_1 <= rva_out_reg_data_46_40_sva_dfm_4_2_3_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_4_3_rsp_0 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_116_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_4_3_rsp_0 <= rva_out_reg_data_55_48_sva_dfm_4_2_7_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_4_3_rsp_1 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_117_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_4_3_rsp_1 <= rva_out_reg_data_55_48_sva_dfm_4_2_3_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_0_sva_dfm_2_7_1 <= 1'b0;
      reg_weight_port_read_out_data_0_0_sva_dfm_2_1_ftd <= 1'b0;
      weight_port_read_out_data_0_1_sva_dfm_2_7_1 <= 1'b0;
      reg_weight_port_read_out_data_0_1_sva_dfm_2_1_ftd <= 3'b000;
      weight_port_read_out_data_0_2_sva_dfm_2_7_1 <= 1'b0;
      weight_port_read_out_data_0_2_sva_dfm_2_6_1 <= 1'b0;
      weight_port_read_out_data_0_3_sva_dfm_2_7_1 <= 1'b0;
      weight_port_read_out_data_0_3_sva_dfm_2_6_4_1 <= 3'b000;
    end
    else if ( weight_port_read_out_data_and_96_ssc ) begin
      weight_port_read_out_data_0_0_sva_dfm_2_7_1 <= weight_port_read_out_data_0_0_sva_dfm_1_7;
      reg_weight_port_read_out_data_0_0_sva_dfm_2_1_ftd <= weight_port_read_out_data_0_0_sva_dfm_1_6;
      weight_port_read_out_data_0_1_sva_dfm_2_7_1 <= weight_port_read_out_data_0_1_sva_dfm_1_7;
      reg_weight_port_read_out_data_0_1_sva_dfm_2_1_ftd <= weight_port_read_out_data_0_1_sva_dfm_1_6_4;
      weight_port_read_out_data_0_2_sva_dfm_2_7_1 <= weight_port_read_out_data_0_2_sva_dfm_1_7;
      weight_port_read_out_data_0_2_sva_dfm_2_6_1 <= weight_port_read_out_data_0_2_sva_dfm_1_6;
      weight_port_read_out_data_0_3_sva_dfm_2_7_1 <= weight_port_read_out_data_0_3_sva_dfm_1_7;
      weight_port_read_out_data_0_3_sva_dfm_2_6_4_1 <= weight_port_read_out_data_0_3_sva_dfm_1_6_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_2_1_ftd_1 <= 6'b000000;
    end
    else if ( weight_port_read_out_data_and_108_enex5 ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_2_1_ftd_1 <= weight_port_read_out_data_0_0_sva_dfm_1_5_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_2_1_ftd_1 <= 4'b0000;
    end
    else if ( weight_port_read_out_data_and_109_enex5 ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_2_1_ftd_1 <= weight_port_read_out_data_0_1_sva_dfm_1_3_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_2_sva_dfm_2_5_0_1 <= 6'b000000;
    end
    else if ( weight_port_read_out_data_and_110_enex5 ) begin
      weight_port_read_out_data_0_2_sva_dfm_2_5_0_1 <= weight_port_read_out_data_0_2_sva_dfm_1_5_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_3_sva_dfm_2_3_0_1 <= 4'b0000;
    end
    else if ( weight_port_read_out_data_and_111_enex5 ) begin
      weight_port_read_out_data_0_3_sva_dfm_2_3_0_1 <= weight_port_read_out_data_0_3_sva_dfm_1_3_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_46_40_sva_dfm_4_2_3_0 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_118_enex5 ) begin
      rva_out_reg_data_46_40_sva_dfm_4_2_3_0 <= rva_out_reg_data_46_40_sva_dfm_4_1_3_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_4_2_7_4 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_119_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_4_2_7_4 <= rva_out_reg_data_55_48_sva_dfm_4_1_7_4;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_55_48_sva_dfm_4_2_3_0 <= 4'b0000;
    end
    else if ( rva_out_reg_data_and_120_enex5 ) begin
      rva_out_reg_data_55_48_sva_dfm_4_2_3_0 <= rva_out_reg_data_55_48_sva_dfm_4_1_3_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_0_sva_dfm_1_7 <= 1'b0;
      weight_port_read_out_data_0_0_sva_dfm_1_6 <= 1'b0;
      weight_port_read_out_data_0_0_sva_dfm_1_5_0 <= 6'b000000;
      weight_port_read_out_data_0_1_sva_dfm_1_7 <= 1'b0;
      weight_port_read_out_data_0_1_sva_dfm_1_6_4 <= 3'b000;
      weight_port_read_out_data_0_1_sva_dfm_1_3_0 <= 4'b0000;
      weight_port_read_out_data_0_2_sva_dfm_1_7 <= 1'b0;
      weight_port_read_out_data_0_2_sva_dfm_1_6 <= 1'b0;
      weight_port_read_out_data_0_2_sva_dfm_1_5_0 <= 6'b000000;
      weight_port_read_out_data_0_3_sva_dfm_1_7 <= 1'b0;
      weight_port_read_out_data_0_3_sva_dfm_1_6_4 <= 3'b000;
      weight_port_read_out_data_0_3_sva_dfm_1_3_0 <= 4'b0000;
    end
    else if ( weight_port_read_out_data_and_100_ssc ) begin
      weight_port_read_out_data_0_0_sva_dfm_1_7 <= MUX1HOT_s_1_3_2(weight_port_read_out_data_0_0_sva_dfm_mx0w0_7,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000004[7]),
          weight_port_read_out_data_0_2_sva_dfm_2_7, {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , while_and_1123_rgt , while_while_nor_259_cse});
      weight_port_read_out_data_0_0_sva_dfm_1_6 <= MUX1HOT_s_1_3_2((weight_port_read_out_data_0_0_sva_dfm_mx0w0_6_0[6]),
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000004[6]),
          weight_port_read_out_data_0_2_sva_dfm_2_6, {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , while_and_1123_rgt , while_while_nor_259_cse});
      weight_port_read_out_data_0_0_sva_dfm_1_5_0 <= MUX1HOT_v_6_3_2((weight_port_read_out_data_0_0_sva_dfm_mx0w0_6_0[5:0]),
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000004[5:0]),
          weight_port_read_out_data_0_2_sva_dfm_2_5_0, {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , while_and_1123_rgt , while_while_nor_259_cse});
      weight_port_read_out_data_0_1_sva_dfm_1_7 <= MUX1HOT_s_1_3_2(weight_port_read_out_data_0_1_sva_dfm_mx0w0_7,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000003[7]),
          weight_port_read_out_data_0_3_sva_dfm_2_7, {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , while_and_1123_rgt , while_while_nor_259_cse});
      weight_port_read_out_data_0_1_sva_dfm_1_6_4 <= MUX1HOT_v_3_3_2((weight_port_read_out_data_0_1_sva_dfm_mx0w0_6_0[6:4]),
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000003[6:4]),
          weight_port_read_out_data_0_3_sva_dfm_2_6_4, {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , while_and_1123_rgt , while_while_nor_259_cse});
      weight_port_read_out_data_0_1_sva_dfm_1_3_0 <= MUX1HOT_v_4_3_2((weight_port_read_out_data_0_1_sva_dfm_mx0w0_6_0[3:0]),
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000003[3:0]),
          weight_port_read_out_data_0_3_sva_dfm_2_3_0, {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , while_and_1123_rgt , while_while_nor_259_cse});
      weight_port_read_out_data_0_2_sva_dfm_1_7 <= MUX1HOT_s_1_3_2(weight_port_read_out_data_0_2_sva_dfm_mx0w0_7,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000002[7]),
          weight_port_read_out_data_0_4_sva_dfm_2_7, {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , while_and_1123_rgt , while_while_nor_259_cse});
      weight_port_read_out_data_0_2_sva_dfm_1_6 <= MUX1HOT_s_1_3_2(weight_port_read_out_data_0_2_sva_dfm_mx0w0_6,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000002[6]),
          weight_port_read_out_data_0_4_sva_dfm_2_6, {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , while_and_1123_rgt , while_while_nor_259_cse});
      weight_port_read_out_data_0_2_sva_dfm_1_5_0 <= MUX1HOT_v_6_3_2(weight_port_read_out_data_0_2_sva_dfm_mx0w0_5_0,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000002[5:0]),
          weight_port_read_out_data_0_4_sva_dfm_2_5_0, {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , while_and_1123_rgt , while_while_nor_259_cse});
      weight_port_read_out_data_0_3_sva_dfm_1_7 <= MUX1HOT_s_1_3_2(weight_port_read_out_data_0_3_sva_dfm_mx0w0_7,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000001[7]),
          (weight_port_read_out_data_0_5_sva_dfm_2_7_4[3]), {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , while_and_1123_rgt , while_while_nor_259_cse});
      weight_port_read_out_data_0_3_sva_dfm_1_6_4 <= MUX1HOT_v_3_3_2(weight_port_read_out_data_0_3_sva_dfm_mx0w0_6_4,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000001[6:4]),
          (weight_port_read_out_data_0_5_sva_dfm_2_7_4[2:0]), {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , while_and_1123_rgt , while_while_nor_259_cse});
      weight_port_read_out_data_0_3_sva_dfm_1_3_0 <= MUX1HOT_v_4_3_2(weight_port_read_out_data_0_3_sva_dfm_mx0w0_3_0,
          (crossbar_spec_PE_Weight_WordType_8U_8U_1_for_1_data_in_tmp_operator_2_for_8_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_sdt_000001[3:0]),
          weight_port_read_out_data_0_5_sva_dfm_2_3_0, {while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5
          , while_and_1123_rgt , while_while_nor_259_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_39_36_sva_dfm_4_1_3 <= 1'b0;
      rva_out_reg_data_39_36_sva_dfm_4_1_2 <= 1'b0;
      rva_out_reg_data_39_36_sva_dfm_4_1_1_0 <= 2'b00;
      rva_out_reg_data_46_40_sva_dfm_4_1_6_4 <= 3'b000;
    end
    else if ( rva_out_reg_data_and_40_cse ) begin
      rva_out_reg_data_39_36_sva_dfm_4_1_3 <= MUX1HOT_s_1_4_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1_3_0[3]),
          rva_out_reg_data_39_36_sva_dfm_6_mx1_3, (input_mem_banks_read_read_data_lpi_1_dfm_1_4[39]),
          weight_port_read_out_data_0_4_sva_dfm_3_7, {PECore_PushAxiRsp_if_asn_61
          , PECore_PushAxiRsp_if_asn_63 , PECore_PushAxiRsp_if_asn_65 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
      rva_out_reg_data_39_36_sva_dfm_4_1_2 <= MUX1HOT_s_1_4_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1_3_0[2]),
          rva_out_reg_data_39_36_sva_dfm_6_mx1_2, (input_mem_banks_read_read_data_lpi_1_dfm_1_4[38]),
          weight_port_read_out_data_0_4_sva_dfm_3_6, {PECore_PushAxiRsp_if_asn_61
          , PECore_PushAxiRsp_if_asn_63 , PECore_PushAxiRsp_if_asn_65 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
      rva_out_reg_data_39_36_sva_dfm_4_1_1_0 <= MUX1HOT_v_2_4_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_14_itm_1_3_0[1:0]),
          rva_out_reg_data_39_36_sva_dfm_6_mx1_1_0, (input_mem_banks_read_read_data_lpi_1_dfm_1_4[37:36]),
          (weight_port_read_out_data_0_4_sva_dfm_3_5_0[5:4]), {PECore_PushAxiRsp_if_asn_61
          , PECore_PushAxiRsp_if_asn_63 , PECore_PushAxiRsp_if_asn_65 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
      rva_out_reg_data_46_40_sva_dfm_4_1_6_4 <= MUX1HOT_v_3_4_2((weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_15_itm_1_6_0[6:4]),
          rva_out_reg_data_46_40_sva_dfm_6_mx1_6_4, (input_mem_banks_read_read_data_lpi_1_dfm_1_4[46:44]),
          (weight_port_read_out_data_0_5_sva_dfm_3_7_4[2:0]), {PECore_PushAxiRsp_if_asn_61
          , PECore_PushAxiRsp_if_asn_63 , PECore_PushAxiRsp_if_asn_65 , crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_46_40_sva_dfm_6_rsp_0 <= 3'b000;
      rva_out_reg_data_39_36_sva_dfm_6_rsp_0 <= 1'b0;
      rva_out_reg_data_39_36_sva_dfm_6_rsp_1 <= 1'b0;
      rva_out_reg_data_39_36_sva_dfm_6_rsp_2 <= 2'b00;
    end
    else if ( rva_out_reg_data_and_45_cse ) begin
      rva_out_reg_data_46_40_sva_dfm_6_rsp_0 <= rva_out_reg_data_46_40_sva_dfm_6_mx1_6_4;
      rva_out_reg_data_39_36_sva_dfm_6_rsp_0 <= rva_out_reg_data_39_36_sva_dfm_6_mx1_3;
      rva_out_reg_data_39_36_sva_dfm_6_rsp_1 <= rva_out_reg_data_39_36_sva_dfm_6_mx1_2;
      rva_out_reg_data_39_36_sva_dfm_6_rsp_2 <= rva_out_reg_data_39_36_sva_dfm_6_mx1_1_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_1_ftd_1_rsp_1
          <= 5'b00000;
    end
    else if ( weight_port_read_out_data_and_112_enex5 ) begin
      reg_weight_port_read_out_data_slc_weight_port_read_out_data_0_0_7_1_itm_1_ftd_1_rsp_1
          <= weight_port_read_out_data_0_0_sva_dfm_3_rsp_1_5_0[5:1];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_0_sva_dfm_3_rsp_1_5_0 <= 6'b000000;
    end
    else if ( weight_port_read_out_data_and_113_enex5 ) begin
      weight_port_read_out_data_0_0_sva_dfm_3_rsp_1_5_0 <= reg_weight_port_read_out_data_0_0_sva_dfm_2_1_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_port_read_out_data_0_1_sva_dfm_3_rsp_1_3_0 <= 4'b0000;
    end
    else if ( weight_port_read_out_data_and_114_enex5 ) begin
      weight_port_read_out_data_0_1_sva_dfm_3_rsp_1_3_0 <= reg_weight_port_read_out_data_0_1_sva_dfm_2_1_ftd_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_8_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_88_enex5 | rva_out_reg_data_and_78_enex5 ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_8_enexo <= rva_out_reg_data_and_88_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_6_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_87_enex5 | rva_out_reg_data_and_79_enex5 ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_6_enexo <= rva_out_reg_data_and_87_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_6_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_86_enex5 | rva_out_reg_data_and_80_enex5 ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_6_enexo <= rva_out_reg_data_and_86_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_90_enex5 | rva_out_reg_data_and_81_enex5 ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_4_3_enexo <= rva_out_reg_data_and_90_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_116_enex5 | rva_out_reg_data_and_82_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_3_enexo <= rva_out_reg_data_and_116_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_3_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_117_enex5 | rva_out_reg_data_and_83_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_3_1_enexo <= rva_out_reg_data_and_117_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_3_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_115_enex5 | rva_out_reg_data_and_84_enex5 ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_3_1_enexo <= rva_out_reg_data_and_115_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_4_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_89_enex5 | rva_out_reg_data_and_85_enex5 ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_4_3_enexo <= rva_out_reg_data_and_89_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_1_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_26_enex5 | input_mem_banks_read_read_data_and_22_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_7_1_itm_1_enexo
          <= input_mem_banks_read_read_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_1_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_27_enex5 | input_mem_banks_read_read_data_and_23_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_15_9_itm_1_enexo
          <= input_mem_banks_read_read_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_1_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_28_enex5 | input_mem_banks_read_read_data_and_24_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_23_17_itm_1_enexo
          <= input_mem_banks_read_read_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_2_sva_dfm_3_2_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_106_enex5 | weight_port_read_out_data_and_104_enex5
        ) begin
      reg_weight_port_read_out_data_0_2_sva_dfm_3_2_enexo <= weight_port_read_out_data_and_106_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_3_2_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_107_enex5 | weight_port_read_out_data_and_105_enex5
        ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_3_2_enexo <= weight_port_read_out_data_and_107_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_1_enexo
          <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_29_enex5 | input_mem_banks_read_read_data_and_25_enex5
        ) begin
      reg_input_mem_banks_read_read_data_slc_input_mem_banks_read_read_data_30_25_itm_1_enexo
          <= input_mem_banks_read_read_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_4_enexo <= 1'b1;
    end
    else if ( input_mem_banks_read_1_read_data_and_7_enex5 | input_mem_banks_read_1_read_data_and_enex5
        ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_4_enexo <= input_mem_banks_read_1_read_data_and_7_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_4_enexo_1 <= 1'b1;
    end
    else if ( input_mem_banks_read_1_read_data_and_7_enex5 | input_mem_banks_read_1_read_data_and_6_enex5
        ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_4_enexo_1 <= input_mem_banks_read_1_read_data_and_7_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_000000
          <= 1'b1;
    end
    else if ( data_in_tmp_operator_2_for_and_tmp | weight_port_read_out_data_and_enex5
        ) begin
      reg_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_3_data_in_tmp_operator_2_for_7_slc_data_in_tmp_operator_2_for_slc_weight_mem_run_3_bank_read_out_data_64_63_0_data_in_tmp_operator_2_for_slc_data_in_tmp_operator_2_for_i_2_0_8_7_0_000000
          <= data_in_tmp_operator_2_for_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_3_enexo <= 1'b1;
    end
    else if ( input_mem_banks_read_1_read_data_and_3_enex5 | input_mem_banks_read_1_read_data_and_7_enex5
        ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_3_enexo <= input_mem_banks_read_1_read_data_and_3_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo <= 1'b1;
    end
    else if ( weight_read_addrs_and_9_cse | weight_read_addrs_and_7_enex5 ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo <= weight_read_addrs_and_9_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1_enexo <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 ) begin
      reg_Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1_enexo <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0_enexo
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_13_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0_enexo
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_13_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_3_enexo
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_26_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_3_enexo
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_26_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1_enexo
          <= 1'b1;
    end
    else if ( Arbiter_8U_Roundrobin_pick_1_and_22_cse | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5
        ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1_enexo
          <= Arbiter_8U_Roundrobin_pick_1_and_22_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0_enexo
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_22_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0_enexo
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_22_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_3_enexo
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_14_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_3_enexo
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_14_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_3_enexo
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_18_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_3_enexo
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_18_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_1 <= 1'b1;
    end
    else if ( weight_read_addrs_and_9_cse | weight_mem_read_arbxbar_xbar_1_for_3_and_enex5
        ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_1 <= weight_read_addrs_and_9_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1_enexo_1 <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 ) begin
      reg_Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1_enexo_1 <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_0_enexo
          <= 1'b1;
    end
    else if ( Arbiter_8U_Roundrobin_pick_1_and_15_cse | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5
        ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_7_1_0_enexo
          <= Arbiter_8U_Roundrobin_pick_1_and_15_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0_enexo_1
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_13_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_5_1_0_enexo_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_13_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_3_enexo_1
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_26_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_1_1_3_enexo_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_26_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1_enexo_1
          <= 1'b1;
    end
    else if ( Arbiter_8U_Roundrobin_pick_1_and_22_cse | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5
        ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_6_1_1_enexo_1
          <= Arbiter_8U_Roundrobin_pick_1_and_22_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0_enexo_1
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_22_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_2_1_0_enexo_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_22_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_3_enexo_1
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_14_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_4_1_3_enexo_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_14_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_3_enexo_1
          <= 1'b1;
    end
    else if ( nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_18_cse
        | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5 ) begin
      reg_nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_7_1_sva_3_1_3_enexo_1
          <= nvhls_set_slc_Arbiter_8U_Roundrobin_Mask_nvhls_nvhls_t_7U_nvuint_t_1_X_temp_and_18_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs_enexo
          <= 1'b1;
    end
    else if ( operator_15_false_1_and_cse | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5
        ) begin
      reg_weight_mem_read_arbxbar_xbar_1_for_3_8_operator_15_false_1_operator_15_false_1_or_svs_enexo
          <= operator_15_false_1_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_2 <= 1'b1;
    end
    else if ( weight_read_addrs_and_9_cse | weight_mem_read_arbxbar_xbar_1_for_3_and_20_enex5
        ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_3_enexo_2 <= weight_read_addrs_and_9_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_7_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_32_enex5 | weight_write_data_data_and_24_enex5
        ) begin
      reg_weight_write_data_data_0_7_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_32_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_6_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_33_enex5 | weight_write_data_data_and_25_enex5
        ) begin
      reg_weight_write_data_data_0_6_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_33_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_5_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_34_enex5 | weight_write_data_data_and_26_enex5
        ) begin
      reg_weight_write_data_data_0_5_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_34_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_4_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_35_enex5 | weight_write_data_data_and_27_enex5
        ) begin
      reg_weight_write_data_data_0_4_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_35_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_3_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_36_enex5 | weight_write_data_data_and_28_enex5
        ) begin
      reg_weight_write_data_data_0_3_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_36_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_2_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_37_enex5 | weight_write_data_data_and_29_enex5
        ) begin
      reg_weight_write_data_data_0_2_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_37_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_1_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_38_enex5 | weight_write_data_data_and_30_enex5
        ) begin
      reg_weight_write_data_data_0_1_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_38_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_0_lpi_1_dfm_1_2_6_enexo <= 1'b1;
    end
    else if ( weight_write_data_data_and_39_enex5 | weight_write_data_data_and_31_enex5
        ) begin
      reg_weight_write_data_data_0_0_lpi_1_dfm_1_2_6_enexo <= weight_write_data_data_and_39_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_addrs_lpi_1_dfm_1_2_enexo <= 1'b1;
    end
    else if ( weight_write_addrs_and_2_enex5 | weight_write_addrs_and_enex5 ) begin
      reg_weight_write_addrs_lpi_1_dfm_1_2_enexo <= weight_write_addrs_and_2_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_7_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_14_cse | weight_write_data_data_and_32_enex5 ) begin
      reg_weight_write_data_data_0_7_lpi_1_dfm_1_1_enexo <= while_if_and_14_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_6_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_14_cse | weight_write_data_data_and_33_enex5 ) begin
      reg_weight_write_data_data_0_6_lpi_1_dfm_1_1_enexo <= while_if_and_14_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_5_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_14_cse | weight_write_data_data_and_34_enex5 ) begin
      reg_weight_write_data_data_0_5_lpi_1_dfm_1_1_enexo <= while_if_and_14_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_4_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_14_cse | weight_write_data_data_and_35_enex5 ) begin
      reg_weight_write_data_data_0_4_lpi_1_dfm_1_1_enexo <= while_if_and_14_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_3_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_14_cse | weight_write_data_data_and_36_enex5 ) begin
      reg_weight_write_data_data_0_3_lpi_1_dfm_1_1_enexo <= while_if_and_14_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_2_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_14_cse | weight_write_data_data_and_37_enex5 ) begin
      reg_weight_write_data_data_0_2_lpi_1_dfm_1_1_enexo <= while_if_and_14_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_1_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_14_cse | weight_write_data_data_and_38_enex5 ) begin
      reg_weight_write_data_data_0_1_lpi_1_dfm_1_1_enexo <= while_if_and_14_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_write_data_data_0_0_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_14_cse | weight_write_data_data_and_39_enex5 ) begin
      reg_weight_write_data_data_0_0_lpi_1_dfm_1_1_enexo <= while_if_and_14_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_pe_manager_base_input_enexo <= 1'b1;
    end
    else if ( pe_manager_base_input_and_tmp | weight_write_addrs_and_2_enex5 ) begin
      reg_pe_manager_base_input_enexo <= pe_manager_base_input_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_read_addrs_0_3_0_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_14_cse | weight_read_addrs_and_28_enex5 ) begin
      reg_weight_read_addrs_0_3_0_lpi_1_dfm_1_1_enexo <= while_if_and_14_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_pe_config_num_output_enexo <= 1'b1;
    end
    else if ( pe_config_num_manager_and_cse | pe_config_UpdateManagerCounter_if_if_and_enex5
        ) begin
      reg_pe_config_num_output_enexo <= pe_config_num_manager_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( while_if_and_14_cse | weight_read_addrs_and_29_enex5 ) begin
      reg_weight_read_addrs_0_14_4_lpi_1_dfm_1_1_enexo <= while_if_and_14_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_in_reg_data_sva_1_enexo <= 1'b1;
    end
    else if ( rva_in_reg_data_and_tmp | PEManager_15U_PEManagerWrite_and_enex5 )
        begin
      reg_rva_in_reg_data_sva_1_enexo <= rva_in_reg_data_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0_enexo <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_18_enex5 | input_mem_banks_read_read_data_and_26_enex5
        ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0_enexo <= input_mem_banks_read_read_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0_enexo_1 <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_18_enex5 | input_mem_banks_read_read_data_and_27_enex5
        ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0_enexo_1 <= input_mem_banks_read_read_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0_enexo_2 <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_18_enex5 | input_mem_banks_read_read_data_and_28_enex5
        ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0_enexo_2 <= input_mem_banks_read_read_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0_enexo_3 <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_18_enex5 | input_mem_banks_read_read_data_and_29_enex5
        ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_6_31_0_enexo_3 <= input_mem_banks_read_read_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_2_enexo <= 1'b1;
    end
    else if ( input_mem_banks_read_1_read_data_and_4_enex5 | input_mem_banks_read_1_read_data_and_3_enex5
        ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_2_enexo <= input_mem_banks_read_1_read_data_and_4_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_5_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_91_enex5 | rva_out_reg_data_and_86_enex5 ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_5_enexo <= rva_out_reg_data_and_91_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_5_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_92_enex5 | rva_out_reg_data_and_87_enex5 ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_5_enexo <= rva_out_reg_data_and_92_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_7_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_93_enex5 | rva_out_reg_data_and_88_enex5 ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_7_enexo <= rva_out_reg_data_and_93_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_94_enex5 | rva_out_reg_data_and_89_enex5 ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_4_2_enexo <= rva_out_reg_data_and_94_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_95_enex5 | rva_out_reg_data_and_90_enex5 ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_4_2_enexo <= rva_out_reg_data_and_95_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_5_31_0_enexo <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_19_enex5 | input_mem_banks_read_read_data_and_18_enex5
        ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_5_31_0_enexo <= input_mem_banks_read_read_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_write_arbxbar_xbar_for_empty_sva_1_enexo <= 1'b1;
    end
    else if ( weight_mem_read_arbxbar_xbar_requests_transpose_and_14_cse | weight_mem_write_arbxbar_xbar_for_empty_and_enex5
        ) begin
      reg_weight_mem_write_arbxbar_xbar_for_empty_sva_1_enexo <= weight_mem_read_arbxbar_xbar_requests_transpose_and_14_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( input_mem_banks_read_1_read_data_and_5_enex5 | input_mem_banks_read_1_read_data_and_4_enex5
        ) begin
      reg_input_mem_banks_read_1_read_data_lpi_1_dfm_1_1_enexo <= input_mem_banks_read_1_read_data_and_5_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_run_3_for_5_mux_12_itm_1_1_enexo <= 1'b1;
    end
    else if ( weight_mem_run_3_for_5_and_209_ssc | rva_out_reg_data_and_91_enex5
        ) begin
      reg_weight_mem_run_3_for_5_mux_12_itm_1_1_enexo <= weight_mem_run_3_for_5_and_209_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_run_3_for_5_mux_11_itm_1_1_enexo <= 1'b1;
    end
    else if ( weight_mem_run_3_for_5_and_209_ssc | rva_out_reg_data_and_92_enex5
        ) begin
      reg_weight_mem_run_3_for_5_mux_11_itm_1_1_enexo <= weight_mem_run_3_for_5_and_209_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_mem_run_3_for_5_mux_10_itm_1_1_enexo <= 1'b1;
    end
    else if ( weight_mem_run_3_for_5_and_209_ssc | rva_out_reg_data_and_93_enex5
        ) begin
      reg_weight_mem_run_3_for_5_mux_10_itm_1_1_enexo <= weight_mem_run_3_for_5_and_209_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( and_1402_cse | rva_out_reg_data_and_94_enex5 ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_4_1_enexo <= and_1402_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( and_1402_cse | rva_out_reg_data_and_95_enex5 ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_4_1_enexo <= and_1402_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_167_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1920_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_167_sva_dfm_2_enexo <= and_1920_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_86_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1677_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_86_sva_dfm_2_enexo <= and_1677_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_242_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2145_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_242_sva_dfm_2_enexo <= and_2145_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_165_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1914_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_165_sva_dfm_2_enexo <= and_1914_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_186_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1977_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_186_sva_dfm_2_enexo <= and_1977_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_110_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1749_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_110_sva_dfm_2_enexo <= and_1749_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_187_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1980_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_187_sva_dfm_2_enexo <= and_1980_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_246_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2157_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_246_sva_dfm_2_enexo <= and_2157_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_129_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1806_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_129_sva_dfm_2_enexo <= and_1806_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_175_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1944_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_175_sva_dfm_2_enexo <= and_1944_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_239_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2136_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_239_sva_dfm_2_enexo <= and_2136_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_227_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2100_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_227_sva_dfm_2_enexo <= and_2100_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_138_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1833_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_138_sva_dfm_2_enexo <= and_1833_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_174_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1941_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_174_sva_dfm_2_enexo <= and_1941_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_11_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1452_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_11_sva_dfm_2_enexo <= and_1452_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_79_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1656_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_79_sva_dfm_2_enexo <= and_1656_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_71_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1632_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_71_sva_dfm_2_enexo <= and_1632_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_82_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1665_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_82_sva_dfm_2_enexo <= and_1665_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_97_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1710_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_97_sva_dfm_2_enexo <= and_1710_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_188_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1983_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_188_sva_dfm_2_enexo <= and_1983_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_162_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1905_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_162_sva_dfm_2_enexo <= and_1905_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_205_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2034_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_205_sva_dfm_2_enexo <= and_2034_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_93_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1698_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_93_sva_dfm_2_enexo <= and_1698_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_54_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1581_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_54_sva_dfm_2_enexo <= and_1581_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_38_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1533_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_38_sva_dfm_2_enexo <= and_1533_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_192_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1995_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_192_sva_dfm_2_enexo <= and_1995_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_209_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2046_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_209_sva_dfm_2_enexo <= and_2046_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_220_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2079_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_220_sva_dfm_2_enexo <= and_2079_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_139_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1836_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_139_sva_dfm_2_enexo <= and_1836_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_196_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2007_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_196_sva_dfm_2_enexo <= and_2007_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_207_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2040_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_207_sva_dfm_2_enexo <= and_2040_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_224_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2091_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_224_sva_dfm_2_enexo <= and_2091_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_204_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2031_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_204_sva_dfm_2_enexo <= and_2031_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_write_req_valid_lpi_1_dfm_1_1_enexo <= 1'b1;
    end
    else if ( rva_in_reg_rw_and_6_cse | input_mem_banks_read_1_read_data_and_5_enex5
        ) begin
      reg_input_write_req_valid_lpi_1_dfm_1_1_enexo <= rva_in_reg_rw_and_6_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_51_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1572_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_51_sva_dfm_2_enexo <= and_1572_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_72_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1635_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_72_sva_dfm_2_enexo <= and_1635_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_111_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1752_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_111_sva_dfm_2_enexo <= and_1752_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_2_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1425_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_2_sva_dfm_2_enexo <= and_1425_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_99_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1716_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_99_sva_dfm_2_enexo <= and_1716_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_65_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1614_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_65_sva_dfm_2_enexo <= and_1614_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_101_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1722_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_101_sva_dfm_2_enexo <= and_1722_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_52_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1575_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_52_sva_dfm_2_enexo <= and_1575_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_182_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1965_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_182_sva_dfm_2_enexo <= and_1965_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_109_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1746_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_109_sva_dfm_2_enexo <= and_1746_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_60_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1599_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_60_sva_dfm_2_enexo <= and_1599_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_83_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1668_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_83_sva_dfm_2_enexo <= and_1668_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_214_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2061_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_214_sva_dfm_2_enexo <= and_2061_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_33_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1518_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_33_sva_dfm_2_enexo <= and_1518_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_23_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1488_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_23_sva_dfm_2_enexo <= and_1488_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_173_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1938_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_173_sva_dfm_2_enexo <= and_1938_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_141_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1842_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_141_sva_dfm_2_enexo <= and_1842_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_114_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1761_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_114_sva_dfm_2_enexo <= and_1761_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_236_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2127_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_236_sva_dfm_2_enexo <= and_2127_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_238_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2133_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_238_sva_dfm_2_enexo <= and_2133_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_151_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1872_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_151_sva_dfm_2_enexo <= and_1872_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_243_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2148_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_243_sva_dfm_2_enexo <= and_2148_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_245_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2154_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_245_sva_dfm_2_enexo <= and_2154_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_131_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1812_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_131_sva_dfm_2_enexo <= and_1812_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_94_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1701_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_94_sva_dfm_2_enexo <= and_1701_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_226_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2097_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_226_sva_dfm_2_enexo <= and_2097_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_168_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1923_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_168_sva_dfm_2_enexo <= and_1923_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_26_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1497_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_26_sva_dfm_2_enexo <= and_1497_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_124_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1791_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_124_sva_dfm_2_enexo <= and_1791_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_45_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1554_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_45_sva_dfm_2_enexo <= and_1554_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_89_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1686_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_89_sva_dfm_2_enexo <= and_1686_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_75_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1644_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_75_sva_dfm_2_enexo <= and_1644_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_163_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1908_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_163_sva_dfm_2_enexo <= and_1908_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_61_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1602_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_61_sva_dfm_2_enexo <= and_1602_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_13_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1458_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_13_sva_dfm_2_enexo <= and_1458_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_62_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1605_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_62_sva_dfm_2_enexo <= and_1605_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_32_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1515_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_32_sva_dfm_2_enexo <= and_1515_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_6_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1437_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_6_sva_dfm_2_enexo <= and_1437_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_210_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2049_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_210_sva_dfm_2_enexo <= and_2049_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_31_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1512_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_31_sva_dfm_2_enexo <= and_1512_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_118_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1773_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_118_sva_dfm_2_enexo <= and_1773_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_230_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2109_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_230_sva_dfm_2_enexo <= and_2109_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_250_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2169_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_250_sva_dfm_2_enexo <= and_2169_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_217_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2070_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_217_sva_dfm_2_enexo <= and_2070_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_253_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2178_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_253_sva_dfm_2_enexo <= and_2178_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_212_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2055_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_212_sva_dfm_2_enexo <= and_2055_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_132_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1815_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_132_sva_dfm_2_enexo <= and_1815_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_43_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1548_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_43_sva_dfm_2_enexo <= and_1548_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_160_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1899_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_160_sva_dfm_2_enexo <= and_1899_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_42_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1545_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_42_sva_dfm_2_enexo <= and_1545_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_85_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1674_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_85_sva_dfm_2_enexo <= and_1674_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_4_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1431_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_4_sva_dfm_2_enexo <= and_1431_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_16_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1467_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_16_sva_dfm_2_enexo <= and_1467_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_25_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1494_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_25_sva_dfm_2_enexo <= and_1494_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_46_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1557_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_46_sva_dfm_2_enexo <= and_1557_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_50_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1569_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_50_sva_dfm_2_enexo <= and_1569_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_40_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1539_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_40_sva_dfm_2_enexo <= and_1539_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_117_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1770_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_117_sva_dfm_2_enexo <= and_1770_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_134_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1821_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_134_sva_dfm_2_enexo <= and_1821_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_155_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1884_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_155_sva_dfm_2_enexo <= and_1884_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_254_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2181_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_254_sva_dfm_2_enexo <= and_2181_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_17_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1470_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_17_sva_dfm_2_enexo <= and_1470_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_208_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2043_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_208_sva_dfm_2_enexo <= and_2043_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_185_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1974_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_185_sva_dfm_2_enexo <= and_1974_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_219_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2076_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_219_sva_dfm_2_enexo <= and_2076_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_125_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1794_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_125_sva_dfm_2_enexo <= and_1794_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_68_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1623_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_68_sva_dfm_2_enexo <= and_1623_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_24_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1491_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_24_sva_dfm_2_enexo <= and_1491_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_12_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1455_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_12_sva_dfm_2_enexo <= and_1455_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_59_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1596_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_59_sva_dfm_2_enexo <= and_1596_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_199_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2016_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_199_sva_dfm_2_enexo <= and_2016_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_156_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1887_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_156_sva_dfm_2_enexo <= and_1887_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_77_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1650_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_77_sva_dfm_2_enexo <= and_1650_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_216_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2067_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_216_sva_dfm_2_enexo <= and_2067_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_34_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1521_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_34_sva_dfm_2_enexo <= and_1521_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_251_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2172_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_251_sva_dfm_2_enexo <= and_2172_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_228_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2103_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_228_sva_dfm_2_enexo <= and_2103_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_78_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1653_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_78_sva_dfm_2_enexo <= and_1653_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_67_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1620_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_67_sva_dfm_2_enexo <= and_1620_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_19_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1476_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_19_sva_dfm_2_enexo <= and_1476_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_27_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1500_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_27_sva_dfm_2_enexo <= and_1500_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_81_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1662_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_81_sva_dfm_2_enexo <= and_1662_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_164_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1911_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_164_sva_dfm_2_enexo <= and_1911_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_183_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1968_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_183_sva_dfm_2_enexo <= and_1968_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_179_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1956_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_179_sva_dfm_2_enexo <= and_1956_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_189_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1986_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_189_sva_dfm_2_enexo <= and_1986_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_213_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2058_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_213_sva_dfm_2_enexo <= and_2058_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_234_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2121_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_234_sva_dfm_2_enexo <= and_2121_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_248_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2163_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_248_sva_dfm_2_enexo <= and_2163_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_249_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2166_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_249_sva_dfm_2_enexo <= and_2166_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_112_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1755_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_112_sva_dfm_2_enexo <= and_1755_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_232_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2115_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_232_sva_dfm_2_enexo <= and_2115_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_read_addrs_sva_1_1_enexo <= 1'b1;
    end
    else if ( PECoreRun_wen | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_read_addrs_sva_1_1_enexo <= PECoreRun_wen;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_181_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1962_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_181_sva_dfm_2_enexo <= and_1962_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_18_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1473_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_18_sva_dfm_2_enexo <= and_1473_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_218_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2073_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_218_sva_dfm_2_enexo <= and_2073_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_80_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1659_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_80_sva_dfm_2_enexo <= and_1659_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_121_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1782_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_121_sva_dfm_2_enexo <= and_1782_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_15_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1464_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_15_sva_dfm_2_enexo <= and_1464_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_92_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1695_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_92_sva_dfm_2_enexo <= and_1695_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_152_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1875_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_152_sva_dfm_2_enexo <= and_1875_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_203_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2028_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_203_sva_dfm_2_enexo <= and_2028_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_0_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1419_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_0_sva_dfm_2_enexo <= and_1419_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_44_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1551_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_44_sva_dfm_2_enexo <= and_1551_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_237_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2130_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_237_sva_dfm_2_enexo <= and_2130_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_105_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1734_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_105_sva_dfm_2_enexo <= and_1734_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_84_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1671_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_84_sva_dfm_2_enexo <= and_1671_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_193_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1998_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_193_sva_dfm_2_enexo <= and_1998_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_225_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2094_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_225_sva_dfm_2_enexo <= and_2094_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_21_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1482_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_21_sva_dfm_2_enexo <= and_1482_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_143_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1848_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_143_sva_dfm_2_enexo <= and_1848_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_57_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1590_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_57_sva_dfm_2_enexo <= and_1590_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_154_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1881_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_154_sva_dfm_2_enexo <= and_1881_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_63_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1608_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_63_sva_dfm_2_enexo <= and_1608_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_106_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1737_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_106_sva_dfm_2_enexo <= and_1737_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_87_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1680_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_87_sva_dfm_2_enexo <= and_1680_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_177_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1950_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_177_sva_dfm_2_enexo <= and_1950_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_201_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2022_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_201_sva_dfm_2_enexo <= and_2022_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_122_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1785_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_122_sva_dfm_2_enexo <= and_1785_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_113_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1758_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_113_sva_dfm_2_enexo <= and_1758_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_88_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1683_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_88_sva_dfm_2_enexo <= and_1683_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_74_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1641_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_74_sva_dfm_2_enexo <= and_1641_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_90_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1689_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_90_sva_dfm_2_enexo <= and_1689_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_41_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1542_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_41_sva_dfm_2_enexo <= and_1542_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_7_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1440_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_7_sva_dfm_2_enexo <= and_1440_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_235_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2124_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_235_sva_dfm_2_enexo <= and_2124_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_126_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1797_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_126_sva_dfm_2_enexo <= and_1797_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_146_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1857_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_146_sva_dfm_2_enexo <= and_1857_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_229_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2106_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_229_sva_dfm_2_enexo <= and_2106_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_223_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2088_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_223_sva_dfm_2_enexo <= and_2088_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_161_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1902_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_161_sva_dfm_2_enexo <= and_1902_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_206_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2037_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_206_sva_dfm_2_enexo <= and_2037_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_130_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1809_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_130_sva_dfm_2_enexo <= and_1809_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_195_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2004_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_195_sva_dfm_2_enexo <= and_2004_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_sva_1_enexo <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_21_tmp | input_mem_banks_read_1_read_data_and_5_enex5
        ) begin
      reg_input_mem_banks_read_read_data_sva_1_enexo <= input_mem_banks_read_read_data_and_21_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_103_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1728_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_103_sva_dfm_2_enexo <= and_1728_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_100_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1719_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_100_sva_dfm_2_enexo <= and_1719_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_157_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1890_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_157_sva_dfm_2_enexo <= and_1890_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_127_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1800_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_127_sva_dfm_2_enexo <= and_1800_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_49_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1566_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_49_sva_dfm_2_enexo <= and_1566_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_47_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1560_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_47_sva_dfm_2_enexo <= and_1560_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_240_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2139_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_240_sva_dfm_2_enexo <= and_2139_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_222_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2085_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_222_sva_dfm_2_enexo <= and_2085_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_120_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1779_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_120_sva_dfm_2_enexo <= and_1779_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_66_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1617_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_66_sva_dfm_2_enexo <= and_1617_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_35_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1524_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_35_sva_dfm_2_enexo <= and_1524_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_133_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1818_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_133_sva_dfm_2_enexo <= and_1818_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_172_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1935_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_172_sva_dfm_2_enexo <= and_1935_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_69_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1626_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_69_sva_dfm_2_enexo <= and_1626_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_108_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1743_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_108_sva_dfm_2_enexo <= and_1743_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_14_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1461_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_14_sva_dfm_2_enexo <= and_1461_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_159_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1896_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_159_sva_dfm_2_enexo <= and_1896_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_76_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1647_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_76_sva_dfm_2_enexo <= and_1647_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_241_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2142_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_241_sva_dfm_2_enexo <= and_2142_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_171_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1932_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_171_sva_dfm_2_enexo <= and_1932_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_200_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2019_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_200_sva_dfm_2_enexo <= and_2019_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_98_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1713_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_98_sva_dfm_2_enexo <= and_1713_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_233_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2118_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_233_sva_dfm_2_enexo <= and_2118_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_148_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1863_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_148_sva_dfm_2_enexo <= and_1863_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_104_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1731_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_104_sva_dfm_2_enexo <= and_1731_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_55_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1584_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_55_sva_dfm_2_enexo <= and_1584_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_123_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1788_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_123_sva_dfm_2_enexo <= and_1788_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_119_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1776_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_119_sva_dfm_2_enexo <= and_1776_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_135_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1824_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_135_sva_dfm_2_enexo <= and_1824_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_116_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1767_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_116_sva_dfm_2_enexo <= and_1767_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_128_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1803_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_128_sva_dfm_2_enexo <= and_1803_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_194_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2001_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_194_sva_dfm_2_enexo <= and_2001_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_30_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1509_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_30_sva_dfm_2_enexo <= and_1509_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_136_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1827_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_136_sva_dfm_2_enexo <= and_1827_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_255_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2184_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_255_sva_dfm_2_enexo <= and_2184_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_221_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2082_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_221_sva_dfm_2_enexo <= and_2082_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_244_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2151_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_244_sva_dfm_2_enexo <= and_2151_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_28_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1503_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_28_sva_dfm_2_enexo <= and_1503_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_231_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2112_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_231_sva_dfm_2_enexo <= and_2112_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_180_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1959_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_180_sva_dfm_2_enexo <= and_1959_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_145_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1854_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_145_sva_dfm_2_enexo <= and_1854_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_150_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1869_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_150_sva_dfm_2_enexo <= and_1869_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_96_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1707_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_96_sva_dfm_2_enexo <= and_1707_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_140_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1839_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_140_sva_dfm_2_enexo <= and_1839_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_8_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1443_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_8_sva_dfm_2_enexo <= and_1443_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_91_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1692_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_91_sva_dfm_2_enexo <= and_1692_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_202_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2025_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_202_sva_dfm_2_enexo <= and_2025_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_20_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1479_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_20_sva_dfm_2_enexo <= and_1479_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_169_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1926_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_169_sva_dfm_2_enexo <= and_1926_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_176_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1947_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_176_sva_dfm_2_enexo <= and_1947_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_158_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1893_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_158_sva_dfm_2_enexo <= and_1893_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_149_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1866_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_149_sva_dfm_2_enexo <= and_1866_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_147_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1860_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_147_sva_dfm_2_enexo <= and_1860_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_53_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1578_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_53_sva_dfm_2_enexo <= and_1578_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_29_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1506_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_29_sva_dfm_2_enexo <= and_1506_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_153_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1878_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_153_sva_dfm_2_enexo <= and_1878_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_252_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2175_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_252_sva_dfm_2_enexo <= and_2175_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_3_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1428_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_3_sva_dfm_2_enexo <= and_1428_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_102_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1725_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_102_sva_dfm_2_enexo <= and_1725_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_107_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1740_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_107_sva_dfm_2_enexo <= and_1740_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_9_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1446_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_9_sva_dfm_2_enexo <= and_1446_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_137_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1830_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_137_sva_dfm_2_enexo <= and_1830_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_115_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1764_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_115_sva_dfm_2_enexo <= and_1764_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_170_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1929_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_170_sva_dfm_2_enexo <= and_1929_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_211_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2052_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_211_sva_dfm_2_enexo <= and_2052_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_10_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1449_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_10_sva_dfm_2_enexo <= and_1449_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_197_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2010_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_197_sva_dfm_2_enexo <= and_2010_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_64_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1611_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_64_sva_dfm_2_enexo <= and_1611_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_166_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1917_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_166_sva_dfm_2_enexo <= and_1917_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_191_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1992_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_191_sva_dfm_2_enexo <= and_1992_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_198_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2013_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_198_sva_dfm_2_enexo <= and_2013_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_190_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1989_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_190_sva_dfm_2_enexo <= and_1989_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_5_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1434_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_5_sva_dfm_2_enexo <= and_1434_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_184_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1971_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_184_sva_dfm_2_enexo <= and_1971_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_215_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2064_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_215_sva_dfm_2_enexo <= and_2064_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_37_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1530_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_37_sva_dfm_2_enexo <= and_1530_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_247_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_2160_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_247_sva_dfm_2_enexo <= and_2160_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_36_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1527_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_36_sva_dfm_2_enexo <= and_1527_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_142_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1845_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_142_sva_dfm_2_enexo <= and_1845_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_178_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1953_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_178_sva_dfm_2_enexo <= and_1953_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_73_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1638_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_73_sva_dfm_2_enexo <= and_1638_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_144_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1851_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_144_sva_dfm_2_enexo <= and_1851_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_22_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1485_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_22_sva_dfm_2_enexo <= and_1485_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_48_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1563_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_48_sva_dfm_2_enexo <= and_1563_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_56_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1587_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_56_sva_dfm_2_enexo <= and_1587_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_39_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1536_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_39_sva_dfm_2_enexo <= and_1536_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_58_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1593_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_58_sva_dfm_2_enexo <= and_1593_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_1_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1422_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_1_sva_dfm_2_enexo <= and_1422_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_95_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1704_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_95_sva_dfm_2_enexo <= and_1704_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_bank_a_70_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( and_1629_tmp | input_mem_banks_read_1_read_data_and_5_enex5 ) begin
      reg_input_mem_banks_bank_a_70_sva_dfm_2_enexo <= and_1629_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo <= 1'b1;
    end
    else if ( input_mem_banks_read_read_data_and_20_tmp | input_mem_banks_read_read_data_and_19_enex5
        ) begin
      reg_input_mem_banks_read_read_data_lpi_1_dfm_1_4_enexo <= input_mem_banks_read_read_data_and_20_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_59_cse | rva_out_reg_data_and_96_enex5 ) begin
      reg_rva_out_reg_data_30_25_sva_dfm_1_enexo <= rva_out_reg_data_and_59_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_59_cse | rva_out_reg_data_and_97_enex5 ) begin
      reg_rva_out_reg_data_23_17_sva_dfm_1_enexo <= rva_out_reg_data_and_59_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_104_enex5 | rva_out_reg_data_and_98_enex5 ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_3_enexo <= rva_out_reg_data_and_104_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_1_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_105_enex5 | rva_out_reg_data_and_99_enex5 ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_1_3_enexo <= rva_out_reg_data_and_105_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_1_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_106_enex5 | rva_out_reg_data_and_100_enex5 ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_1_3_enexo <= rva_out_reg_data_and_106_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_1_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_107_enex5 | rva_out_reg_data_and_101_enex5 ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_1_3_enexo <= rva_out_reg_data_and_107_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_1_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_108_enex5 | rva_out_reg_data_and_102_enex5 ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_1_3_enexo <= rva_out_reg_data_and_108_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_1_3_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_109_enex5 | rva_out_reg_data_and_103_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_1_3_enexo <= rva_out_reg_data_and_109_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_67_enex5 | rva_out_reg_data_and_104_enex5 ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_2_enexo <= rva_out_reg_data_and_67_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_1_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_110_enex5 | rva_out_reg_data_and_105_enex5 ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_1_2_enexo <= rva_out_reg_data_and_110_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_1_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_111_enex5 | rva_out_reg_data_and_106_enex5 ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_1_2_enexo <= rva_out_reg_data_and_111_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_1_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_112_enex5 | rva_out_reg_data_and_107_enex5 ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_1_2_enexo <= rva_out_reg_data_and_112_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_1_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_113_enex5 | rva_out_reg_data_and_108_enex5 ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_1_2_enexo <= rva_out_reg_data_and_113_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_1_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_114_enex5 | rva_out_reg_data_and_109_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_1_2_enexo <= rva_out_reg_data_and_114_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_1_enexo <= 1'b1;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_37_cse | rva_out_reg_data_and_67_enex5
        ) begin
      reg_rva_out_reg_data_15_9_sva_dfm_1_enexo <= PECore_DecodeAxiRead_case_4_switch_lp_and_37_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_41_cse | rva_out_reg_data_and_110_enex5
        ) begin
      reg_rva_out_reg_data_35_32_sva_dfm_1_1_enexo <= PECore_DecodeAxiRead_case_4_switch_lp_and_41_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_41_cse | rva_out_reg_data_and_111_enex5
        ) begin
      reg_rva_out_reg_data_39_36_sva_dfm_1_1_enexo <= PECore_DecodeAxiRead_case_4_switch_lp_and_41_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_41_cse | rva_out_reg_data_and_112_enex5
        ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_1_1_enexo <= PECore_DecodeAxiRead_case_4_switch_lp_and_41_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_1_1_enexo <= 1'b1;
    end
    else if ( PECore_DecodeAxiRead_case_4_switch_lp_and_41_cse | rva_out_reg_data_and_113_enex5
        ) begin
      reg_rva_out_reg_data_62_56_sva_dfm_1_1_enexo <= PECore_DecodeAxiRead_case_4_switch_lp_and_41_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_pe_config_input_counter_sva_dfm_1_enexo <= 1'b1;
    end
    else if ( and_1217_tmp | rva_out_reg_data_and_114_enex5 ) begin
      reg_pe_config_input_counter_sva_dfm_1_enexo <= and_1217_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_2_sva_dfm_2_2_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_110_enex5 | weight_port_read_out_data_and_106_enex5
        ) begin
      reg_weight_port_read_out_data_0_2_sva_dfm_2_2_enexo <= weight_port_read_out_data_and_110_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_2_2_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_111_enex5 | weight_port_read_out_data_and_107_enex5
        ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_2_2_enexo <= weight_port_read_out_data_and_111_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_2_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_118_enex5 | rva_out_reg_data_and_115_enex5 ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_2_1_enexo <= rva_out_reg_data_and_118_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_2_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_119_enex5 | rva_out_reg_data_and_116_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_2_enexo <= rva_out_reg_data_and_119_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_2_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_120_enex5 | rva_out_reg_data_and_117_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_2_1_enexo <= rva_out_reg_data_and_120_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_1_2_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_100_ssc | weight_port_read_out_data_and_108_enex5
        ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_1_2_enexo <= weight_port_read_out_data_and_100_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_1_2_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_100_ssc | weight_port_read_out_data_and_109_enex5
        ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_1_2_enexo <= weight_port_read_out_data_and_100_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_2_sva_dfm_1_2_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_100_ssc | weight_port_read_out_data_and_110_enex5
        ) begin
      reg_weight_port_read_out_data_0_2_sva_dfm_1_2_enexo <= weight_port_read_out_data_and_100_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_1_2_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_100_ssc | weight_port_read_out_data_and_111_enex5
        ) begin
      reg_weight_port_read_out_data_0_3_sva_dfm_1_2_enexo <= weight_port_read_out_data_and_100_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_1_1_enexo <= 1'b1;
    end
    else if ( and_1402_cse | rva_out_reg_data_and_118_enex5 ) begin
      reg_rva_out_reg_data_46_40_sva_dfm_4_1_1_enexo <= and_1402_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_1_enexo <= 1'b1;
    end
    else if ( and_1402_cse | rva_out_reg_data_and_119_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_1_enexo <= and_1402_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_1_1_enexo <= 1'b1;
    end
    else if ( and_1402_cse | rva_out_reg_data_and_120_enex5 ) begin
      reg_rva_out_reg_data_55_48_sva_dfm_4_1_1_enexo <= and_1402_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_3_2_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_113_enex5 | weight_port_read_out_data_and_112_enex5
        ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_3_2_enexo <= weight_port_read_out_data_and_113_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_2_2_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_108_enex5 | weight_port_read_out_data_and_113_enex5
        ) begin
      reg_weight_port_read_out_data_0_0_sva_dfm_2_2_enexo <= weight_port_read_out_data_and_108_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_2_2_enexo <= 1'b1;
    end
    else if ( weight_port_read_out_data_and_109_enex5 | weight_port_read_out_data_and_114_enex5
        ) begin
      reg_weight_port_read_out_data_0_1_sva_dfm_2_2_enexo <= weight_port_read_out_data_and_109_enex5;
    end
  end
  assign nl_operator_4_false_acc_nl = pe_config_manager_counter_sva_mx1 + 4'b0001;
  assign operator_4_false_acc_nl = nl_operator_4_false_acc_nl[3:0];
  assign pe_config_UpdateManagerCounter_if_not_7_nl = ~ pe_config_UpdateManagerCounter_pe_config_UpdateManagerCounter_if_nor_svs_1_1;
  assign nl_input_read_addrs_sva_1_1  = pe_config_input_counter_sva_mx1 + pe_manager_base_input_sva_mx1_7_0;
  assign while_if_while_if_and_12_nl = PECore_DecodeAxiRead_switch_lp_equal_tmp_3_mx0w0
      & (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt);
  assign nl_PECore_RunScale_if_for_8_mul_1_nl = $signed(accum_vector_data_7_sva)
      * $signed(9'b010100111);
  assign PECore_RunScale_if_for_8_mul_1_nl = nl_PECore_RunScale_if_for_8_mul_1_nl[30:0];
  assign nl_PECore_RunScale_if_for_1_mul_1_nl = $signed(accum_vector_data_0_sva)
      * $signed(9'b010100111);
  assign PECore_RunScale_if_for_1_mul_1_nl = nl_PECore_RunScale_if_for_1_mul_1_nl[30:0];
  assign nl_PECore_RunScale_if_for_7_mul_1_nl = $signed(accum_vector_data_6_sva)
      * $signed(9'b010100111);
  assign PECore_RunScale_if_for_7_mul_1_nl = nl_PECore_RunScale_if_for_7_mul_1_nl[30:0];
  assign nl_PECore_RunScale_if_for_2_mul_1_nl = $signed(accum_vector_data_1_sva)
      * $signed(9'b010100111);
  assign PECore_RunScale_if_for_2_mul_1_nl = nl_PECore_RunScale_if_for_2_mul_1_nl[30:0];
  assign nl_PECore_RunScale_if_for_6_mul_1_nl = $signed(accum_vector_data_5_sva)
      * $signed(9'b010100111);
  assign PECore_RunScale_if_for_6_mul_1_nl = nl_PECore_RunScale_if_for_6_mul_1_nl[30:0];
  assign nl_PECore_RunScale_if_for_3_mul_1_nl = $signed(accum_vector_data_2_sva)
      * $signed(9'b010100111);
  assign PECore_RunScale_if_for_3_mul_1_nl = nl_PECore_RunScale_if_for_3_mul_1_nl[30:0];
  assign nl_PECore_RunScale_if_for_5_mul_1_nl = $signed(accum_vector_data_4_sva)
      * $signed(9'b010100111);
  assign PECore_RunScale_if_for_5_mul_1_nl = nl_PECore_RunScale_if_for_5_mul_1_nl[30:0];
  assign nl_PECore_RunScale_if_for_4_mul_1_nl = $signed(accum_vector_data_3_sva)
      * $signed(9'b010100111);
  assign PECore_RunScale_if_for_4_mul_1_nl = nl_PECore_RunScale_if_for_4_mul_1_nl[30:0];
  assign accum_vector_data_mux_62_nl = MUX_v_23_2_2(accum_vector_data_7_sva_6_mx1w0,
      accum_vector_data_7_sva_6, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7);
  assign accum_vector_data_mux_59_nl = MUX_v_23_2_2(accum_vector_data_7_sva_7_mx1w0,
      accum_vector_data_7_sva_7, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7);
  assign nl_accum_vector_data_acc_30_itm_1  = accum_vector_data_mux_62_nl + accum_vector_data_mux_59_nl;
  assign accum_vector_data_mux_68_nl = MUX_v_23_2_2(accum_vector_data_6_sva_6_mx1w0,
      accum_vector_data_6_sva_6, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7);
  assign accum_vector_data_mux_65_nl = MUX_v_23_2_2(accum_vector_data_6_sva_7_mx1w0,
      accum_vector_data_6_sva_7, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7);
  assign nl_accum_vector_data_acc_28_itm_1  = accum_vector_data_mux_68_nl + accum_vector_data_mux_65_nl;
  assign accum_vector_data_mux_74_nl = MUX_v_23_2_2(accum_vector_data_5_sva_6_mx1w0,
      accum_vector_data_5_sva_6, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7);
  assign accum_vector_data_mux_71_nl = MUX_v_23_2_2(accum_vector_data_5_sva_7_mx1w0,
      accum_vector_data_5_sva_7, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7);
  assign nl_accum_vector_data_acc_25_itm_1  = accum_vector_data_mux_74_nl + accum_vector_data_mux_71_nl;
  assign accum_vector_data_mux_80_nl = MUX_v_23_2_2(accum_vector_data_4_sva_6_mx1w0,
      accum_vector_data_4_sva_6, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7);
  assign accum_vector_data_mux_77_nl = MUX_v_23_2_2(accum_vector_data_4_sva_7_mx1w0,
      accum_vector_data_4_sva_7, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7);
  assign nl_accum_vector_data_acc_22_itm_1  = accum_vector_data_mux_80_nl + accum_vector_data_mux_77_nl;
  assign accum_vector_data_mux_86_nl = MUX_v_23_2_2(accum_vector_data_3_sva_6_mx1w0,
      accum_vector_data_3_sva_6, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7);
  assign accum_vector_data_mux_83_nl = MUX_v_23_2_2(accum_vector_data_3_sva_7_mx1w0,
      accum_vector_data_3_sva_7, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7);
  assign nl_accum_vector_data_acc_19_itm_1  = accum_vector_data_mux_86_nl + accum_vector_data_mux_83_nl;
  assign accum_vector_data_mux_92_nl = MUX_v_23_2_2(accum_vector_data_1_sva_6_mx1w0,
      accum_vector_data_1_sva_6, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7);
  assign accum_vector_data_mux_89_nl = MUX_v_23_2_2(accum_vector_data_1_sva_7_mx1w0,
      accum_vector_data_1_sva_7, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7);
  assign nl_accum_vector_data_acc_13_itm_1  = accum_vector_data_mux_92_nl + accum_vector_data_mux_89_nl;
  assign accum_vector_data_mux_98_nl = MUX_v_23_2_2(accum_vector_data_0_sva_6_mx1w0,
      accum_vector_data_0_sva_6, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7);
  assign accum_vector_data_mux_95_nl = MUX_v_23_2_2(accum_vector_data_0_sva_7_mx1w0,
      accum_vector_data_0_sva_7, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7);
  assign nl_accum_vector_data_acc_10_itm_1  = accum_vector_data_mux_98_nl + accum_vector_data_mux_95_nl;
  assign mux_6_nl = MUX_s_1_2_2(or_tmp_5, and_tmp, weight_mem_run_3_for_land_3_lpi_1_dfm_1);
  assign or_21_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_63_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_78_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_68_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_for_and_49_tmp | nor_tmp_1;
  assign mux_7_nl = MUX_s_1_2_2(weight_mem_run_3_for_land_5_lpi_1_dfm_1, or_21_nl,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign or_22_nl = (~ weight_mem_run_3_for_land_7_lpi_1_dfm_1) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4;
  assign mux_8_nl = MUX_s_1_2_2(or_tmp_5, and_tmp, weight_mem_run_3_for_land_7_lpi_1_dfm_1);
  assign mux_9_nl = MUX_s_1_2_2(or_22_nl, mux_8_nl, PECore_DecodeAxiRead_switch_lp_equal_tmp_1_3);
  assign weight_mem_run_3_for_5_and_100_nl = (weight_read_addrs_7_lpi_1_dfm_2_2_0==3'b011)
      & weight_mem_run_3_for_land_lpi_1_dfm_1;
  assign mux_10_nl = MUX_s_1_2_2(weight_mem_run_3_for_land_4_lpi_1_dfm_1, (~ rva_in_reg_rw_sva_st_1_4),
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_20_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2==3'b011)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_6_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2==3'b101)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_15_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2==3'b110)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_16_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2==3'b111)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_1;
  assign or_1483_nl = reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_6_cse
      | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_5_cse | reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_4_cse
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_3 | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_2
      | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_1 | Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_0
      | mux_tmp_483;
  assign mux_511_nl = MUX_s_1_2_2(mux_tmp_483, or_1483_nl, Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1);
  assign or_1485_nl = (~ while_stage_0_5) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | (~(Arbiter_8U_Roundrobin_pick_return_1_0_lpi_1_dfm_1_1 | Arbiter_8U_Roundrobin_pick_return_1_0_7_lpi_1_dfm_1_1
      | Arbiter_8U_Roundrobin_pick_return_1_0_6_lpi_1_dfm_1_1 | Arbiter_8U_Roundrobin_pick_return_1_0_5_lpi_1_dfm_1_1
      | Arbiter_8U_Roundrobin_pick_return_1_0_4_lpi_1_dfm_1_1 | Arbiter_8U_Roundrobin_pick_return_1_0_3_lpi_1_dfm_1_1
      | Arbiter_8U_Roundrobin_pick_return_1_0_2_lpi_1_dfm_1_1 | Arbiter_8U_Roundrobin_pick_return_1_0_1_lpi_1_dfm_1_1
      | mux_511_nl));
  assign or_1466_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | (~(weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_1_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1));
  assign mux_512_nl = MUX_s_1_2_2(or_1485_nl, or_1466_nl, while_stage_0_6);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_123_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_24_nl
      = MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[7:0]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_123_nl);
  assign nor_331_nl = ~(weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | (~ weight_mem_read_arbxbar_xbar_1_for_3_3_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1)
      | weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
  assign mux_12_nl = MUX_s_1_2_2(nor_331_nl, crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_44_itm_1,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_109_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_40_nl
      = MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[7:0]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_109_nl);
  assign nor_332_nl = ~(weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | (~ weight_mem_read_arbxbar_xbar_1_for_3_5_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1)
      | weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
  assign mux_13_nl = MUX_s_1_2_2(nor_332_nl, crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_76_itm_1,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign or_32_nl = (~ weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp)
      | (~ while_stage_0_5) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3;
  assign or_31_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | (~ weight_mem_read_arbxbar_xbar_1_for_3_8_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
  assign mux_14_nl = MUX_s_1_2_2(or_32_nl, or_31_nl, while_stage_0_6);
  assign or_34_nl = (~ weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_tmp)
      | (~ while_stage_0_5) | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3;
  assign or_33_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      | (~ weight_mem_read_arbxbar_xbar_1_for_3_7_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
  assign mux_15_nl = MUX_s_1_2_2(or_34_nl, or_33_nl, while_stage_0_6);
  assign mux_16_nl = MUX_s_1_2_2(PECore_RunMac_PECore_RunMac_if_and_svs_st_3, ProductSum_for_asn_25_itm_3,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign nor_900_nl = ~((~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17])
      | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt) | (~ reg_rva_in_PopNB_mioi_iswt0_cse)
      | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[15]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[14])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[13]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[12])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[10])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[9]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[8])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]));
  assign nor_901_nl = ~((~ PECore_DecodeAxiWrite_case_4_switch_lp_equal_tmp_1_1)
      | PECore_DecodeAxiWrite_switch_lp_equal_tmp_1 | PECore_DecodeAxiWrite_switch_lp_nor_tmp_1
      | PECore_DecodeAxiWrite_switch_lp_equal_tmp_2 | nand_372_cse);
  assign mux_513_nl = MUX_s_1_2_2(nor_900_nl, nor_901_nl, while_stage_0_3);
  assign mux_514_nl = MUX_s_1_2_2(mux_513_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2,
      while_stage_0_4);
  assign PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_6_nl
      = MUX_v_11_2_2(11'b00000000000, PEManager_15U_GetWeightAddr_else_acc_2_psp_sva_1,
      PECore_DecodeAxiRead_switch_lp_equal_tmp_2_2);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_49_nl = weight_mem_read_arbxbar_arbiters_next_7_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[7]);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_42_nl = weight_mem_read_arbxbar_arbiters_next_6_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[6]);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_35_nl = weight_mem_read_arbxbar_arbiters_next_5_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[5]);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_28_nl = weight_mem_read_arbxbar_arbiters_next_4_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[4]);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_21_nl = weight_mem_read_arbxbar_arbiters_next_3_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[3]);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_14_nl = weight_mem_read_arbxbar_arbiters_next_2_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[2]);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_7_nl = weight_mem_read_arbxbar_arbiters_next_1_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[1]);
  assign Arbiter_8U_Roundrobin_pick_Arbiter_8U_Roundrobin_pick_or_nl = weight_mem_read_arbxbar_arbiters_next_0_7_sva_mx0
      | (weight_mem_read_arbxbar_xbar_for_1_lshift_tmp[0]);
  assign PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_and_nl
      = MUX_v_4_2_2(4'b0000, pe_config_manager_counter_sva_mx1, PECore_DecodeAxiWrite_case_4_switch_lp_or_cse_1);
  assign and_601_nl = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[18]) & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[19]))
      & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16])) & rva_in_PopNB_mioi_return_rsc_z_mxwt
      & and_dcpl_211 & (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[17]));
  assign PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_or_nl = (state_mux_1_cse!=2'b00)
      | state_0_sva_mx1;
  assign PECore_UpdateFSM_switch_lp_or_nl = PECore_UpdateFSM_switch_lp_equal_tmp_6
      | PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_and_1_cse_1;
  assign PECore_UpdateFSM_switch_lp_mux1h_18_nl = MUX1HOT_v_2_3_2((signext_2_1(PECore_UpdateFSM_switch_lp_PECore_UpdateFSM_switch_lp_or_nl)),
      2'b01, 2'b10, {PECore_RunFSM_switch_lp_PECore_RunFSM_switch_lp_nor_1_cse_1
      , PECore_UpdateFSM_switch_lp_or_nl , PECore_RunScale_PECore_RunScale_if_and_1_svs_1});
  assign PECore_UpdateFSM_switch_lp_nor_8_nl = ~(PECore_PushOutput_PECore_PushOutput_if_and_svs_1
      | PECore_UpdateFSM_switch_lp_nor_tmp_1);
  assign PECore_UpdateFSM_switch_lp_and_1_nl = MUX_v_2_2_2(2'b00, PECore_UpdateFSM_switch_lp_mux1h_18_nl,
      PECore_UpdateFSM_switch_lp_nor_8_nl);
  assign mux_515_nl = MUX_s_1_2_2(PECore_UpdateFSM_switch_lp_equal_tmp_3_1, nor_912_cse,
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign mux_516_nl = MUX_s_1_2_2(and_2257_cse, nor_912_cse, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1);
  assign nl_operator_8_false_acc_sdt_sva_1  = conv_u2s_8_9(pe_config_num_output_sva)
      + 9'b111111111;
  assign accum_vector_data_mux_12_nl = MUX_v_23_2_2(accum_vector_data_7_sva_4_mx0w0,
      accum_vector_data_7_sva_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign accum_vector_data_mux_9_nl = MUX_v_23_2_2(accum_vector_data_7_sva_5_mx1w0,
      accum_vector_data_7_sva_5, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign nl_accum_vector_data_acc_29_nl = accum_vector_data_mux_12_nl + accum_vector_data_mux_9_nl;
  assign accum_vector_data_acc_29_nl = nl_accum_vector_data_acc_29_nl[22:0];
  assign nl_accum_vector_data_7_sva  = accum_vector_data_acc_29_nl + accum_vector_data_acc_30_itm_1;
  assign accum_vector_data_mux_54_nl = MUX_v_23_2_2(accum_vector_data_0_sva_4_mx1w0,
      accum_vector_data_0_sva_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign accum_vector_data_mux_51_nl = MUX_v_23_2_2(accum_vector_data_0_sva_5_mx1w0,
      accum_vector_data_0_sva_5, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign nl_accum_vector_data_acc_9_nl = accum_vector_data_mux_54_nl + accum_vector_data_mux_51_nl;
  assign accum_vector_data_acc_9_nl = nl_accum_vector_data_acc_9_nl[22:0];
  assign nl_accum_vector_data_0_sva  = accum_vector_data_acc_9_nl + accum_vector_data_acc_10_itm_1;
  assign accum_vector_data_mux_17_nl = MUX_v_23_2_2(accum_vector_data_6_sva_4_mx0w0,
      accum_vector_data_6_sva_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign accum_vector_data_mux_14_nl = MUX_v_23_2_2(accum_vector_data_6_sva_5_mx1w0,
      accum_vector_data_6_sva_5, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign nl_accum_vector_data_acc_27_nl = accum_vector_data_mux_17_nl + accum_vector_data_mux_14_nl;
  assign accum_vector_data_acc_27_nl = nl_accum_vector_data_acc_27_nl[22:0];
  assign nl_accum_vector_data_6_sva  = accum_vector_data_acc_27_nl + accum_vector_data_acc_28_itm_1;
  assign accum_vector_data_mux_48_nl = MUX_v_23_2_2(accum_vector_data_1_sva_4_mx1w0,
      accum_vector_data_1_sva_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign accum_vector_data_mux_45_nl = MUX_v_23_2_2(accum_vector_data_1_sva_5_mx1w0,
      accum_vector_data_1_sva_5, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign nl_accum_vector_data_acc_12_nl = accum_vector_data_mux_48_nl + accum_vector_data_mux_45_nl;
  assign accum_vector_data_acc_12_nl = nl_accum_vector_data_acc_12_nl[22:0];
  assign nl_accum_vector_data_1_sva  = accum_vector_data_acc_12_nl + accum_vector_data_acc_13_itm_1;
  assign accum_vector_data_mux_21_nl = MUX_v_23_2_2(accum_vector_data_5_sva_4_mx1w0,
      accum_vector_data_5_sva_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign accum_vector_data_mux_19_nl = MUX_v_23_2_2(accum_vector_data_5_sva_5_mx0w0,
      accum_vector_data_5_sva_5, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign nl_accum_vector_data_acc_24_nl = accum_vector_data_mux_21_nl + accum_vector_data_mux_19_nl;
  assign accum_vector_data_acc_24_nl = nl_accum_vector_data_acc_24_nl[22:0];
  assign nl_accum_vector_data_5_sva  = accum_vector_data_acc_24_nl + accum_vector_data_acc_25_itm_1;
  assign accum_vector_data_mux_42_nl = MUX_v_23_2_2(accum_vector_data_2_sva_4_mx1w0,
      accum_vector_data_2_sva_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign accum_vector_data_mux_39_nl = MUX_v_23_2_2(accum_vector_data_2_sva_5_mx1w0,
      accum_vector_data_2_sva_5, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign nl_accum_vector_data_acc_15_nl = accum_vector_data_mux_42_nl + accum_vector_data_mux_39_nl;
  assign accum_vector_data_acc_15_nl = nl_accum_vector_data_acc_15_nl[22:0];
  assign accum_vector_data_mux_36_nl = MUX_v_23_2_2(accum_vector_data_2_sva_6_mx1w0,
      accum_vector_data_2_sva_6, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign nl_accum_vector_data_acc_16_nl = accum_vector_data_mux_36_nl + accum_vector_data_2_sva_7;
  assign accum_vector_data_acc_16_nl = nl_accum_vector_data_acc_16_nl[22:0];
  assign nl_accum_vector_data_2_sva  = accum_vector_data_acc_15_nl + accum_vector_data_acc_16_nl;
  assign accum_vector_data_mux_27_nl = MUX_v_23_2_2(accum_vector_data_4_sva_4_mx1w0,
      accum_vector_data_4_sva_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign accum_vector_data_mux_24_nl = MUX_v_23_2_2(accum_vector_data_4_sva_5_mx1w0,
      accum_vector_data_4_sva_5, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign nl_accum_vector_data_acc_21_nl = accum_vector_data_mux_27_nl + accum_vector_data_mux_24_nl;
  assign accum_vector_data_acc_21_nl = nl_accum_vector_data_acc_21_nl[22:0];
  assign nl_accum_vector_data_4_sva  = accum_vector_data_acc_21_nl + accum_vector_data_acc_22_itm_1;
  assign accum_vector_data_mux_33_nl = MUX_v_23_2_2(accum_vector_data_3_sva_4_mx1w0,
      accum_vector_data_3_sva_4, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign accum_vector_data_mux_30_nl = MUX_v_23_2_2(accum_vector_data_3_sva_5_mx1w0,
      accum_vector_data_3_sva_5, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_8);
  assign nl_accum_vector_data_acc_18_nl = accum_vector_data_mux_33_nl + accum_vector_data_mux_30_nl;
  assign accum_vector_data_acc_18_nl = nl_accum_vector_data_acc_18_nl[22:0];
  assign nl_accum_vector_data_3_sva  = accum_vector_data_acc_18_nl + accum_vector_data_acc_19_itm_1;
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_122_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_125_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_128_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_76_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_108_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_111_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_112_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_114_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_130_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_134_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_20_nl
      = pe_manager_base_input_sva_mx1_7_0 & ({{7{and_321_cse}}, and_321_cse}) & ({{7{PECore_DecodeAxiRead_switch_lp_nor_13_cse_1}},
      PECore_DecodeAxiRead_switch_lp_nor_13_cse_1});
  assign PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_and_1_nl
      = MUX_v_8_2_2(8'b00000000, pe_config_input_counter_sva_mx1, PECore_DecodeAxiWrite_case_4_switch_lp_or_cse_1);
  assign PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_mux_6_nl
      = MUX_s_1_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[8]), pe_config_is_zero_first_sva_mx1,
      PECore_DecodeAxiWrite_case_4_switch_lp_or_cse_1);
  assign PECore_DecodeAxiWrite_switch_lp_PECore_DecodeAxiWrite_switch_lp_mux_19_nl
      = MUX_s_1_2_2(PECore_DecodeAxiWrite_case_4_switch_lp_PECore_DecodeAxiWrite_case_4_switch_lp_mux_6_nl,
      pe_config_is_zero_first_sva_mx1, PECore_DecodeAxiWrite_switch_lp_or_5_cse_1);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_crossbar_spec_PE_Weight_WordType_8U_8U_for_nor_1_nl
      = ~((crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1!=3'b000));
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_and_7_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1==3'b101)
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_and_9_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1==3'b111)
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_7_nl = (weight_read_addrs_1_lpi_1_dfm_1[2:0]==3'b110)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_1_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_and_16_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1==3'b110)
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_14_nl = (weight_read_addrs_1_lpi_1_dfm_1[2:0]==3'b101)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_1_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_4_nl = (weight_read_addrs_1_lpi_1_dfm_1[2:0]==3'b011)
      & weight_mem_run_3_for_land_2_lpi_1_dfm_1_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_for_and_5_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_1==3'b011)
      & crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_28_nl = (pe_manager_base_weight_sva[2])
      & pe_manager_base_weight_slc_pe_manager_base_weight_2_0_122_itm_1 & (pe_manager_base_weight_sva[0])
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_35_nl = pe_manager_base_weight_slc_pe_manager_base_weight_2_0_95_itm_1
      & (pe_manager_base_weight_sva[1:0]==2'b10) & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_34_nl = (pe_manager_base_weight_sva[2])
      & pe_manager_base_weight_slc_pe_manager_base_weight_2_0_93_itm_1 & (~ (pe_manager_base_weight_sva[1]))
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_26_nl = pe_manager_base_weight_slc_pe_manager_base_weight_2_0_95_itm_1
      & pe_manager_base_weight_slc_pe_manager_base_weight_2_0_93_itm_1 & (~ (pe_manager_base_weight_sva[1]))
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_24_nl = (pe_manager_base_weight_sva[1])
      & pe_manager_base_weight_slc_pe_manager_base_weight_2_0_93_itm_1 & (~ (pe_manager_base_weight_sva[2]))
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign nor_338_nl = ~(while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3
      | mux_tmp_25);
  assign mux_30_nl = MUX_s_1_2_2(or_tmp_43, nor_338_nl, weight_mem_read_arbxbar_xbar_requests_transpose_slc_weight_mem_read_arbxbar_xbar_requests_transpose_0_6_1_itm_1);
  assign mux_31_nl = MUX_s_1_2_2(mux_30_nl, or_tmp_43, ProductSum_for_asn_64_itm_3);
  assign or_1593_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7
      | (~ or_tmp_745);
  assign mux_538_nl = MUX_s_1_2_2(mux_537_cse, or_1593_nl, while_stage_0_9);
  assign or_1612_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7
      | (~ or_tmp_762);
  assign mux_546_nl = MUX_s_1_2_2(mux_545_cse, or_1612_nl, while_stage_0_9);
  assign or_1632_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_7
      | (~ or_tmp_779);
  assign mux_554_nl = MUX_s_1_2_2(mux_553_cse, or_1632_nl, while_stage_0_9);
  assign accum_vector_operator_1_for_not_13_nl = ~ accum_vector_operator_1_for_asn_25_itm_6;
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_131_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_117_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[2]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_124_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_96_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_110_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_132_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_133_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_135_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_banks_load_store_for_else_mux1h_11_nl = MUX1HOT_s_1_3_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[63]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[39]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[39]),
      {and_dcpl_580 , and_dcpl_582 , and_dcpl_584});
  assign weight_mem_banks_load_store_for_else_mux1h_38_nl = MUX1HOT_v_7_4_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[62:56]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[38:32]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[38:32]),
      rva_out_reg_data_46_40_sva_dfm_1_4, {and_dcpl_580 , and_dcpl_582 , and_dcpl_584
      , (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2)});
  assign not_2441_nl = ~ or_dcpl_679;
  assign weight_mem_banks_load_store_for_else_mux1h_18_nl = MUX1HOT_v_4_3_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[47:44]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[31:28]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[31:28]),
      {and_dcpl_580 , and_dcpl_582 , and_dcpl_584});
  assign not_2442_nl = ~ or_dcpl_679;
  assign weight_mem_banks_load_store_for_else_mux1h_39_nl = MUX1HOT_v_4_4_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[43:40]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[27:24]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[27:24]),
      rva_out_reg_data_35_32_sva_dfm_1_4, {and_dcpl_580 , and_dcpl_582 , and_dcpl_584
      , (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2)});
  assign not_2443_nl = ~ or_dcpl_679;
  assign and_918_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1])
      & (~ or_1401_tmp);
  assign and_919_nl = nor_464_cse & (~ or_1401_tmp);
  assign and_612_nl = (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1:0]==2'b01)
      & (~ or_1401_tmp);
  assign mux1h_2_nl = MUX1HOT_v_8_3_2((weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[63:56]),
      (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[63:56]), (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[15:8]),
      {and_918_nl , and_919_nl , and_612_nl});
  assign not_2450_nl = ~ or_1401_tmp;
  assign mux_109_nl = MUX_s_1_2_2((crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2]),
      (~ (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2])), crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1]);
  assign nor_350_nl = ~((crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2:1]!=2'b00));
  assign mux_110_nl = MUX_s_1_2_2(mux_109_nl, nor_350_nl, crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0]);
  assign and_613_nl = while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1]);
  assign and_615_nl = and_dcpl_588 & (~ (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0]));
  assign and_619_nl = and_dcpl_592 & (~(weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      | while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4));
  assign and_623_nl = weight_mem_read_arbxbar_xbar_1_for_3_4_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      & (~ weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1)
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign and_624_nl = weight_mem_read_arbxbar_xbar_1_for_3_6_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1
      & (~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4);
  assign weight_mem_banks_load_store_for_else_mux1h_20_nl = MUX1HOT_v_8_5_2((weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[47:40]),
      (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[47:40]), (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[7:0]),
      (weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d[7:0]), (weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d[7:0]),
      {and_613_nl , and_615_nl , and_619_nl , and_623_nl , and_624_nl});
  assign and_616_nl = and_dcpl_588 & (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0]);
  assign weight_mem_banks_load_store_for_else_or_nl = MUX_v_8_2_2(weight_mem_banks_load_store_for_else_mux1h_20_nl,
      8'b11111111, and_616_nl);
  assign or_1404_nl = ((~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[1])) & (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0])
      & and_dcpl_588) | ((~ while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4)
      & and_dcpl_592 & weight_mem_read_arbxbar_xbar_1_for_3_2_weight_mem_read_arbxbar_xbar_1_for_3_if_1_operator_8_false_3_or_mdf_sva_1);
  assign mux_489_nl = MUX_v_8_2_2(weight_mem_banks_load_store_for_else_or_nl, (weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[7:0]),
      or_1404_nl);
  assign or_1402_nl = (~ (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0]))
      | (weight_mem_write_arbxbar_xbar_for_empty_sva_2[1]);
  assign mux_475_nl = MUX_s_1_2_2(nor_tmp, or_1402_nl, weight_mem_write_arbxbar_xbar_for_empty_sva_2[4]);
  assign nor_522_nl = ~((mux_475_nl & and_dcpl_588) | ((weight_mem_write_arbxbar_xbar_for_empty_sva_2[2])
      & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_4
      & (crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1])));
  assign mux_115_nl = MUX_s_1_2_2(or_tmp_215, (~ mux_tmp_108), crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2]);
  assign mux_114_nl = MUX_s_1_2_2((~ mux_tmp_108), or_tmp_215, crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[2]);
  assign mux_116_nl = MUX_s_1_2_2(mux_115_nl, mux_114_nl, crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[1]);
  assign mux_113_nl = MUX_s_1_2_2((~ mux_tmp_108), or_tmp_215, or_362_cse);
  assign mux_117_nl = MUX_s_1_2_2(mux_116_nl, mux_113_nl, crossbar_spec_PE_Weight_WordType_8U_8U_source_tmp_1_lpi_1_dfm_2[0]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_126_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_127_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[3]);
  assign weight_mem_banks_load_store_for_else_mux1h_25_nl = MUX1HOT_v_2_3_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[39:38]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[23:22]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[23:22]),
      {and_dcpl_580 , and_dcpl_582 , and_dcpl_584});
  assign not_2444_nl = ~ or_dcpl_679;
  assign weight_mem_banks_load_store_for_else_mux1h_40_nl = MUX1HOT_v_6_4_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[37:32]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[21:16]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[21:16]),
      rva_out_reg_data_30_25_sva_dfm_2, {and_dcpl_580 , and_dcpl_582 , and_dcpl_584
      , (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2)});
  assign not_2445_nl = ~ or_dcpl_679;
  assign weight_mem_banks_load_store_for_else_mux1h_30_nl = MUX1HOT_s_1_3_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[31]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[15]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[15]),
      {and_dcpl_580 , and_dcpl_582 , and_dcpl_584});
  assign weight_mem_banks_load_store_for_else_mux1h_41_nl = MUX1HOT_v_7_4_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[30:24]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[14:8]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[14:8]),
      rva_out_reg_data_23_17_sva_dfm_2, {and_dcpl_580 , and_dcpl_582 , and_dcpl_584
      , (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2)});
  assign not_2447_nl = ~ or_dcpl_679;
  assign weight_mem_banks_load_store_for_else_mux1h_35_nl = MUX1HOT_s_1_3_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[23]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[7]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[7]),
      {and_dcpl_580 , and_dcpl_582 , and_dcpl_584});
  assign weight_mem_banks_load_store_for_else_mux1h_42_nl = MUX1HOT_v_7_4_2((weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d[22:16]),
      (weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d[6:0]), (weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d[6:0]),
      rva_out_reg_data_15_9_sva_dfm_4, {and_dcpl_580 , and_dcpl_582 , and_dcpl_584
      , (~ crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_2)});
  assign not_2449_nl = ~ or_dcpl_679;
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_113_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_72_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[5]);
  assign weight_mem_write_arbxbar_xbar_for_1_for_not_129_nl = ~ (weight_mem_write_arbxbar_xbar_for_empty_sva_2[0]);
  assign weight_mem_banks_load_store_for_else_weight_mem_banks_load_store_for_else_and_1_nl
      = MUX_v_8_2_2(8'b00000000, (weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d[15:8]),
      weight_mem_write_arbxbar_xbar_for_1_for_not_129_nl);
  assign mux_122_nl = MUX_s_1_2_2(weight_mem_run_3_for_land_1_lpi_1_dfm_1, (~ pe_manager_base_weight_slc_pe_manager_base_weight_2_0_178_itm_1),
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign input_mem_banks_read_1_for_mux_4_nl = MUX_v_64_256_2(input_mem_banks_bank_a_0_sva_dfm_2,
      input_mem_banks_bank_a_1_sva_dfm_2, input_mem_banks_bank_a_2_sva_dfm_2, input_mem_banks_bank_a_3_sva_dfm_2,
      input_mem_banks_bank_a_4_sva_dfm_2, input_mem_banks_bank_a_5_sva_dfm_2, input_mem_banks_bank_a_6_sva_dfm_2,
      input_mem_banks_bank_a_7_sva_dfm_2, input_mem_banks_bank_a_8_sva_dfm_2, input_mem_banks_bank_a_9_sva_dfm_2,
      input_mem_banks_bank_a_10_sva_dfm_2, input_mem_banks_bank_a_11_sva_dfm_2, input_mem_banks_bank_a_12_sva_dfm_2,
      input_mem_banks_bank_a_13_sva_dfm_2, input_mem_banks_bank_a_14_sva_dfm_2, input_mem_banks_bank_a_15_sva_dfm_2,
      input_mem_banks_bank_a_16_sva_dfm_2, input_mem_banks_bank_a_17_sva_dfm_2, input_mem_banks_bank_a_18_sva_dfm_2,
      input_mem_banks_bank_a_19_sva_dfm_2, input_mem_banks_bank_a_20_sva_dfm_2, input_mem_banks_bank_a_21_sva_dfm_2,
      input_mem_banks_bank_a_22_sva_dfm_2, input_mem_banks_bank_a_23_sva_dfm_2, input_mem_banks_bank_a_24_sva_dfm_2,
      input_mem_banks_bank_a_25_sva_dfm_2, input_mem_banks_bank_a_26_sva_dfm_2, input_mem_banks_bank_a_27_sva_dfm_2,
      input_mem_banks_bank_a_28_sva_dfm_2, input_mem_banks_bank_a_29_sva_dfm_2, input_mem_banks_bank_a_30_sva_dfm_2,
      input_mem_banks_bank_a_31_sva_dfm_2, input_mem_banks_bank_a_32_sva_dfm_2, input_mem_banks_bank_a_33_sva_dfm_2,
      input_mem_banks_bank_a_34_sva_dfm_2, input_mem_banks_bank_a_35_sva_dfm_2, input_mem_banks_bank_a_36_sva_dfm_2,
      input_mem_banks_bank_a_37_sva_dfm_2, input_mem_banks_bank_a_38_sva_dfm_2, input_mem_banks_bank_a_39_sva_dfm_2,
      input_mem_banks_bank_a_40_sva_dfm_2, input_mem_banks_bank_a_41_sva_dfm_2, input_mem_banks_bank_a_42_sva_dfm_2,
      input_mem_banks_bank_a_43_sva_dfm_2, input_mem_banks_bank_a_44_sva_dfm_2, input_mem_banks_bank_a_45_sva_dfm_2,
      input_mem_banks_bank_a_46_sva_dfm_2, input_mem_banks_bank_a_47_sva_dfm_2, input_mem_banks_bank_a_48_sva_dfm_2,
      input_mem_banks_bank_a_49_sva_dfm_2, input_mem_banks_bank_a_50_sva_dfm_2, input_mem_banks_bank_a_51_sva_dfm_2,
      input_mem_banks_bank_a_52_sva_dfm_2, input_mem_banks_bank_a_53_sva_dfm_2, input_mem_banks_bank_a_54_sva_dfm_2,
      input_mem_banks_bank_a_55_sva_dfm_2, input_mem_banks_bank_a_56_sva_dfm_2, input_mem_banks_bank_a_57_sva_dfm_2,
      input_mem_banks_bank_a_58_sva_dfm_2, input_mem_banks_bank_a_59_sva_dfm_2, input_mem_banks_bank_a_60_sva_dfm_2,
      input_mem_banks_bank_a_61_sva_dfm_2, input_mem_banks_bank_a_62_sva_dfm_2, input_mem_banks_bank_a_63_sva_dfm_2,
      input_mem_banks_bank_a_64_sva_dfm_2, input_mem_banks_bank_a_65_sva_dfm_2, input_mem_banks_bank_a_66_sva_dfm_2,
      input_mem_banks_bank_a_67_sva_dfm_2, input_mem_banks_bank_a_68_sva_dfm_2, input_mem_banks_bank_a_69_sva_dfm_2,
      input_mem_banks_bank_a_70_sva_dfm_2, input_mem_banks_bank_a_71_sva_dfm_2, input_mem_banks_bank_a_72_sva_dfm_2,
      input_mem_banks_bank_a_73_sva_dfm_2, input_mem_banks_bank_a_74_sva_dfm_2, input_mem_banks_bank_a_75_sva_dfm_2,
      input_mem_banks_bank_a_76_sva_dfm_2, input_mem_banks_bank_a_77_sva_dfm_2, input_mem_banks_bank_a_78_sva_dfm_2,
      input_mem_banks_bank_a_79_sva_dfm_2, input_mem_banks_bank_a_80_sva_dfm_2, input_mem_banks_bank_a_81_sva_dfm_2,
      input_mem_banks_bank_a_82_sva_dfm_2, input_mem_banks_bank_a_83_sva_dfm_2, input_mem_banks_bank_a_84_sva_dfm_2,
      input_mem_banks_bank_a_85_sva_dfm_2, input_mem_banks_bank_a_86_sva_dfm_2, input_mem_banks_bank_a_87_sva_dfm_2,
      input_mem_banks_bank_a_88_sva_dfm_2, input_mem_banks_bank_a_89_sva_dfm_2, input_mem_banks_bank_a_90_sva_dfm_2,
      input_mem_banks_bank_a_91_sva_dfm_2, input_mem_banks_bank_a_92_sva_dfm_2, input_mem_banks_bank_a_93_sva_dfm_2,
      input_mem_banks_bank_a_94_sva_dfm_2, input_mem_banks_bank_a_95_sva_dfm_2, input_mem_banks_bank_a_96_sva_dfm_2,
      input_mem_banks_bank_a_97_sva_dfm_2, input_mem_banks_bank_a_98_sva_dfm_2, input_mem_banks_bank_a_99_sva_dfm_2,
      input_mem_banks_bank_a_100_sva_dfm_2, input_mem_banks_bank_a_101_sva_dfm_2,
      input_mem_banks_bank_a_102_sva_dfm_2, input_mem_banks_bank_a_103_sva_dfm_2,
      input_mem_banks_bank_a_104_sva_dfm_2, input_mem_banks_bank_a_105_sva_dfm_2,
      input_mem_banks_bank_a_106_sva_dfm_2, input_mem_banks_bank_a_107_sva_dfm_2,
      input_mem_banks_bank_a_108_sva_dfm_2, input_mem_banks_bank_a_109_sva_dfm_2,
      input_mem_banks_bank_a_110_sva_dfm_2, input_mem_banks_bank_a_111_sva_dfm_2,
      input_mem_banks_bank_a_112_sva_dfm_2, input_mem_banks_bank_a_113_sva_dfm_2,
      input_mem_banks_bank_a_114_sva_dfm_2, input_mem_banks_bank_a_115_sva_dfm_2,
      input_mem_banks_bank_a_116_sva_dfm_2, input_mem_banks_bank_a_117_sva_dfm_2,
      input_mem_banks_bank_a_118_sva_dfm_2, input_mem_banks_bank_a_119_sva_dfm_2,
      input_mem_banks_bank_a_120_sva_dfm_2, input_mem_banks_bank_a_121_sva_dfm_2,
      input_mem_banks_bank_a_122_sva_dfm_2, input_mem_banks_bank_a_123_sva_dfm_2,
      input_mem_banks_bank_a_124_sva_dfm_2, input_mem_banks_bank_a_125_sva_dfm_2,
      input_mem_banks_bank_a_126_sva_dfm_2, input_mem_banks_bank_a_127_sva_dfm_2,
      input_mem_banks_bank_a_128_sva_dfm_2, input_mem_banks_bank_a_129_sva_dfm_2,
      input_mem_banks_bank_a_130_sva_dfm_2, input_mem_banks_bank_a_131_sva_dfm_2,
      input_mem_banks_bank_a_132_sva_dfm_2, input_mem_banks_bank_a_133_sva_dfm_2,
      input_mem_banks_bank_a_134_sva_dfm_2, input_mem_banks_bank_a_135_sva_dfm_2,
      input_mem_banks_bank_a_136_sva_dfm_2, input_mem_banks_bank_a_137_sva_dfm_2,
      input_mem_banks_bank_a_138_sva_dfm_2, input_mem_banks_bank_a_139_sva_dfm_2,
      input_mem_banks_bank_a_140_sva_dfm_2, input_mem_banks_bank_a_141_sva_dfm_2,
      input_mem_banks_bank_a_142_sva_dfm_2, input_mem_banks_bank_a_143_sva_dfm_2,
      input_mem_banks_bank_a_144_sva_dfm_2, input_mem_banks_bank_a_145_sva_dfm_2,
      input_mem_banks_bank_a_146_sva_dfm_2, input_mem_banks_bank_a_147_sva_dfm_2,
      input_mem_banks_bank_a_148_sva_dfm_2, input_mem_banks_bank_a_149_sva_dfm_2,
      input_mem_banks_bank_a_150_sva_dfm_2, input_mem_banks_bank_a_151_sva_dfm_2,
      input_mem_banks_bank_a_152_sva_dfm_2, input_mem_banks_bank_a_153_sva_dfm_2,
      input_mem_banks_bank_a_154_sva_dfm_2, input_mem_banks_bank_a_155_sva_dfm_2,
      input_mem_banks_bank_a_156_sva_dfm_2, input_mem_banks_bank_a_157_sva_dfm_2,
      input_mem_banks_bank_a_158_sva_dfm_2, input_mem_banks_bank_a_159_sva_dfm_2,
      input_mem_banks_bank_a_160_sva_dfm_2, input_mem_banks_bank_a_161_sva_dfm_2,
      input_mem_banks_bank_a_162_sva_dfm_2, input_mem_banks_bank_a_163_sva_dfm_2,
      input_mem_banks_bank_a_164_sva_dfm_2, input_mem_banks_bank_a_165_sva_dfm_2,
      input_mem_banks_bank_a_166_sva_dfm_2, input_mem_banks_bank_a_167_sva_dfm_2,
      input_mem_banks_bank_a_168_sva_dfm_2, input_mem_banks_bank_a_169_sva_dfm_2,
      input_mem_banks_bank_a_170_sva_dfm_2, input_mem_banks_bank_a_171_sva_dfm_2,
      input_mem_banks_bank_a_172_sva_dfm_2, input_mem_banks_bank_a_173_sva_dfm_2,
      input_mem_banks_bank_a_174_sva_dfm_2, input_mem_banks_bank_a_175_sva_dfm_2,
      input_mem_banks_bank_a_176_sva_dfm_2, input_mem_banks_bank_a_177_sva_dfm_2,
      input_mem_banks_bank_a_178_sva_dfm_2, input_mem_banks_bank_a_179_sva_dfm_2,
      input_mem_banks_bank_a_180_sva_dfm_2, input_mem_banks_bank_a_181_sva_dfm_2,
      input_mem_banks_bank_a_182_sva_dfm_2, input_mem_banks_bank_a_183_sva_dfm_2,
      input_mem_banks_bank_a_184_sva_dfm_2, input_mem_banks_bank_a_185_sva_dfm_2,
      input_mem_banks_bank_a_186_sva_dfm_2, input_mem_banks_bank_a_187_sva_dfm_2,
      input_mem_banks_bank_a_188_sva_dfm_2, input_mem_banks_bank_a_189_sva_dfm_2,
      input_mem_banks_bank_a_190_sva_dfm_2, input_mem_banks_bank_a_191_sva_dfm_2,
      input_mem_banks_bank_a_192_sva_dfm_2, input_mem_banks_bank_a_193_sva_dfm_2,
      input_mem_banks_bank_a_194_sva_dfm_2, input_mem_banks_bank_a_195_sva_dfm_2,
      input_mem_banks_bank_a_196_sva_dfm_2, input_mem_banks_bank_a_197_sva_dfm_2,
      input_mem_banks_bank_a_198_sva_dfm_2, input_mem_banks_bank_a_199_sva_dfm_2,
      input_mem_banks_bank_a_200_sva_dfm_2, input_mem_banks_bank_a_201_sva_dfm_2,
      input_mem_banks_bank_a_202_sva_dfm_2, input_mem_banks_bank_a_203_sva_dfm_2,
      input_mem_banks_bank_a_204_sva_dfm_2, input_mem_banks_bank_a_205_sva_dfm_2,
      input_mem_banks_bank_a_206_sva_dfm_2, input_mem_banks_bank_a_207_sva_dfm_2,
      input_mem_banks_bank_a_208_sva_dfm_2, input_mem_banks_bank_a_209_sva_dfm_2,
      input_mem_banks_bank_a_210_sva_dfm_2, input_mem_banks_bank_a_211_sva_dfm_2,
      input_mem_banks_bank_a_212_sva_dfm_2, input_mem_banks_bank_a_213_sva_dfm_2,
      input_mem_banks_bank_a_214_sva_dfm_2, input_mem_banks_bank_a_215_sva_dfm_2,
      input_mem_banks_bank_a_216_sva_dfm_2, input_mem_banks_bank_a_217_sva_dfm_2,
      input_mem_banks_bank_a_218_sva_dfm_2, input_mem_banks_bank_a_219_sva_dfm_2,
      input_mem_banks_bank_a_220_sva_dfm_2, input_mem_banks_bank_a_221_sva_dfm_2,
      input_mem_banks_bank_a_222_sva_dfm_2, input_mem_banks_bank_a_223_sva_dfm_2,
      input_mem_banks_bank_a_224_sva_dfm_2, input_mem_banks_bank_a_225_sva_dfm_2,
      input_mem_banks_bank_a_226_sva_dfm_2, input_mem_banks_bank_a_227_sva_dfm_2,
      input_mem_banks_bank_a_228_sva_dfm_2, input_mem_banks_bank_a_229_sva_dfm_2,
      input_mem_banks_bank_a_230_sva_dfm_2, input_mem_banks_bank_a_231_sva_dfm_2,
      input_mem_banks_bank_a_232_sva_dfm_2, input_mem_banks_bank_a_233_sva_dfm_2,
      input_mem_banks_bank_a_234_sva_dfm_2, input_mem_banks_bank_a_235_sva_dfm_2,
      input_mem_banks_bank_a_236_sva_dfm_2, input_mem_banks_bank_a_237_sva_dfm_2,
      input_mem_banks_bank_a_238_sva_dfm_2, input_mem_banks_bank_a_239_sva_dfm_2,
      input_mem_banks_bank_a_240_sva_dfm_2, input_mem_banks_bank_a_241_sva_dfm_2,
      input_mem_banks_bank_a_242_sva_dfm_2, input_mem_banks_bank_a_243_sva_dfm_2,
      input_mem_banks_bank_a_244_sva_dfm_2, input_mem_banks_bank_a_245_sva_dfm_2,
      input_mem_banks_bank_a_246_sva_dfm_2, input_mem_banks_bank_a_247_sva_dfm_2,
      input_mem_banks_bank_a_248_sva_dfm_2, input_mem_banks_bank_a_249_sva_dfm_2,
      input_mem_banks_bank_a_250_sva_dfm_2, input_mem_banks_bank_a_251_sva_dfm_2,
      input_mem_banks_bank_a_252_sva_dfm_2, input_mem_banks_bank_a_253_sva_dfm_2,
      input_mem_banks_bank_a_254_sva_dfm_2, input_mem_banks_bank_a_255_sva_dfm_2,
      input_read_addrs_sva_1_1);
  assign and_629_nl = (~ input_write_req_valid_lpi_1_dfm_1_1) & while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_1;
  assign weight_port_read_out_data_mux_20_nl = MUX_s_1_2_2(PECore_PushAxiRsp_if_else_mux_13_mx0w2,
      weight_port_read_out_data_0_7_sva_dfm_3_7, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign while_if_while_if_and_2_nl = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[14:0])
      & ({{14{PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0}}, PECore_DecodeAxiRead_switch_lp_equal_tmp_2_mx0w0})
      & ({{14{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt});
  assign or_1096_nl = or_dcpl_91 | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[16]) |
      (~ rva_in_PopNB_mioi_return_rsc_z_mxwt) | or_dcpl_658;
  assign mux_177_nl = MUX_s_1_2_2(PECore_RunMac_PECore_RunMac_if_and_svs_st_2, (weight_mem_write_arbxbar_xbar_for_lshift_tmp[3]),
      while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_2);
  assign and_699_nl = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_7_1 & Arbiter_8U_Roundrobin_pick_return_1_7_1_lpi_1_dfm_1_1
      & PECore_RunFSM_switch_lp_equal_tmp_1_2;
  assign mux_178_nl = MUX_s_1_2_2(and_699_nl, PECore_RunFSM_switch_lp_equal_tmp_1_2,
      and_700_cse);
  assign or_921_nl = Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_76_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_52_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_88_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_64_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_112_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_100_tmp;
  assign mux_179_nl = MUX_s_1_2_2(mux_178_nl, PECore_RunFSM_switch_lp_equal_tmp_1_2,
      or_921_nl);
  assign mux_180_nl = MUX_s_1_2_2(mux_179_nl, (~ or_tmp_334), while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign and_701_nl = Arbiter_8U_Roundrobin_pick_1_unequal_tmp_6_1 & reg_Arbiter_8U_Roundrobin_pick_return_1_7_1_7_lpi_1_dfm_1_5_cse
      & PECore_RunFSM_switch_lp_equal_tmp_1_2;
  assign mux_181_nl = MUX_s_1_2_2(and_701_nl, PECore_RunFSM_switch_lp_equal_tmp_1_2,
      and_702_cse);
  assign mux_182_nl = MUX_s_1_2_2(mux_181_nl, PECore_RunFSM_switch_lp_equal_tmp_1_2,
      and_703_cse);
  assign or_923_nl = Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_89_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_53_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_65_tmp
      | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_77_tmp | Arbiter_8U_Roundrobin_pick_1_Arbiter_8U_Roundrobin_pick_1_and_101_tmp;
  assign mux_183_nl = MUX_s_1_2_2(mux_182_nl, PECore_RunFSM_switch_lp_equal_tmp_1_2,
      or_923_nl);
  assign nor_354_nl = ~((~ PECore_DecodeAxiRead_switch_lp_equal_tmp_1_2) | rva_in_reg_rw_sva_3
      | input_read_req_valid_lpi_1_dfm_1_3 | crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_1
      | pe_manager_base_weight_slc_pe_manager_base_weight_2_0_178_itm_1);
  assign mux_184_nl = MUX_s_1_2_2(mux_183_nl, nor_354_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_3);
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_nl = pe_manager_base_weight_slc_pe_manager_base_weight_2_0_95_itm_1
      & (pe_manager_base_weight_sva[0]) & crossbar_spec_PE_Weight_WordType_8U_8U_1_for_not_1_itm_1
      & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_16_nl = pe_manager_base_weight_slc_pe_manager_base_weight_2_0_122_itm_1
      & (pe_manager_base_weight_sva[0]) & (~ (pe_manager_base_weight_sva[2])) & weight_mem_run_3_for_land_1_lpi_1_dfm_1;
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux_2_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_case_4_switch_lp_asn_2_itm_2,
      (pe_manager_base_weight_sva_mx1_3_0[0]), PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_2);
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux_3_nl = MUX_s_1_2_2(PECore_DecodeAxiRead_case_4_switch_lp_asn_1_itm_2,
      (pe_manager_base_weight_sva_mx2[8]), PECore_DecodeAxiRead_case_4_switch_lp_equal_tmp_1_2);
  assign PECore_DecodeAxiRead_switch_lp_PECore_DecodeAxiRead_switch_lp_and_1_nl =
      (while_if_slc_while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_23_4_3_itm_1[2])
      & PECore_DecodeAxiRead_switch_lp_nor_2_cse;
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux_7_nl = MUX_s_1_2_2(pe_config_is_valid_sva,
      pe_manager_zero_active_sva, and_321_cse);
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux_8_nl = MUX_s_1_2_2(pe_config_is_zero_first_sva_mx1,
      (pe_manager_num_input_sva[0]), and_321_cse);
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux_9_nl = MUX_v_4_2_2(pe_config_num_manager_sva,
      (pe_manager_base_bias_sva[3:0]), and_321_cse);
  assign PECore_DecodeAxiRead_case_4_switch_lp_mux_10_nl = MUX_v_7_2_2((pe_config_num_output_sva[6:0]),
      (pe_manager_base_bias_sva[14:8]), and_321_cse);
  assign and_2582_nl = (reg_weight_mem_run_3_for_5_and_168_itm_2_cse | reg_weight_mem_run_3_for_5_and_167_itm_2_cse
      | reg_weight_mem_run_3_for_5_and_166_itm_2_cse | reg_weight_mem_run_3_for_5_and_165_itm_2_cse
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_56_itm_2 | reg_weight_mem_run_3_for_5_and_163_itm_2_cse
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_54_itm_2 | reg_weight_mem_run_3_for_5_weight_mem_run_3_for_5_nor_20_itm_2_cse)
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign mux_1256_nl = MUX_s_1_2_2(and_2582_nl, or_3653_cse, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign or_3662_nl = reg_weight_mem_run_3_for_5_and_168_itm_2_cse | reg_weight_mem_run_3_for_5_and_167_itm_2_cse
      | reg_weight_mem_run_3_for_5_and_166_itm_2_cse | reg_weight_mem_run_3_for_5_and_165_itm_2_cse
      | weight_mem_run_3_for_5_and_164_itm_2 | reg_weight_mem_run_3_for_5_and_163_itm_2_cse
      | weight_mem_run_3_for_5_and_162_itm_2 | weight_mem_run_3_for_5_and_161_cse;
  assign mux_1257_nl = MUX_s_1_2_2(or_3659_cse, or_3658_cse, reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[2]);
  assign mux_1258_nl = MUX_s_1_2_2(mux_1257_nl, or_3657_cse, reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[0]);
  assign or_3660_nl = or_tmp_2762 | (crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3
      & mux_1258_nl);
  assign mux_1259_nl = MUX_s_1_2_2(or_3662_nl, or_3660_nl, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign and_2584_nl = (reg_weight_mem_run_3_for_5_and_168_itm_2_cse | reg_weight_mem_run_3_for_5_and_167_itm_2_cse
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_10_itm_2 | reg_weight_mem_run_3_for_5_and_165_itm_2_cse
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_56_itm_2 | reg_weight_mem_run_3_for_5_and_163_itm_2_cse
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_and_54_itm_2 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_crossbar_spec_PE_Weight_WordType_8U_8U_1_for_nor_itm_3)
      & weight_mem_run_3_for_land_1_lpi_1_dfm_3;
  assign mux_1262_nl = MUX_s_1_2_2(and_2584_nl, or_3653_cse, while_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_st_5);
  assign mux_1279_nl = MUX_s_1_2_2(not_tmp_1925, or_tmp_2778, or_3659_cse);
  assign mux_1278_nl = MUX_s_1_2_2(not_tmp_1925, or_tmp_2778, or_3658_cse);
  assign mux_1280_nl = MUX_s_1_2_2(mux_1279_nl, mux_1278_nl, reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[2]);
  assign mux_1277_nl = MUX_s_1_2_2(not_tmp_1925, or_tmp_2778, or_3657_cse);
  assign mux_1281_nl = MUX_s_1_2_2(mux_1280_nl, mux_1277_nl, reg_weight_read_addrs_1_lpi_1_dfm_3_2_0_cse[0]);
  assign mux_1282_nl = MUX_s_1_2_2(not_tmp_1925, mux_1281_nl, crossbar_spec_PE_Weight_WordType_8U_8U_for_land_1_lpi_1_dfm_3);
  assign or_3684_nl = crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_62_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_71_itm_1 | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_72_itm_1
      | crossbar_spec_PE_Weight_WordType_8U_8U_1_for_if_1_and_47_itm_1;
  assign mux_1283_nl = MUX_s_1_2_2(mux_1282_nl, or_tmp_2778, or_3684_nl);
  assign mux_1290_nl = MUX_s_1_2_2(mux_1268_cse, or_tmp_2778, or_tmp_2755);
  assign mux_1297_nl = MUX_s_1_2_2(mux_1268_cse, or_tmp_2778, or_tmp_2762);

  function automatic  MUX1HOT_s_1_1_2;
    input  input_0;
    input  sel;
    reg  result;
  begin
    result = input_0 & sel;
    MUX1HOT_s_1_1_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_3_2;
    input  input_2;
    input  input_1;
    input  input_0;
    input [2:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_4_2;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [3:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_7_2;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [6:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    MUX1HOT_s_1_7_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_8_2;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [7:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    MUX1HOT_s_1_8_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_9_2;
    input  input_8;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [8:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    MUX1HOT_s_1_9_2 = result;
  end
  endfunction


  function automatic [10:0] MUX1HOT_v_11_8_2;
    input [10:0] input_7;
    input [10:0] input_6;
    input [10:0] input_5;
    input [10:0] input_4;
    input [10:0] input_3;
    input [10:0] input_2;
    input [10:0] input_1;
    input [10:0] input_0;
    input [7:0] sel;
    reg [10:0] result;
  begin
    result = input_0 & {11{sel[0]}};
    result = result | (input_1 & {11{sel[1]}});
    result = result | (input_2 & {11{sel[2]}});
    result = result | (input_3 & {11{sel[3]}});
    result = result | (input_4 & {11{sel[4]}});
    result = result | (input_5 & {11{sel[5]}});
    result = result | (input_6 & {11{sel[6]}});
    result = result | (input_7 & {11{sel[7]}});
    MUX1HOT_v_11_8_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_3_2;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [2:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    MUX1HOT_v_2_3_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_4_2;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [3:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    result = result | (input_3 & {2{sel[3]}});
    MUX1HOT_v_2_4_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_3_2;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [2:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | (input_1 & {3{sel[1]}});
    result = result | (input_2 & {3{sel[2]}});
    MUX1HOT_v_3_3_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_4_2;
    input [2:0] input_3;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [3:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | (input_1 & {3{sel[1]}});
    result = result | (input_2 & {3{sel[2]}});
    result = result | (input_3 & {3{sel[3]}});
    MUX1HOT_v_3_4_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_8_2;
    input [2:0] input_7;
    input [2:0] input_6;
    input [2:0] input_5;
    input [2:0] input_4;
    input [2:0] input_3;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [7:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | (input_1 & {3{sel[1]}});
    result = result | (input_2 & {3{sel[2]}});
    result = result | (input_3 & {3{sel[3]}});
    result = result | (input_4 & {3{sel[4]}});
    result = result | (input_5 & {3{sel[5]}});
    result = result | (input_6 & {3{sel[6]}});
    result = result | (input_7 & {3{sel[7]}});
    MUX1HOT_v_3_8_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_3_2;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [2:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    MUX1HOT_v_4_3_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_4_2;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [3:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    MUX1HOT_v_4_4_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_8_2;
    input [3:0] input_7;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [7:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    result = result | (input_5 & {4{sel[5]}});
    result = result | (input_6 & {4{sel[6]}});
    result = result | (input_7 & {4{sel[7]}});
    MUX1HOT_v_4_8_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_4_2;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [3:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    result = result | (input_3 & {5{sel[3]}});
    MUX1HOT_v_5_4_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_3_2;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [2:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | (input_1 & {64{sel[1]}});
    result = result | (input_2 & {64{sel[2]}});
    MUX1HOT_v_64_3_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_3_2;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [2:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | (input_1 & {6{sel[1]}});
    result = result | (input_2 & {6{sel[2]}});
    MUX1HOT_v_6_3_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_4_2;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [3:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | (input_1 & {6{sel[1]}});
    result = result | (input_2 & {6{sel[2]}});
    result = result | (input_3 & {6{sel[3]}});
    MUX1HOT_v_6_4_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_8_2;
    input [5:0] input_7;
    input [5:0] input_6;
    input [5:0] input_5;
    input [5:0] input_4;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [7:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | (input_1 & {6{sel[1]}});
    result = result | (input_2 & {6{sel[2]}});
    result = result | (input_3 & {6{sel[3]}});
    result = result | (input_4 & {6{sel[4]}});
    result = result | (input_5 & {6{sel[5]}});
    result = result | (input_6 & {6{sel[6]}});
    result = result | (input_7 & {6{sel[7]}});
    MUX1HOT_v_6_8_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_3_2;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [2:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | (input_1 & {7{sel[1]}});
    result = result | (input_2 & {7{sel[2]}});
    MUX1HOT_v_7_3_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_4_2;
    input [6:0] input_3;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [3:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | (input_1 & {7{sel[1]}});
    result = result | (input_2 & {7{sel[2]}});
    result = result | (input_3 & {7{sel[3]}});
    MUX1HOT_v_7_4_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_8_2;
    input [6:0] input_7;
    input [6:0] input_6;
    input [6:0] input_5;
    input [6:0] input_4;
    input [6:0] input_3;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [7:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | (input_1 & {7{sel[1]}});
    result = result | (input_2 & {7{sel[2]}});
    result = result | (input_3 & {7{sel[3]}});
    result = result | (input_4 & {7{sel[4]}});
    result = result | (input_5 & {7{sel[5]}});
    result = result | (input_6 & {7{sel[6]}});
    result = result | (input_7 & {7{sel[7]}});
    MUX1HOT_v_7_8_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_9_2;
    input [6:0] input_8;
    input [6:0] input_7;
    input [6:0] input_6;
    input [6:0] input_5;
    input [6:0] input_4;
    input [6:0] input_3;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [8:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | (input_1 & {7{sel[1]}});
    result = result | (input_2 & {7{sel[2]}});
    result = result | (input_3 & {7{sel[3]}});
    result = result | (input_4 & {7{sel[4]}});
    result = result | (input_5 & {7{sel[5]}});
    result = result | (input_6 & {7{sel[6]}});
    result = result | (input_7 & {7{sel[7]}});
    result = result | (input_8 & {7{sel[8]}});
    MUX1HOT_v_7_9_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_3_2;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [2:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    MUX1HOT_v_8_3_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_5_2;
    input [7:0] input_4;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [4:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    result = result | (input_3 & {8{sel[3]}});
    result = result | (input_4 & {8{sel[4]}});
    MUX1HOT_v_8_5_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_6_2;
    input [7:0] input_5;
    input [7:0] input_4;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [5:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    result = result | (input_3 & {8{sel[3]}});
    result = result | (input_4 & {8{sel[4]}});
    result = result | (input_5 & {8{sel[5]}});
    MUX1HOT_v_8_6_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_8_2;
    input [7:0] input_7;
    input [7:0] input_6;
    input [7:0] input_5;
    input [7:0] input_4;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [7:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    result = result | (input_3 & {8{sel[3]}});
    result = result | (input_4 & {8{sel[4]}});
    result = result | (input_5 & {8{sel[5]}});
    result = result | (input_6 & {8{sel[6]}});
    result = result | (input_7 & {8{sel[7]}});
    MUX1HOT_v_8_8_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_9_2;
    input [7:0] input_8;
    input [7:0] input_7;
    input [7:0] input_6;
    input [7:0] input_5;
    input [7:0] input_4;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [8:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    result = result | (input_3 & {8{sel[3]}});
    result = result | (input_4 & {8{sel[4]}});
    result = result | (input_5 & {8{sel[5]}});
    result = result | (input_6 & {8{sel[6]}});
    result = result | (input_7 & {8{sel[7]}});
    result = result | (input_8 & {8{sel[8]}});
    MUX1HOT_v_8_9_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_8_2;
    input  input_0;
    input  input_1;
    input  input_2;
    input  input_3;
    input  input_4;
    input  input_5;
    input  input_6;
    input  input_7;
    input [2:0] sel;
    reg  result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_s_1_8_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_2_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input  sel;
    reg [10:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_11_2_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_8_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input [10:0] input_2;
    input [10:0] input_3;
    input [10:0] input_4;
    input [10:0] input_5;
    input [10:0] input_6;
    input [10:0] input_7;
    input [2:0] sel;
    reg [10:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_11_8_2 = result;
  end
  endfunction


  function automatic [12:0] MUX_v_13_2_2;
    input [12:0] input_0;
    input [12:0] input_1;
    input  sel;
    reg [12:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_13_2_2 = result;
  end
  endfunction


  function automatic [13:0] MUX_v_14_2_2;
    input [13:0] input_0;
    input [13:0] input_1;
    input  sel;
    reg [13:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_14_2_2 = result;
  end
  endfunction


  function automatic [14:0] MUX_v_15_2_2;
    input [14:0] input_0;
    input [14:0] input_1;
    input  sel;
    reg [14:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_15_2_2 = result;
  end
  endfunction


  function automatic [19:0] MUX_v_20_2_2;
    input [19:0] input_0;
    input [19:0] input_1;
    input  sel;
    reg [19:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_20_2_2 = result;
  end
  endfunction


  function automatic [22:0] MUX_v_23_2_2;
    input [22:0] input_0;
    input [22:0] input_1;
    input  sel;
    reg [22:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_23_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input  sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input  sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input  sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_8_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [3:0] input_2;
    input [3:0] input_3;
    input [3:0] input_4;
    input [3:0] input_5;
    input [3:0] input_6;
    input [3:0] input_7;
    input [2:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_4_8_2 = result;
  end
  endfunction


  function automatic [55:0] MUX_v_56_2_2;
    input [55:0] input_0;
    input [55:0] input_1;
    input  sel;
    reg [55:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_56_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input  sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_256_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [63:0] input_2;
    input [63:0] input_3;
    input [63:0] input_4;
    input [63:0] input_5;
    input [63:0] input_6;
    input [63:0] input_7;
    input [63:0] input_8;
    input [63:0] input_9;
    input [63:0] input_10;
    input [63:0] input_11;
    input [63:0] input_12;
    input [63:0] input_13;
    input [63:0] input_14;
    input [63:0] input_15;
    input [63:0] input_16;
    input [63:0] input_17;
    input [63:0] input_18;
    input [63:0] input_19;
    input [63:0] input_20;
    input [63:0] input_21;
    input [63:0] input_22;
    input [63:0] input_23;
    input [63:0] input_24;
    input [63:0] input_25;
    input [63:0] input_26;
    input [63:0] input_27;
    input [63:0] input_28;
    input [63:0] input_29;
    input [63:0] input_30;
    input [63:0] input_31;
    input [63:0] input_32;
    input [63:0] input_33;
    input [63:0] input_34;
    input [63:0] input_35;
    input [63:0] input_36;
    input [63:0] input_37;
    input [63:0] input_38;
    input [63:0] input_39;
    input [63:0] input_40;
    input [63:0] input_41;
    input [63:0] input_42;
    input [63:0] input_43;
    input [63:0] input_44;
    input [63:0] input_45;
    input [63:0] input_46;
    input [63:0] input_47;
    input [63:0] input_48;
    input [63:0] input_49;
    input [63:0] input_50;
    input [63:0] input_51;
    input [63:0] input_52;
    input [63:0] input_53;
    input [63:0] input_54;
    input [63:0] input_55;
    input [63:0] input_56;
    input [63:0] input_57;
    input [63:0] input_58;
    input [63:0] input_59;
    input [63:0] input_60;
    input [63:0] input_61;
    input [63:0] input_62;
    input [63:0] input_63;
    input [63:0] input_64;
    input [63:0] input_65;
    input [63:0] input_66;
    input [63:0] input_67;
    input [63:0] input_68;
    input [63:0] input_69;
    input [63:0] input_70;
    input [63:0] input_71;
    input [63:0] input_72;
    input [63:0] input_73;
    input [63:0] input_74;
    input [63:0] input_75;
    input [63:0] input_76;
    input [63:0] input_77;
    input [63:0] input_78;
    input [63:0] input_79;
    input [63:0] input_80;
    input [63:0] input_81;
    input [63:0] input_82;
    input [63:0] input_83;
    input [63:0] input_84;
    input [63:0] input_85;
    input [63:0] input_86;
    input [63:0] input_87;
    input [63:0] input_88;
    input [63:0] input_89;
    input [63:0] input_90;
    input [63:0] input_91;
    input [63:0] input_92;
    input [63:0] input_93;
    input [63:0] input_94;
    input [63:0] input_95;
    input [63:0] input_96;
    input [63:0] input_97;
    input [63:0] input_98;
    input [63:0] input_99;
    input [63:0] input_100;
    input [63:0] input_101;
    input [63:0] input_102;
    input [63:0] input_103;
    input [63:0] input_104;
    input [63:0] input_105;
    input [63:0] input_106;
    input [63:0] input_107;
    input [63:0] input_108;
    input [63:0] input_109;
    input [63:0] input_110;
    input [63:0] input_111;
    input [63:0] input_112;
    input [63:0] input_113;
    input [63:0] input_114;
    input [63:0] input_115;
    input [63:0] input_116;
    input [63:0] input_117;
    input [63:0] input_118;
    input [63:0] input_119;
    input [63:0] input_120;
    input [63:0] input_121;
    input [63:0] input_122;
    input [63:0] input_123;
    input [63:0] input_124;
    input [63:0] input_125;
    input [63:0] input_126;
    input [63:0] input_127;
    input [63:0] input_128;
    input [63:0] input_129;
    input [63:0] input_130;
    input [63:0] input_131;
    input [63:0] input_132;
    input [63:0] input_133;
    input [63:0] input_134;
    input [63:0] input_135;
    input [63:0] input_136;
    input [63:0] input_137;
    input [63:0] input_138;
    input [63:0] input_139;
    input [63:0] input_140;
    input [63:0] input_141;
    input [63:0] input_142;
    input [63:0] input_143;
    input [63:0] input_144;
    input [63:0] input_145;
    input [63:0] input_146;
    input [63:0] input_147;
    input [63:0] input_148;
    input [63:0] input_149;
    input [63:0] input_150;
    input [63:0] input_151;
    input [63:0] input_152;
    input [63:0] input_153;
    input [63:0] input_154;
    input [63:0] input_155;
    input [63:0] input_156;
    input [63:0] input_157;
    input [63:0] input_158;
    input [63:0] input_159;
    input [63:0] input_160;
    input [63:0] input_161;
    input [63:0] input_162;
    input [63:0] input_163;
    input [63:0] input_164;
    input [63:0] input_165;
    input [63:0] input_166;
    input [63:0] input_167;
    input [63:0] input_168;
    input [63:0] input_169;
    input [63:0] input_170;
    input [63:0] input_171;
    input [63:0] input_172;
    input [63:0] input_173;
    input [63:0] input_174;
    input [63:0] input_175;
    input [63:0] input_176;
    input [63:0] input_177;
    input [63:0] input_178;
    input [63:0] input_179;
    input [63:0] input_180;
    input [63:0] input_181;
    input [63:0] input_182;
    input [63:0] input_183;
    input [63:0] input_184;
    input [63:0] input_185;
    input [63:0] input_186;
    input [63:0] input_187;
    input [63:0] input_188;
    input [63:0] input_189;
    input [63:0] input_190;
    input [63:0] input_191;
    input [63:0] input_192;
    input [63:0] input_193;
    input [63:0] input_194;
    input [63:0] input_195;
    input [63:0] input_196;
    input [63:0] input_197;
    input [63:0] input_198;
    input [63:0] input_199;
    input [63:0] input_200;
    input [63:0] input_201;
    input [63:0] input_202;
    input [63:0] input_203;
    input [63:0] input_204;
    input [63:0] input_205;
    input [63:0] input_206;
    input [63:0] input_207;
    input [63:0] input_208;
    input [63:0] input_209;
    input [63:0] input_210;
    input [63:0] input_211;
    input [63:0] input_212;
    input [63:0] input_213;
    input [63:0] input_214;
    input [63:0] input_215;
    input [63:0] input_216;
    input [63:0] input_217;
    input [63:0] input_218;
    input [63:0] input_219;
    input [63:0] input_220;
    input [63:0] input_221;
    input [63:0] input_222;
    input [63:0] input_223;
    input [63:0] input_224;
    input [63:0] input_225;
    input [63:0] input_226;
    input [63:0] input_227;
    input [63:0] input_228;
    input [63:0] input_229;
    input [63:0] input_230;
    input [63:0] input_231;
    input [63:0] input_232;
    input [63:0] input_233;
    input [63:0] input_234;
    input [63:0] input_235;
    input [63:0] input_236;
    input [63:0] input_237;
    input [63:0] input_238;
    input [63:0] input_239;
    input [63:0] input_240;
    input [63:0] input_241;
    input [63:0] input_242;
    input [63:0] input_243;
    input [63:0] input_244;
    input [63:0] input_245;
    input [63:0] input_246;
    input [63:0] input_247;
    input [63:0] input_248;
    input [63:0] input_249;
    input [63:0] input_250;
    input [63:0] input_251;
    input [63:0] input_252;
    input [63:0] input_253;
    input [63:0] input_254;
    input [63:0] input_255;
    input [7:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      8'b00000000 : begin
        result = input_0;
      end
      8'b00000001 : begin
        result = input_1;
      end
      8'b00000010 : begin
        result = input_2;
      end
      8'b00000011 : begin
        result = input_3;
      end
      8'b00000100 : begin
        result = input_4;
      end
      8'b00000101 : begin
        result = input_5;
      end
      8'b00000110 : begin
        result = input_6;
      end
      8'b00000111 : begin
        result = input_7;
      end
      8'b00001000 : begin
        result = input_8;
      end
      8'b00001001 : begin
        result = input_9;
      end
      8'b00001010 : begin
        result = input_10;
      end
      8'b00001011 : begin
        result = input_11;
      end
      8'b00001100 : begin
        result = input_12;
      end
      8'b00001101 : begin
        result = input_13;
      end
      8'b00001110 : begin
        result = input_14;
      end
      8'b00001111 : begin
        result = input_15;
      end
      8'b00010000 : begin
        result = input_16;
      end
      8'b00010001 : begin
        result = input_17;
      end
      8'b00010010 : begin
        result = input_18;
      end
      8'b00010011 : begin
        result = input_19;
      end
      8'b00010100 : begin
        result = input_20;
      end
      8'b00010101 : begin
        result = input_21;
      end
      8'b00010110 : begin
        result = input_22;
      end
      8'b00010111 : begin
        result = input_23;
      end
      8'b00011000 : begin
        result = input_24;
      end
      8'b00011001 : begin
        result = input_25;
      end
      8'b00011010 : begin
        result = input_26;
      end
      8'b00011011 : begin
        result = input_27;
      end
      8'b00011100 : begin
        result = input_28;
      end
      8'b00011101 : begin
        result = input_29;
      end
      8'b00011110 : begin
        result = input_30;
      end
      8'b00011111 : begin
        result = input_31;
      end
      8'b00100000 : begin
        result = input_32;
      end
      8'b00100001 : begin
        result = input_33;
      end
      8'b00100010 : begin
        result = input_34;
      end
      8'b00100011 : begin
        result = input_35;
      end
      8'b00100100 : begin
        result = input_36;
      end
      8'b00100101 : begin
        result = input_37;
      end
      8'b00100110 : begin
        result = input_38;
      end
      8'b00100111 : begin
        result = input_39;
      end
      8'b00101000 : begin
        result = input_40;
      end
      8'b00101001 : begin
        result = input_41;
      end
      8'b00101010 : begin
        result = input_42;
      end
      8'b00101011 : begin
        result = input_43;
      end
      8'b00101100 : begin
        result = input_44;
      end
      8'b00101101 : begin
        result = input_45;
      end
      8'b00101110 : begin
        result = input_46;
      end
      8'b00101111 : begin
        result = input_47;
      end
      8'b00110000 : begin
        result = input_48;
      end
      8'b00110001 : begin
        result = input_49;
      end
      8'b00110010 : begin
        result = input_50;
      end
      8'b00110011 : begin
        result = input_51;
      end
      8'b00110100 : begin
        result = input_52;
      end
      8'b00110101 : begin
        result = input_53;
      end
      8'b00110110 : begin
        result = input_54;
      end
      8'b00110111 : begin
        result = input_55;
      end
      8'b00111000 : begin
        result = input_56;
      end
      8'b00111001 : begin
        result = input_57;
      end
      8'b00111010 : begin
        result = input_58;
      end
      8'b00111011 : begin
        result = input_59;
      end
      8'b00111100 : begin
        result = input_60;
      end
      8'b00111101 : begin
        result = input_61;
      end
      8'b00111110 : begin
        result = input_62;
      end
      8'b00111111 : begin
        result = input_63;
      end
      8'b01000000 : begin
        result = input_64;
      end
      8'b01000001 : begin
        result = input_65;
      end
      8'b01000010 : begin
        result = input_66;
      end
      8'b01000011 : begin
        result = input_67;
      end
      8'b01000100 : begin
        result = input_68;
      end
      8'b01000101 : begin
        result = input_69;
      end
      8'b01000110 : begin
        result = input_70;
      end
      8'b01000111 : begin
        result = input_71;
      end
      8'b01001000 : begin
        result = input_72;
      end
      8'b01001001 : begin
        result = input_73;
      end
      8'b01001010 : begin
        result = input_74;
      end
      8'b01001011 : begin
        result = input_75;
      end
      8'b01001100 : begin
        result = input_76;
      end
      8'b01001101 : begin
        result = input_77;
      end
      8'b01001110 : begin
        result = input_78;
      end
      8'b01001111 : begin
        result = input_79;
      end
      8'b01010000 : begin
        result = input_80;
      end
      8'b01010001 : begin
        result = input_81;
      end
      8'b01010010 : begin
        result = input_82;
      end
      8'b01010011 : begin
        result = input_83;
      end
      8'b01010100 : begin
        result = input_84;
      end
      8'b01010101 : begin
        result = input_85;
      end
      8'b01010110 : begin
        result = input_86;
      end
      8'b01010111 : begin
        result = input_87;
      end
      8'b01011000 : begin
        result = input_88;
      end
      8'b01011001 : begin
        result = input_89;
      end
      8'b01011010 : begin
        result = input_90;
      end
      8'b01011011 : begin
        result = input_91;
      end
      8'b01011100 : begin
        result = input_92;
      end
      8'b01011101 : begin
        result = input_93;
      end
      8'b01011110 : begin
        result = input_94;
      end
      8'b01011111 : begin
        result = input_95;
      end
      8'b01100000 : begin
        result = input_96;
      end
      8'b01100001 : begin
        result = input_97;
      end
      8'b01100010 : begin
        result = input_98;
      end
      8'b01100011 : begin
        result = input_99;
      end
      8'b01100100 : begin
        result = input_100;
      end
      8'b01100101 : begin
        result = input_101;
      end
      8'b01100110 : begin
        result = input_102;
      end
      8'b01100111 : begin
        result = input_103;
      end
      8'b01101000 : begin
        result = input_104;
      end
      8'b01101001 : begin
        result = input_105;
      end
      8'b01101010 : begin
        result = input_106;
      end
      8'b01101011 : begin
        result = input_107;
      end
      8'b01101100 : begin
        result = input_108;
      end
      8'b01101101 : begin
        result = input_109;
      end
      8'b01101110 : begin
        result = input_110;
      end
      8'b01101111 : begin
        result = input_111;
      end
      8'b01110000 : begin
        result = input_112;
      end
      8'b01110001 : begin
        result = input_113;
      end
      8'b01110010 : begin
        result = input_114;
      end
      8'b01110011 : begin
        result = input_115;
      end
      8'b01110100 : begin
        result = input_116;
      end
      8'b01110101 : begin
        result = input_117;
      end
      8'b01110110 : begin
        result = input_118;
      end
      8'b01110111 : begin
        result = input_119;
      end
      8'b01111000 : begin
        result = input_120;
      end
      8'b01111001 : begin
        result = input_121;
      end
      8'b01111010 : begin
        result = input_122;
      end
      8'b01111011 : begin
        result = input_123;
      end
      8'b01111100 : begin
        result = input_124;
      end
      8'b01111101 : begin
        result = input_125;
      end
      8'b01111110 : begin
        result = input_126;
      end
      8'b01111111 : begin
        result = input_127;
      end
      8'b10000000 : begin
        result = input_128;
      end
      8'b10000001 : begin
        result = input_129;
      end
      8'b10000010 : begin
        result = input_130;
      end
      8'b10000011 : begin
        result = input_131;
      end
      8'b10000100 : begin
        result = input_132;
      end
      8'b10000101 : begin
        result = input_133;
      end
      8'b10000110 : begin
        result = input_134;
      end
      8'b10000111 : begin
        result = input_135;
      end
      8'b10001000 : begin
        result = input_136;
      end
      8'b10001001 : begin
        result = input_137;
      end
      8'b10001010 : begin
        result = input_138;
      end
      8'b10001011 : begin
        result = input_139;
      end
      8'b10001100 : begin
        result = input_140;
      end
      8'b10001101 : begin
        result = input_141;
      end
      8'b10001110 : begin
        result = input_142;
      end
      8'b10001111 : begin
        result = input_143;
      end
      8'b10010000 : begin
        result = input_144;
      end
      8'b10010001 : begin
        result = input_145;
      end
      8'b10010010 : begin
        result = input_146;
      end
      8'b10010011 : begin
        result = input_147;
      end
      8'b10010100 : begin
        result = input_148;
      end
      8'b10010101 : begin
        result = input_149;
      end
      8'b10010110 : begin
        result = input_150;
      end
      8'b10010111 : begin
        result = input_151;
      end
      8'b10011000 : begin
        result = input_152;
      end
      8'b10011001 : begin
        result = input_153;
      end
      8'b10011010 : begin
        result = input_154;
      end
      8'b10011011 : begin
        result = input_155;
      end
      8'b10011100 : begin
        result = input_156;
      end
      8'b10011101 : begin
        result = input_157;
      end
      8'b10011110 : begin
        result = input_158;
      end
      8'b10011111 : begin
        result = input_159;
      end
      8'b10100000 : begin
        result = input_160;
      end
      8'b10100001 : begin
        result = input_161;
      end
      8'b10100010 : begin
        result = input_162;
      end
      8'b10100011 : begin
        result = input_163;
      end
      8'b10100100 : begin
        result = input_164;
      end
      8'b10100101 : begin
        result = input_165;
      end
      8'b10100110 : begin
        result = input_166;
      end
      8'b10100111 : begin
        result = input_167;
      end
      8'b10101000 : begin
        result = input_168;
      end
      8'b10101001 : begin
        result = input_169;
      end
      8'b10101010 : begin
        result = input_170;
      end
      8'b10101011 : begin
        result = input_171;
      end
      8'b10101100 : begin
        result = input_172;
      end
      8'b10101101 : begin
        result = input_173;
      end
      8'b10101110 : begin
        result = input_174;
      end
      8'b10101111 : begin
        result = input_175;
      end
      8'b10110000 : begin
        result = input_176;
      end
      8'b10110001 : begin
        result = input_177;
      end
      8'b10110010 : begin
        result = input_178;
      end
      8'b10110011 : begin
        result = input_179;
      end
      8'b10110100 : begin
        result = input_180;
      end
      8'b10110101 : begin
        result = input_181;
      end
      8'b10110110 : begin
        result = input_182;
      end
      8'b10110111 : begin
        result = input_183;
      end
      8'b10111000 : begin
        result = input_184;
      end
      8'b10111001 : begin
        result = input_185;
      end
      8'b10111010 : begin
        result = input_186;
      end
      8'b10111011 : begin
        result = input_187;
      end
      8'b10111100 : begin
        result = input_188;
      end
      8'b10111101 : begin
        result = input_189;
      end
      8'b10111110 : begin
        result = input_190;
      end
      8'b10111111 : begin
        result = input_191;
      end
      8'b11000000 : begin
        result = input_192;
      end
      8'b11000001 : begin
        result = input_193;
      end
      8'b11000010 : begin
        result = input_194;
      end
      8'b11000011 : begin
        result = input_195;
      end
      8'b11000100 : begin
        result = input_196;
      end
      8'b11000101 : begin
        result = input_197;
      end
      8'b11000110 : begin
        result = input_198;
      end
      8'b11000111 : begin
        result = input_199;
      end
      8'b11001000 : begin
        result = input_200;
      end
      8'b11001001 : begin
        result = input_201;
      end
      8'b11001010 : begin
        result = input_202;
      end
      8'b11001011 : begin
        result = input_203;
      end
      8'b11001100 : begin
        result = input_204;
      end
      8'b11001101 : begin
        result = input_205;
      end
      8'b11001110 : begin
        result = input_206;
      end
      8'b11001111 : begin
        result = input_207;
      end
      8'b11010000 : begin
        result = input_208;
      end
      8'b11010001 : begin
        result = input_209;
      end
      8'b11010010 : begin
        result = input_210;
      end
      8'b11010011 : begin
        result = input_211;
      end
      8'b11010100 : begin
        result = input_212;
      end
      8'b11010101 : begin
        result = input_213;
      end
      8'b11010110 : begin
        result = input_214;
      end
      8'b11010111 : begin
        result = input_215;
      end
      8'b11011000 : begin
        result = input_216;
      end
      8'b11011001 : begin
        result = input_217;
      end
      8'b11011010 : begin
        result = input_218;
      end
      8'b11011011 : begin
        result = input_219;
      end
      8'b11011100 : begin
        result = input_220;
      end
      8'b11011101 : begin
        result = input_221;
      end
      8'b11011110 : begin
        result = input_222;
      end
      8'b11011111 : begin
        result = input_223;
      end
      8'b11100000 : begin
        result = input_224;
      end
      8'b11100001 : begin
        result = input_225;
      end
      8'b11100010 : begin
        result = input_226;
      end
      8'b11100011 : begin
        result = input_227;
      end
      8'b11100100 : begin
        result = input_228;
      end
      8'b11100101 : begin
        result = input_229;
      end
      8'b11100110 : begin
        result = input_230;
      end
      8'b11100111 : begin
        result = input_231;
      end
      8'b11101000 : begin
        result = input_232;
      end
      8'b11101001 : begin
        result = input_233;
      end
      8'b11101010 : begin
        result = input_234;
      end
      8'b11101011 : begin
        result = input_235;
      end
      8'b11101100 : begin
        result = input_236;
      end
      8'b11101101 : begin
        result = input_237;
      end
      8'b11101110 : begin
        result = input_238;
      end
      8'b11101111 : begin
        result = input_239;
      end
      8'b11110000 : begin
        result = input_240;
      end
      8'b11110001 : begin
        result = input_241;
      end
      8'b11110010 : begin
        result = input_242;
      end
      8'b11110011 : begin
        result = input_243;
      end
      8'b11110100 : begin
        result = input_244;
      end
      8'b11110101 : begin
        result = input_245;
      end
      8'b11110110 : begin
        result = input_246;
      end
      8'b11110111 : begin
        result = input_247;
      end
      8'b11111000 : begin
        result = input_248;
      end
      8'b11111001 : begin
        result = input_249;
      end
      8'b11111010 : begin
        result = input_250;
      end
      8'b11111011 : begin
        result = input_251;
      end
      8'b11111100 : begin
        result = input_252;
      end
      8'b11111101 : begin
        result = input_253;
      end
      8'b11111110 : begin
        result = input_254;
      end
      default : begin
        result = input_255;
      end
    endcase
    MUX_v_64_256_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input  sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function automatic [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input  sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input  sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_8_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [7:0] input_2;
    input [7:0] input_3;
    input [7:0] input_4;
    input [7:0] input_5;
    input [7:0] input_6;
    input [7:0] input_7;
    input [2:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_8_8_2 = result;
  end
  endfunction


  function automatic [19:0] readslicef_31_20_11;
    input [30:0] vector;
    reg [30:0] tmp;
  begin
    tmp = vector >> 11;
    readslicef_31_20_11 = tmp[19:0];
  end
  endfunction


  function automatic [10:0] signext_11_1;
    input  vector;
  begin
    signext_11_1= {{10{vector}}, vector};
  end
  endfunction


  function automatic [255:0] signext_256_244;
    input [243:0] vector;
  begin
    signext_256_244= {{12{vector[243]}}, vector};
  end
  endfunction


  function automatic [1:0] signext_2_1;
    input  vector;
  begin
    signext_2_1= {{1{vector}}, vector};
  end
  endfunction


  function automatic [3:0] signext_4_1;
    input  vector;
  begin
    signext_4_1= {{3{vector}}, vector};
  end
  endfunction


  function automatic [4:0] signext_5_1;
    input  vector;
  begin
    signext_5_1= {{4{vector}}, vector};
  end
  endfunction


  function automatic [6:0] signext_7_1;
    input  vector;
  begin
    signext_7_1= {{6{vector}}, vector};
  end
  endfunction


  function automatic [4:0] conv_u2s_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2s_4_5 =  {1'b0, vector};
  end
  endfunction


  function automatic [8:0] conv_u2s_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2s_8_9 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    PECore
// ------------------------------------------------------------------


module PECore (
  clk, rst, start_vld, start_rdy, start_dat, input_port_vld, input_port_rdy, input_port_dat,
      rva_in_vld, rva_in_rdy, rva_in_dat, rva_out_vld, rva_out_rdy, rva_out_dat,
      act_port_vld, act_port_rdy, act_port_dat, SC_SRAM_CONFIG
);
  input clk;
  input rst;
  input start_vld;
  output start_rdy;
  input start_dat;
  input input_port_vld;
  output input_port_rdy;
  input [73:0] input_port_dat;
  input rva_in_vld;
  output rva_in_rdy;
  input [96:0] rva_in_dat;
  output rva_out_vld;
  input rva_out_rdy;
  output [63:0] rva_out_dat;
  output act_port_vld;
  input act_port_rdy;
  output [255:0] act_port_dat;
  input [31:0] SC_SRAM_CONFIG;


  // Interconnect Declarations
  wire weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d;
  wire [63:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_d_d;
  wire [63:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_radr_d;
  wire weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d;
  wire [63:0] weight_mem_banks_bank_a0_a0_a1_a_rsci_d_d;
  wire [63:0] weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a0_a0_a1_a_rsci_radr_d;
  wire weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d;
  wire [63:0] weight_mem_banks_bank_a0_a1_a0_a_rsci_d_d;
  wire [63:0] weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a0_a1_a0_a_rsci_radr_d;
  wire weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d;
  wire [63:0] weight_mem_banks_bank_a0_a1_a1_a_rsci_d_d;
  wire [63:0] weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a0_a1_a1_a_rsci_radr_d;
  wire weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d;
  wire [63:0] weight_mem_banks_bank_a1_a0_a0_a_rsci_d_d;
  wire [63:0] weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a1_a0_a0_a_rsci_radr_d;
  wire weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d;
  wire [63:0] weight_mem_banks_bank_a1_a0_a1_a_rsci_d_d;
  wire [63:0] weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a1_a0_a1_a_rsci_radr_d;
  wire weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d;
  wire [63:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_d_d;
  wire [63:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_radr_d;
  wire weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d;
  wire [63:0] weight_mem_banks_bank_a1_a1_a1_a_rsci_d_d;
  wire [63:0] weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d;
  wire [11:0] weight_mem_banks_bank_a1_a1_a1_a_rsci_radr_d;
  wire [7:0] ProductSum_for_acc_11_cmp_a;
  wire ProductSum_for_acc_11_cmp_en;
  wire [22:0] ProductSum_for_acc_11_cmp_z;
  wire [7:0] ProductSum_for_acc_10_cmp_a;
  wire [22:0] ProductSum_for_acc_10_cmp_z;
  wire [7:0] ProductSum_for_acc_9_cmp_a0;
  wire [7:0] ProductSum_for_acc_9_cmp_b0;
  wire [7:0] ProductSum_for_acc_9_cmp_c0;
  wire ProductSum_for_acc_9_cmp_en;
  wire [22:0] ProductSum_for_acc_9_cmp_z;
  wire [7:0] ProductSum_for_acc_8_cmp_a0;
  wire [7:0] ProductSum_for_acc_8_cmp_b0;
  wire [7:0] ProductSum_for_acc_8_cmp_c0;
  wire [22:0] ProductSum_for_acc_8_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_a;
  wire [22:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_4_cmp_a;
  wire [22:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_4_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_c0;
  wire [22:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_c0;
  wire [22:0] PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_a;
  wire [22:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_4_cmp_a;
  wire [22:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_4_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_c0;
  wire [22:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_c0;
  wire [22:0] PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_a;
  wire [22:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_4_cmp_a;
  wire [22:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_4_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_c0;
  wire [22:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_c0;
  wire [22:0] PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_a;
  wire [22:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_4_cmp_a;
  wire [22:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_4_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_c0;
  wire [22:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_c0;
  wire [22:0] PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_a;
  wire PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_load;
  wire [22:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_a;
  wire [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_b;
  wire [22:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_c0;
  wire [22:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_c0;
  wire [22:0] PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_a;
  wire [22:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_4_cmp_a;
  wire [22:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_4_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_c0;
  wire [22:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_c0;
  wire [22:0] PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_a;
  wire [22:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_a;
  wire [22:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_c0;
  wire [22:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_z;
  wire [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_a0;
  wire [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_b0;
  wire [7:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_c0;
  wire [22:0] PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_z;
  wire weight_mem_banks_bank_a0_a0_a0_a_rsc_clken;
  wire [63:0] weight_mem_banks_bank_a0_a0_a0_a_rsc_q;
  wire weight_mem_banks_bank_a0_a0_a0_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a0_a0_a0_a_rsc_radr;
  wire weight_mem_banks_bank_a0_a0_a0_a_rsc_we;
  wire [63:0] weight_mem_banks_bank_a0_a0_a0_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a0_a0_a0_a_rsc_wadr;
  wire weight_mem_banks_bank_a0_a0_a1_a_rsc_clken;
  wire [63:0] weight_mem_banks_bank_a0_a0_a1_a_rsc_q;
  wire weight_mem_banks_bank_a0_a0_a1_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a0_a0_a1_a_rsc_radr;
  wire weight_mem_banks_bank_a0_a0_a1_a_rsc_we;
  wire [63:0] weight_mem_banks_bank_a0_a0_a1_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a0_a0_a1_a_rsc_wadr;
  wire weight_mem_banks_bank_a0_a1_a0_a_rsc_clken;
  wire [63:0] weight_mem_banks_bank_a0_a1_a0_a_rsc_q;
  wire weight_mem_banks_bank_a0_a1_a0_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a0_a1_a0_a_rsc_radr;
  wire weight_mem_banks_bank_a0_a1_a0_a_rsc_we;
  wire [63:0] weight_mem_banks_bank_a0_a1_a0_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a0_a1_a0_a_rsc_wadr;
  wire weight_mem_banks_bank_a0_a1_a1_a_rsc_clken;
  wire [63:0] weight_mem_banks_bank_a0_a1_a1_a_rsc_q;
  wire weight_mem_banks_bank_a0_a1_a1_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a0_a1_a1_a_rsc_radr;
  wire weight_mem_banks_bank_a0_a1_a1_a_rsc_we;
  wire [63:0] weight_mem_banks_bank_a0_a1_a1_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a0_a1_a1_a_rsc_wadr;
  wire weight_mem_banks_bank_a1_a0_a0_a_rsc_clken;
  wire [63:0] weight_mem_banks_bank_a1_a0_a0_a_rsc_q;
  wire weight_mem_banks_bank_a1_a0_a0_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a1_a0_a0_a_rsc_radr;
  wire weight_mem_banks_bank_a1_a0_a0_a_rsc_we;
  wire [63:0] weight_mem_banks_bank_a1_a0_a0_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a1_a0_a0_a_rsc_wadr;
  wire weight_mem_banks_bank_a1_a0_a1_a_rsc_clken;
  wire [63:0] weight_mem_banks_bank_a1_a0_a1_a_rsc_q;
  wire weight_mem_banks_bank_a1_a0_a1_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a1_a0_a1_a_rsc_radr;
  wire weight_mem_banks_bank_a1_a0_a1_a_rsc_we;
  wire [63:0] weight_mem_banks_bank_a1_a0_a1_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a1_a0_a1_a_rsc_wadr;
  wire weight_mem_banks_bank_a1_a1_a0_a_rsc_clken;
  wire [63:0] weight_mem_banks_bank_a1_a1_a0_a_rsc_q;
  wire weight_mem_banks_bank_a1_a1_a0_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a1_a1_a0_a_rsc_radr;
  wire weight_mem_banks_bank_a1_a1_a0_a_rsc_we;
  wire [63:0] weight_mem_banks_bank_a1_a1_a0_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a1_a1_a0_a_rsc_wadr;
  wire weight_mem_banks_bank_a1_a1_a1_a_rsc_clken;
  wire [63:0] weight_mem_banks_bank_a1_a1_a1_a_rsc_q;
  wire weight_mem_banks_bank_a1_a1_a1_a_rsc_re;
  wire [11:0] weight_mem_banks_bank_a1_a1_a1_a_rsc_radr;
  wire weight_mem_banks_bank_a1_a1_a1_a_rsc_we;
  wire [63:0] weight_mem_banks_bank_a1_a1_a1_a_rsc_d;
  wire [11:0] weight_mem_banks_bank_a1_a1_a1_a_rsc_wadr;
  wire [7:0] ProductSum_for_acc_11_cmp_b_iff;
  wire ProductSum_for_acc_11_cmp_load_iff;
  wire ProductSum_for_acc_11_cmp_datavalid_iff;
  wire [7:0] ProductSum_for_acc_10_cmp_b_iff;
  wire [7:0] ProductSum_for_acc_9_cmp_a1_iff;
  wire [7:0] ProductSum_for_acc_9_cmp_b1_iff;
  wire [7:0] ProductSum_for_acc_9_cmp_c1_iff;
  wire ProductSum_for_acc_9_cmp_load_iff;
  wire ProductSum_for_acc_9_cmp_datavalid_iff;
  wire [7:0] ProductSum_for_acc_8_cmp_a1_iff;
  wire [7:0] ProductSum_for_acc_8_cmp_b1_iff;
  wire [7:0] ProductSum_for_acc_8_cmp_c1_iff;
  wire PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_load_iff;
  wire PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_load_iff;
  wire PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_load_iff;
  wire PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_load_iff;
  wire PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_load_iff;
  wire PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_load_iff;
  wire PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_load_iff;
  wire PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_load_iff;
  wire PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_load_iff;
  wire PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_load_iff;
  wire PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_load_iff;
  wire PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_load_iff;
  wire PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_load_iff;
  wire weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_iff;
  wire [11:0] weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff;
  wire weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_iff;
  wire weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_iff;
  wire weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_iff;
  wire weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_iff;
  wire weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_iff;
  wire weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_iff;
  wire weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_iff;
  wire weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_iff;
  wire weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_iff;
  wire weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_iff;
  wire weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_iff;
  wire weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_iff;
  wire [11:0] weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_iff;
  wire weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_iff;
  wire weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_iff;
  wire weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_iff;


  // Interconnect Declarations for Component Instantiations 
  PECore_mgc_mulacc_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd23),
  .signd_c(32'sd1),
  .width_d(32'sd0),
  .signd_d(32'sd1),
  .width_z(32'sd23),
  .add_d(32'sd1),
  .is_square(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) ProductSum_for_acc_11_cmp (
      .a(ProductSum_for_acc_11_cmp_a),
      .b(ProductSum_for_acc_11_cmp_b_iff),
      .c(23'b00000000000000000000000),
      .load(ProductSum_for_acc_11_cmp_load_iff),
      .datavalid(ProductSum_for_acc_11_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_11_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(ProductSum_for_acc_11_cmp_z),
      .d(2'b0)
    );
  PECore_mgc_mulacc_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd23),
  .signd_c(32'sd1),
  .width_d(32'sd0),
  .signd_d(32'sd1),
  .width_z(32'sd23),
  .add_d(32'sd1),
  .is_square(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) ProductSum_for_acc_10_cmp (
      .a(ProductSum_for_acc_10_cmp_a),
      .b(ProductSum_for_acc_10_cmp_b_iff),
      .c(23'b00000000000000000000000),
      .load(ProductSum_for_acc_11_cmp_load_iff),
      .datavalid(ProductSum_for_acc_11_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_11_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(ProductSum_for_acc_10_cmp_z),
      .d(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd23),
  .signd_e(32'sd1),
  .width_z(32'sd23),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) ProductSum_for_acc_9_cmp (
      .a0(ProductSum_for_acc_9_cmp_a0),
      .a1(ProductSum_for_acc_9_cmp_a1_iff),
      .b0(ProductSum_for_acc_9_cmp_b0),
      .b1(ProductSum_for_acc_9_cmp_b1_iff),
      .c0(ProductSum_for_acc_9_cmp_c0),
      .c1(ProductSum_for_acc_9_cmp_c1_iff),
      .e(23'b00000000000000000000000),
      .load(ProductSum_for_acc_9_cmp_load_iff),
      .datavalid(ProductSum_for_acc_9_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(ProductSum_for_acc_9_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd23),
  .signd_e(32'sd1),
  .width_z(32'sd23),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) ProductSum_for_acc_8_cmp (
      .a0(ProductSum_for_acc_8_cmp_a0),
      .a1(ProductSum_for_acc_8_cmp_a1_iff),
      .b0(ProductSum_for_acc_8_cmp_b0),
      .b1(ProductSum_for_acc_8_cmp_b1_iff),
      .c0(ProductSum_for_acc_8_cmp_c0),
      .c1(ProductSum_for_acc_8_cmp_c1_iff),
      .e(23'b00000000000000000000000),
      .load(ProductSum_for_acc_9_cmp_load_iff),
      .datavalid(ProductSum_for_acc_9_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(ProductSum_for_acc_8_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mulacc_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd23),
  .signd_c(32'sd1),
  .width_d(32'sd0),
  .signd_d(32'sd1),
  .width_z(32'sd23),
  .add_d(32'sd1),
  .is_square(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp (
      .a(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_a),
      .b(ProductSum_for_acc_11_cmp_b_iff),
      .c(23'b00000000000000000000000),
      .load(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_load_iff),
      .datavalid(ProductSum_for_acc_11_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_11_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_z),
      .d(2'b0)
    );
  PECore_mgc_mulacc_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd23),
  .signd_c(32'sd1),
  .width_d(32'sd0),
  .signd_d(32'sd1),
  .width_z(32'sd23),
  .add_d(32'sd1),
  .is_square(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_4_cmp (
      .a(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_4_cmp_a),
      .b(ProductSum_for_acc_10_cmp_b_iff),
      .c(23'b00000000000000000000000),
      .load(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_load_iff),
      .datavalid(ProductSum_for_acc_11_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_11_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_4_cmp_z),
      .d(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd23),
  .signd_e(32'sd1),
  .width_z(32'sd23),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp (
      .a0(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_a0),
      .a1(ProductSum_for_acc_9_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_b0),
      .b1(ProductSum_for_acc_9_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_c0),
      .c1(ProductSum_for_acc_9_cmp_c1_iff),
      .e(23'b00000000000000000000000),
      .load(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_load_iff),
      .datavalid(ProductSum_for_acc_9_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd23),
  .signd_e(32'sd1),
  .width_z(32'sd23),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp (
      .a0(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_a0),
      .a1(ProductSum_for_acc_8_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_b0),
      .b1(ProductSum_for_acc_8_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_c0),
      .c1(ProductSum_for_acc_8_cmp_c1_iff),
      .e(23'b00000000000000000000000),
      .load(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_load_iff),
      .datavalid(ProductSum_for_acc_9_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mulacc_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd23),
  .signd_c(32'sd1),
  .width_d(32'sd0),
  .signd_d(32'sd1),
  .width_z(32'sd23),
  .add_d(32'sd1),
  .is_square(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp (
      .a(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_a),
      .b(ProductSum_for_acc_11_cmp_b_iff),
      .c(23'b00000000000000000000000),
      .load(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_load_iff),
      .datavalid(ProductSum_for_acc_11_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_11_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_z),
      .d(2'b0)
    );
  PECore_mgc_mulacc_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd23),
  .signd_c(32'sd1),
  .width_d(32'sd0),
  .signd_d(32'sd1),
  .width_z(32'sd23),
  .add_d(32'sd1),
  .is_square(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_4_cmp (
      .a(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_4_cmp_a),
      .b(ProductSum_for_acc_10_cmp_b_iff),
      .c(23'b00000000000000000000000),
      .load(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_load_iff),
      .datavalid(ProductSum_for_acc_11_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_11_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_4_cmp_z),
      .d(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd23),
  .signd_e(32'sd1),
  .width_z(32'sd23),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp (
      .a0(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_a0),
      .a1(ProductSum_for_acc_9_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_b0),
      .b1(ProductSum_for_acc_9_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_c0),
      .c1(ProductSum_for_acc_9_cmp_c1_iff),
      .e(23'b00000000000000000000000),
      .load(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_load_iff),
      .datavalid(ProductSum_for_acc_9_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd23),
  .signd_e(32'sd1),
  .width_z(32'sd23),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp (
      .a0(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_a0),
      .a1(ProductSum_for_acc_8_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_b0),
      .b1(ProductSum_for_acc_8_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_c0),
      .c1(ProductSum_for_acc_8_cmp_c1_iff),
      .e(23'b00000000000000000000000),
      .load(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_load_iff),
      .datavalid(ProductSum_for_acc_9_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mulacc_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd23),
  .signd_c(32'sd1),
  .width_d(32'sd0),
  .signd_d(32'sd1),
  .width_z(32'sd23),
  .add_d(32'sd1),
  .is_square(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp (
      .a(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_a),
      .b(ProductSum_for_acc_11_cmp_b_iff),
      .c(23'b00000000000000000000000),
      .load(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_load_iff),
      .datavalid(ProductSum_for_acc_11_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_11_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_z),
      .d(2'b0)
    );
  PECore_mgc_mulacc_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd23),
  .signd_c(32'sd1),
  .width_d(32'sd0),
  .signd_d(32'sd1),
  .width_z(32'sd23),
  .add_d(32'sd1),
  .is_square(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_4_cmp (
      .a(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_4_cmp_a),
      .b(ProductSum_for_acc_10_cmp_b_iff),
      .c(23'b00000000000000000000000),
      .load(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_load_iff),
      .datavalid(ProductSum_for_acc_11_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_11_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_4_cmp_z),
      .d(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd23),
  .signd_e(32'sd1),
  .width_z(32'sd23),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp (
      .a0(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_a0),
      .a1(ProductSum_for_acc_9_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_b0),
      .b1(ProductSum_for_acc_9_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_c0),
      .c1(ProductSum_for_acc_9_cmp_c1_iff),
      .e(23'b00000000000000000000000),
      .load(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_load_iff),
      .datavalid(ProductSum_for_acc_9_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd23),
  .signd_e(32'sd1),
  .width_z(32'sd23),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp (
      .a0(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_a0),
      .a1(ProductSum_for_acc_8_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_b0),
      .b1(ProductSum_for_acc_8_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_c0),
      .c1(ProductSum_for_acc_8_cmp_c1_iff),
      .e(23'b00000000000000000000000),
      .load(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_load_iff),
      .datavalid(ProductSum_for_acc_9_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mulacc_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd23),
  .signd_c(32'sd1),
  .width_d(32'sd0),
  .signd_d(32'sd1),
  .width_z(32'sd23),
  .add_d(32'sd1),
  .is_square(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp (
      .a(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_a),
      .b(ProductSum_for_acc_11_cmp_b_iff),
      .c(23'b00000000000000000000000),
      .load(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_load_iff),
      .datavalid(ProductSum_for_acc_11_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_11_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_z),
      .d(2'b0)
    );
  PECore_mgc_mulacc_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd23),
  .signd_c(32'sd1),
  .width_d(32'sd0),
  .signd_d(32'sd1),
  .width_z(32'sd23),
  .add_d(32'sd1),
  .is_square(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_4_cmp (
      .a(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_4_cmp_a),
      .b(ProductSum_for_acc_10_cmp_b_iff),
      .c(23'b00000000000000000000000),
      .load(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_load_iff),
      .datavalid(ProductSum_for_acc_11_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_11_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_4_cmp_z),
      .d(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd23),
  .signd_e(32'sd1),
  .width_z(32'sd23),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp (
      .a0(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_a0),
      .a1(ProductSum_for_acc_9_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_b0),
      .b1(ProductSum_for_acc_9_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_c0),
      .c1(ProductSum_for_acc_9_cmp_c1_iff),
      .e(23'b00000000000000000000000),
      .load(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_load_iff),
      .datavalid(ProductSum_for_acc_9_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd23),
  .signd_e(32'sd1),
  .width_z(32'sd23),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp (
      .a0(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_a0),
      .a1(ProductSum_for_acc_8_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_b0),
      .b1(ProductSum_for_acc_8_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_c0),
      .c1(ProductSum_for_acc_8_cmp_c1_iff),
      .e(23'b00000000000000000000000),
      .load(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_load_iff),
      .datavalid(ProductSum_for_acc_9_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mulacc_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd23),
  .signd_c(32'sd1),
  .width_d(32'sd0),
  .signd_d(32'sd1),
  .width_z(32'sd23),
  .add_d(32'sd1),
  .is_square(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp (
      .a(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_a),
      .b(ProductSum_for_acc_11_cmp_b_iff),
      .c(23'b00000000000000000000000),
      .load(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_load),
      .datavalid(ProductSum_for_acc_11_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_11_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_z),
      .d(2'b0)
    );
  PECore_mgc_mulacc_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd23),
  .signd_c(32'sd1),
  .width_d(32'sd0),
  .signd_d(32'sd1),
  .width_z(32'sd23),
  .add_d(32'sd1),
  .is_square(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp (
      .a(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_a),
      .b(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_b),
      .c(23'b00000000000000000000000),
      .load(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_load_iff),
      .datavalid(ProductSum_for_acc_9_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_z),
      .d(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd23),
  .signd_e(32'sd1),
  .width_z(32'sd23),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp (
      .a0(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_a0),
      .a1(ProductSum_for_acc_9_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_b0),
      .b1(ProductSum_for_acc_9_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_c0),
      .c1(ProductSum_for_acc_9_cmp_c1_iff),
      .e(23'b00000000000000000000000),
      .load(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_load_iff),
      .datavalid(ProductSum_for_acc_9_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd23),
  .signd_e(32'sd1),
  .width_z(32'sd23),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp (
      .a0(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_a0),
      .a1(ProductSum_for_acc_8_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_b0),
      .b1(ProductSum_for_acc_8_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_c0),
      .c1(ProductSum_for_acc_8_cmp_c1_iff),
      .e(23'b00000000000000000000000),
      .load(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_load_iff),
      .datavalid(ProductSum_for_acc_9_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mulacc_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd23),
  .signd_c(32'sd1),
  .width_d(32'sd0),
  .signd_d(32'sd1),
  .width_z(32'sd23),
  .add_d(32'sd1),
  .is_square(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp (
      .a(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_a),
      .b(ProductSum_for_acc_11_cmp_b_iff),
      .c(23'b00000000000000000000000),
      .load(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_load_iff),
      .datavalid(ProductSum_for_acc_11_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_11_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_z),
      .d(2'b0)
    );
  PECore_mgc_mulacc_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd23),
  .signd_c(32'sd1),
  .width_d(32'sd0),
  .signd_d(32'sd1),
  .width_z(32'sd23),
  .add_d(32'sd1),
  .is_square(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_4_cmp (
      .a(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_4_cmp_a),
      .b(ProductSum_for_acc_10_cmp_b_iff),
      .c(23'b00000000000000000000000),
      .load(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_load_iff),
      .datavalid(ProductSum_for_acc_11_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_11_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_4_cmp_z),
      .d(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd23),
  .signd_e(32'sd1),
  .width_z(32'sd23),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp (
      .a0(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_a0),
      .a1(ProductSum_for_acc_9_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_b0),
      .b1(ProductSum_for_acc_9_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_c0),
      .c1(ProductSum_for_acc_9_cmp_c1_iff),
      .e(23'b00000000000000000000000),
      .load(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_load_iff),
      .datavalid(ProductSum_for_acc_9_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd23),
  .signd_e(32'sd1),
  .width_z(32'sd23),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp (
      .a0(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_a0),
      .a1(ProductSum_for_acc_8_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_b0),
      .b1(ProductSum_for_acc_8_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_c0),
      .c1(ProductSum_for_acc_8_cmp_c1_iff),
      .e(23'b00000000000000000000000),
      .load(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_load_iff),
      .datavalid(ProductSum_for_acc_9_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mulacc_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd23),
  .signd_c(32'sd1),
  .width_d(32'sd0),
  .signd_d(32'sd1),
  .width_z(32'sd23),
  .add_d(32'sd1),
  .is_square(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp (
      .a(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_a),
      .b(ProductSum_for_acc_11_cmp_b_iff),
      .c(23'b00000000000000000000000),
      .load(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_load_iff),
      .datavalid(ProductSum_for_acc_11_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_11_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_z),
      .d(2'b0)
    );
  PECore_mgc_mulacc_pipe #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_b(32'sd8),
  .signd_b(32'sd0),
  .width_c(32'sd23),
  .signd_c(32'sd1),
  .width_d(32'sd0),
  .signd_d(32'sd1),
  .width_z(32'sd23),
  .add_d(32'sd1),
  .is_square(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp (
      .a(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_a),
      .b(ProductSum_for_acc_10_cmp_b_iff),
      .c(23'b00000000000000000000000),
      .load(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_load_iff),
      .datavalid(ProductSum_for_acc_11_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_11_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_z),
      .d(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd23),
  .signd_e(32'sd1),
  .width_z(32'sd23),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp (
      .a0(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_a0),
      .a1(ProductSum_for_acc_9_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_b0),
      .b1(ProductSum_for_acc_9_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_c0),
      .c1(ProductSum_for_acc_9_cmp_c1_iff),
      .e(23'b00000000000000000000000),
      .load(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_load_iff),
      .datavalid(ProductSum_for_acc_9_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  PECore_mgc_mul4acc_pipe #(.width_a0(32'sd8),
  .signd_a0(32'sd0),
  .width_a1(32'sd8),
  .signd_a1(32'sd0),
  .width_b0(32'sd8),
  .signd_b0(32'sd0),
  .width_b1(32'sd8),
  .signd_b1(32'sd0),
  .width_c0(32'sd8),
  .signd_c0(32'sd0),
  .width_c1(32'sd8),
  .signd_c1(32'sd0),
  .width_d0(32'sd0),
  .signd_d0(32'sd0),
  .width_d1(32'sd0),
  .signd_d1(32'sd0),
  .width_e(32'sd23),
  .signd_e(32'sd1),
  .width_z(32'sd23),
  .add_a(32'sd1),
  .add_b(32'sd1),
  .add_c(32'sd1),
  .min_fb_size(32'sd0),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp (
      .a0(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_a0),
      .a1(ProductSum_for_acc_8_cmp_a1_iff),
      .b0(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_b0),
      .b1(ProductSum_for_acc_8_cmp_b1_iff),
      .c0(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_c0),
      .c1(ProductSum_for_acc_8_cmp_c1_iff),
      .e(23'b00000000000000000000000),
      .load(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_load_iff),
      .datavalid(ProductSum_for_acc_9_cmp_datavalid_iff),
      .clk(clk),
      .en(ProductSum_for_acc_9_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_z),
      .d0(2'b0),
      .d1(2'b0)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd64),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a0_a0_a0_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a0_a0_a0_a_rsc_clken),
      .d(weight_mem_banks_bank_a0_a0_a0_a_rsc_d),
      .q(weight_mem_banks_bank_a0_a0_a0_a_rsc_q),
      .radr(weight_mem_banks_bank_a0_a0_a0_a_rsc_radr),
      .re(weight_mem_banks_bank_a0_a0_a0_a_rsc_re),
      .wadr(weight_mem_banks_bank_a0_a0_a0_a_rsc_wadr),
      .we(weight_mem_banks_bank_a0_a0_a0_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd64),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a0_a0_a1_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a0_a0_a1_a_rsc_clken),
      .d(weight_mem_banks_bank_a0_a0_a1_a_rsc_d),
      .q(weight_mem_banks_bank_a0_a0_a1_a_rsc_q),
      .radr(weight_mem_banks_bank_a0_a0_a1_a_rsc_radr),
      .re(weight_mem_banks_bank_a0_a0_a1_a_rsc_re),
      .wadr(weight_mem_banks_bank_a0_a0_a1_a_rsc_wadr),
      .we(weight_mem_banks_bank_a0_a0_a1_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd64),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a0_a1_a0_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a0_a1_a0_a_rsc_clken),
      .d(weight_mem_banks_bank_a0_a1_a0_a_rsc_d),
      .q(weight_mem_banks_bank_a0_a1_a0_a_rsc_q),
      .radr(weight_mem_banks_bank_a0_a1_a0_a_rsc_radr),
      .re(weight_mem_banks_bank_a0_a1_a0_a_rsc_re),
      .wadr(weight_mem_banks_bank_a0_a1_a0_a_rsc_wadr),
      .we(weight_mem_banks_bank_a0_a1_a0_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd64),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a0_a1_a1_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a0_a1_a1_a_rsc_clken),
      .d(weight_mem_banks_bank_a0_a1_a1_a_rsc_d),
      .q(weight_mem_banks_bank_a0_a1_a1_a_rsc_q),
      .radr(weight_mem_banks_bank_a0_a1_a1_a_rsc_radr),
      .re(weight_mem_banks_bank_a0_a1_a1_a_rsc_re),
      .wadr(weight_mem_banks_bank_a0_a1_a1_a_rsc_wadr),
      .we(weight_mem_banks_bank_a0_a1_a1_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd64),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a1_a0_a0_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a1_a0_a0_a_rsc_clken),
      .d(weight_mem_banks_bank_a1_a0_a0_a_rsc_d),
      .q(weight_mem_banks_bank_a1_a0_a0_a_rsc_q),
      .radr(weight_mem_banks_bank_a1_a0_a0_a_rsc_radr),
      .re(weight_mem_banks_bank_a1_a0_a0_a_rsc_re),
      .wadr(weight_mem_banks_bank_a1_a0_a0_a_rsc_wadr),
      .we(weight_mem_banks_bank_a1_a0_a0_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd64),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a1_a0_a1_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a1_a0_a1_a_rsc_clken),
      .d(weight_mem_banks_bank_a1_a0_a1_a_rsc_d),
      .q(weight_mem_banks_bank_a1_a0_a1_a_rsc_q),
      .radr(weight_mem_banks_bank_a1_a0_a1_a_rsc_radr),
      .re(weight_mem_banks_bank_a1_a0_a1_a_rsc_re),
      .wadr(weight_mem_banks_bank_a1_a0_a1_a_rsc_wadr),
      .we(weight_mem_banks_bank_a1_a0_a1_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd64),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a1_a1_a0_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a1_a1_a0_a_rsc_clken),
      .d(weight_mem_banks_bank_a1_a1_a0_a_rsc_d),
      .q(weight_mem_banks_bank_a1_a1_a0_a_rsc_q),
      .radr(weight_mem_banks_bank_a1_a1_a0_a_rsc_radr),
      .re(weight_mem_banks_bank_a1_a1_a0_a_rsc_re),
      .wadr(weight_mem_banks_bank_a1_a1_a0_a_rsc_wadr),
      .we(weight_mem_banks_bank_a1_a1_a0_a_rsc_we)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd12),
  .data_width(32'sd64),
  .depth(32'sd4096),
  .latency(32'sd1),
  .suppress_sim_read_addr_range_errs(32'sd1)) weight_mem_banks_bank_a1_a1_a1_a_rsc_comp
      (
      .clk(clk),
      .clken(weight_mem_banks_bank_a1_a1_a1_a_rsc_clken),
      .d(weight_mem_banks_bank_a1_a1_a1_a_rsc_d),
      .q(weight_mem_banks_bank_a1_a1_a1_a_rsc_q),
      .radr(weight_mem_banks_bank_a1_a1_a1_a_rsc_radr),
      .re(weight_mem_banks_bank_a1_a1_a1_a_rsc_re),
      .wadr(weight_mem_banks_bank_a1_a1_a1_a_rsc_wadr),
      .we(weight_mem_banks_bank_a1_a1_a1_a_rsc_we)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_139_12_64_4096_1_4096_64_1_gen
      weight_mem_banks_bank_a0_a0_a0_a_rsci (
      .clken(weight_mem_banks_bank_a0_a0_a0_a_rsc_clken),
      .q(weight_mem_banks_bank_a0_a0_a0_a_rsc_q),
      .re(weight_mem_banks_bank_a0_a0_a0_a_rsc_re),
      .radr(weight_mem_banks_bank_a0_a0_a0_a_rsc_radr),
      .we(weight_mem_banks_bank_a0_a0_a0_a_rsc_we),
      .d(weight_mem_banks_bank_a0_a0_a0_a_rsc_d),
      .wadr(weight_mem_banks_bank_a0_a0_a0_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_iff)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_140_12_64_4096_1_4096_64_1_gen
      weight_mem_banks_bank_a0_a0_a1_a_rsci (
      .clken(weight_mem_banks_bank_a0_a0_a1_a_rsc_clken),
      .q(weight_mem_banks_bank_a0_a0_a1_a_rsc_q),
      .re(weight_mem_banks_bank_a0_a0_a1_a_rsc_re),
      .radr(weight_mem_banks_bank_a0_a0_a1_a_rsc_radr),
      .we(weight_mem_banks_bank_a0_a0_a1_a_rsc_we),
      .d(weight_mem_banks_bank_a0_a0_a1_a_rsc_d),
      .wadr(weight_mem_banks_bank_a0_a0_a1_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_iff)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_141_12_64_4096_1_4096_64_1_gen
      weight_mem_banks_bank_a0_a1_a0_a_rsci (
      .clken(weight_mem_banks_bank_a0_a1_a0_a_rsc_clken),
      .q(weight_mem_banks_bank_a0_a1_a0_a_rsc_q),
      .re(weight_mem_banks_bank_a0_a1_a0_a_rsc_re),
      .radr(weight_mem_banks_bank_a0_a1_a0_a_rsc_radr),
      .we(weight_mem_banks_bank_a0_a1_a0_a_rsc_we),
      .d(weight_mem_banks_bank_a0_a1_a0_a_rsc_d),
      .wadr(weight_mem_banks_bank_a0_a1_a0_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_iff)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_142_12_64_4096_1_4096_64_1_gen
      weight_mem_banks_bank_a0_a1_a1_a_rsci (
      .clken(weight_mem_banks_bank_a0_a1_a1_a_rsc_clken),
      .q(weight_mem_banks_bank_a0_a1_a1_a_rsc_q),
      .re(weight_mem_banks_bank_a0_a1_a1_a_rsc_re),
      .radr(weight_mem_banks_bank_a0_a1_a1_a_rsc_radr),
      .we(weight_mem_banks_bank_a0_a1_a1_a_rsc_we),
      .d(weight_mem_banks_bank_a0_a1_a1_a_rsc_d),
      .wadr(weight_mem_banks_bank_a0_a1_a1_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_iff)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_143_12_64_4096_1_4096_64_1_gen
      weight_mem_banks_bank_a1_a0_a0_a_rsci (
      .clken(weight_mem_banks_bank_a1_a0_a0_a_rsc_clken),
      .q(weight_mem_banks_bank_a1_a0_a0_a_rsc_q),
      .re(weight_mem_banks_bank_a1_a0_a0_a_rsc_re),
      .radr(weight_mem_banks_bank_a1_a0_a0_a_rsc_radr),
      .we(weight_mem_banks_bank_a1_a0_a0_a_rsc_we),
      .d(weight_mem_banks_bank_a1_a0_a0_a_rsc_d),
      .wadr(weight_mem_banks_bank_a1_a0_a0_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_iff)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_144_12_64_4096_1_4096_64_1_gen
      weight_mem_banks_bank_a1_a0_a1_a_rsci (
      .clken(weight_mem_banks_bank_a1_a0_a1_a_rsc_clken),
      .q(weight_mem_banks_bank_a1_a0_a1_a_rsc_q),
      .re(weight_mem_banks_bank_a1_a0_a1_a_rsc_re),
      .radr(weight_mem_banks_bank_a1_a0_a1_a_rsc_radr),
      .we(weight_mem_banks_bank_a1_a0_a1_a_rsc_we),
      .d(weight_mem_banks_bank_a1_a0_a1_a_rsc_d),
      .wadr(weight_mem_banks_bank_a1_a0_a1_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_iff)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_145_12_64_4096_1_4096_64_1_gen
      weight_mem_banks_bank_a1_a1_a0_a_rsci (
      .clken(weight_mem_banks_bank_a1_a1_a0_a_rsc_clken),
      .q(weight_mem_banks_bank_a1_a1_a0_a_rsc_q),
      .re(weight_mem_banks_bank_a1_a1_a0_a_rsc_re),
      .radr(weight_mem_banks_bank_a1_a1_a0_a_rsc_radr),
      .we(weight_mem_banks_bank_a1_a1_a0_a_rsc_we),
      .d(weight_mem_banks_bank_a1_a1_a0_a_rsc_d),
      .wadr(weight_mem_banks_bank_a1_a1_a0_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_iff)
    );
  PECore_PECore_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_146_12_64_4096_1_4096_64_1_gen
      weight_mem_banks_bank_a1_a1_a1_a_rsci (
      .clken(weight_mem_banks_bank_a1_a1_a1_a_rsc_clken),
      .q(weight_mem_banks_bank_a1_a1_a1_a_rsc_q),
      .re(weight_mem_banks_bank_a1_a1_a1_a_rsc_re),
      .radr(weight_mem_banks_bank_a1_a1_a1_a_rsc_radr),
      .we(weight_mem_banks_bank_a1_a1_a1_a_rsc_we),
      .d(weight_mem_banks_bank_a1_a1_a1_a_rsc_d),
      .wadr(weight_mem_banks_bank_a1_a1_a1_a_rsc_wadr),
      .clken_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d),
      .d_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_d_d),
      .q_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d),
      .radr_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_radr_d),
      .re_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_iff),
      .wadr_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_iff),
      .we_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_iff)
    );
  PECore_PECore_PECoreRun PECore_PECoreRun_inst (
      .clk(clk),
      .rst(rst),
      .start_vld(start_vld),
      .start_rdy(start_rdy),
      .start_dat(start_dat),
      .input_port_vld(input_port_vld),
      .input_port_rdy(input_port_rdy),
      .input_port_dat(input_port_dat),
      .rva_in_vld(rva_in_vld),
      .rva_in_rdy(rva_in_rdy),
      .rva_in_dat(rva_in_dat),
      .rva_out_vld(rva_out_vld),
      .rva_out_rdy(rva_out_rdy),
      .rva_out_dat(rva_out_dat),
      .act_port_vld(act_port_vld),
      .act_port_rdy(act_port_rdy),
      .act_port_dat(act_port_dat),
      .SC_SRAM_CONFIG(SC_SRAM_CONFIG),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_d_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_d_d),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_q_d),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_radr_d(weight_mem_banks_bank_a0_a0_a0_a_rsci_radr_d),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_clken_d),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_d_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_d_d),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_q_d),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_radr_d(weight_mem_banks_bank_a0_a0_a1_a_rsci_radr_d),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_d_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_d_d),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_q_d),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_radr_d(weight_mem_banks_bank_a0_a1_a0_a_rsci_radr_d),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_clken_d),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_d_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_d_d),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_q_d),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_radr_d(weight_mem_banks_bank_a0_a1_a1_a_rsci_radr_d),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_d_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_d_d),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_q_d),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_radr_d(weight_mem_banks_bank_a1_a0_a0_a_rsci_radr_d),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_d_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_d_d),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_q_d),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_radr_d(weight_mem_banks_bank_a1_a0_a1_a_rsci_radr_d),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_d_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_d_d),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_q_d),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_radr_d(weight_mem_banks_bank_a1_a1_a0_a_rsci_radr_d),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_clken_d),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_d_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_d_d),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_q_d),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_radr_d(weight_mem_banks_bank_a1_a1_a1_a_rsci_radr_d),
      .ProductSum_for_acc_11_cmp_a(ProductSum_for_acc_11_cmp_a),
      .ProductSum_for_acc_11_cmp_en(ProductSum_for_acc_11_cmp_en),
      .ProductSum_for_acc_11_cmp_z(ProductSum_for_acc_11_cmp_z),
      .ProductSum_for_acc_10_cmp_a(ProductSum_for_acc_10_cmp_a),
      .ProductSum_for_acc_10_cmp_z(ProductSum_for_acc_10_cmp_z),
      .ProductSum_for_acc_9_cmp_a0(ProductSum_for_acc_9_cmp_a0),
      .ProductSum_for_acc_9_cmp_b0(ProductSum_for_acc_9_cmp_b0),
      .ProductSum_for_acc_9_cmp_c0(ProductSum_for_acc_9_cmp_c0),
      .ProductSum_for_acc_9_cmp_en(ProductSum_for_acc_9_cmp_en),
      .ProductSum_for_acc_9_cmp_z(ProductSum_for_acc_9_cmp_z),
      .ProductSum_for_acc_8_cmp_a0(ProductSum_for_acc_8_cmp_a0),
      .ProductSum_for_acc_8_cmp_b0(ProductSum_for_acc_8_cmp_b0),
      .ProductSum_for_acc_8_cmp_c0(ProductSum_for_acc_8_cmp_c0),
      .ProductSum_for_acc_8_cmp_z(ProductSum_for_acc_8_cmp_z),
      .PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_a(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_a),
      .PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_z(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_z),
      .PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_4_cmp_a(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_4_cmp_a),
      .PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_4_cmp_z(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_4_cmp_z),
      .PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_a0(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_a0),
      .PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_b0(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_b0),
      .PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_c0(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_c0),
      .PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_z(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_z),
      .PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_a0(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_a0),
      .PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_b0(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_b0),
      .PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_c0(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_c0),
      .PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_z(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_2_cmp_z),
      .PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_a(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_a),
      .PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_z(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_z),
      .PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_4_cmp_a(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_4_cmp_a),
      .PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_4_cmp_z(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_4_cmp_z),
      .PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_a0(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_a0),
      .PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_b0(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_b0),
      .PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_c0(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_c0),
      .PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_z(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_z),
      .PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_a0(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_a0),
      .PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_b0(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_b0),
      .PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_c0(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_c0),
      .PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_z(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_2_cmp_z),
      .PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_a(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_a),
      .PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_z(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_z),
      .PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_4_cmp_a(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_4_cmp_a),
      .PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_4_cmp_z(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_4_cmp_z),
      .PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_a0(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_a0),
      .PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_b0(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_b0),
      .PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_c0(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_c0),
      .PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_z(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_z),
      .PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_a0(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_a0),
      .PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_b0(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_b0),
      .PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_c0(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_c0),
      .PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_z(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_2_cmp_z),
      .PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_a(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_a),
      .PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_z(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_z),
      .PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_4_cmp_a(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_4_cmp_a),
      .PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_4_cmp_z(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_4_cmp_z),
      .PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_a0(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_a0),
      .PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_b0(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_b0),
      .PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_c0(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_c0),
      .PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_z(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_z),
      .PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_a0(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_a0),
      .PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_b0(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_b0),
      .PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_c0(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_c0),
      .PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_z(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_2_cmp_z),
      .PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_a(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_a),
      .PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_load(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_load),
      .PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_z(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_5_cmp_z),
      .PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_a(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_a),
      .PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_b(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_b),
      .PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_z(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_z),
      .PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_a0(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_a0),
      .PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_b0(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_b0),
      .PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_c0(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_c0),
      .PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_z(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_3_cmp_z),
      .PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_a0(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_a0),
      .PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_b0(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_b0),
      .PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_c0(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_c0),
      .PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_z(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_2_cmp_z),
      .PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_a(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_a),
      .PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_z(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_z),
      .PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_4_cmp_a(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_4_cmp_a),
      .PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_4_cmp_z(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_4_cmp_z),
      .PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_a0(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_a0),
      .PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_b0(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_b0),
      .PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_c0(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_c0),
      .PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_z(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_z),
      .PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_a0(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_a0),
      .PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_b0(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_b0),
      .PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_c0(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_c0),
      .PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_z(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_2_cmp_z),
      .PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_a(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_a),
      .PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_z(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_z),
      .PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_a(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_a),
      .PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_z(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_4_cmp_z),
      .PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_a0(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_a0),
      .PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_b0(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_b0),
      .PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_c0(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_c0),
      .PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_z(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_z),
      .PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_a0(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_a0),
      .PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_b0(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_b0),
      .PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_c0(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_c0),
      .PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_z(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_2_cmp_z),
      .ProductSum_for_acc_11_cmp_b_pff(ProductSum_for_acc_11_cmp_b_iff),
      .ProductSum_for_acc_11_cmp_load_pff(ProductSum_for_acc_11_cmp_load_iff),
      .ProductSum_for_acc_11_cmp_datavalid_pff(ProductSum_for_acc_11_cmp_datavalid_iff),
      .ProductSum_for_acc_10_cmp_b_pff(ProductSum_for_acc_10_cmp_b_iff),
      .ProductSum_for_acc_9_cmp_a1_pff(ProductSum_for_acc_9_cmp_a1_iff),
      .ProductSum_for_acc_9_cmp_b1_pff(ProductSum_for_acc_9_cmp_b1_iff),
      .ProductSum_for_acc_9_cmp_c1_pff(ProductSum_for_acc_9_cmp_c1_iff),
      .ProductSum_for_acc_9_cmp_load_pff(ProductSum_for_acc_9_cmp_load_iff),
      .ProductSum_for_acc_9_cmp_datavalid_pff(ProductSum_for_acc_9_cmp_datavalid_iff),
      .ProductSum_for_acc_8_cmp_a1_pff(ProductSum_for_acc_8_cmp_a1_iff),
      .ProductSum_for_acc_8_cmp_b1_pff(ProductSum_for_acc_8_cmp_b1_iff),
      .ProductSum_for_acc_8_cmp_c1_pff(ProductSum_for_acc_8_cmp_c1_iff),
      .PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_load_pff(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_5_cmp_load_iff),
      .PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_load_pff(PECore_RunMac_if_for_1_7_PECore_RunMac_if_for_1_acc_3_cmp_load_iff),
      .PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_load_pff(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_5_cmp_load_iff),
      .PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_load_pff(PECore_RunMac_if_for_1_6_PECore_RunMac_if_for_1_acc_3_cmp_load_iff),
      .PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_load_pff(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_5_cmp_load_iff),
      .PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_load_pff(PECore_RunMac_if_for_1_5_PECore_RunMac_if_for_1_acc_3_cmp_load_iff),
      .PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_load_pff(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_5_cmp_load_iff),
      .PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_load_pff(PECore_RunMac_if_for_1_4_PECore_RunMac_if_for_1_acc_3_cmp_load_iff),
      .PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_load_pff(PECore_RunMac_if_for_1_3_PECore_RunMac_if_for_1_acc_4_cmp_load_iff),
      .PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_load_pff(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_5_cmp_load_iff),
      .PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_load_pff(PECore_RunMac_if_for_1_2_PECore_RunMac_if_for_1_acc_3_cmp_load_iff),
      .PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_load_pff(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_5_cmp_load_iff),
      .PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_load_pff(PECore_RunMac_if_for_1_1_PECore_RunMac_if_for_1_acc_3_cmp_load_iff),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_pff(weight_mem_banks_bank_a0_a0_a0_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_pff(weight_mem_banks_bank_a0_a0_a0_a_rsci_wadr_d_iff),
      .weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_pff(weight_mem_banks_bank_a0_a0_a0_a_rsci_we_d_iff),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_pff(weight_mem_banks_bank_a0_a0_a1_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_pff(weight_mem_banks_bank_a0_a0_a1_a_rsci_we_d_iff),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_pff(weight_mem_banks_bank_a0_a1_a0_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_pff(weight_mem_banks_bank_a0_a1_a0_a_rsci_we_d_iff),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_pff(weight_mem_banks_bank_a0_a1_a1_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_pff(weight_mem_banks_bank_a0_a1_a1_a_rsci_we_d_iff),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_pff(weight_mem_banks_bank_a1_a0_a0_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_pff(weight_mem_banks_bank_a1_a0_a0_a_rsci_we_d_iff),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_pff(weight_mem_banks_bank_a1_a0_a1_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_pff(weight_mem_banks_bank_a1_a0_a1_a_rsci_we_d_iff),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_pff(weight_mem_banks_bank_a1_a1_a0_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_pff(weight_mem_banks_bank_a1_a1_a0_a_rsci_wadr_d_iff),
      .weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_pff(weight_mem_banks_bank_a1_a1_a0_a_rsci_we_d_iff),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_pff(weight_mem_banks_bank_a1_a1_a1_a_rsci_re_d_iff),
      .weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_pff(weight_mem_banks_bank_a1_a1_a1_a_rsci_we_d_iff)
    );
endmodule



