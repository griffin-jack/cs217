
//------> ./ActUnit_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ActUnit_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ./ActUnit_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ActUnit_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./ActUnit_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   code@iron-06
//  Generated date: Mon Jan 26 19:49:32 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_core
// ------------------------------------------------------------------


module ActUnit_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_core
    (
  this_vld, this_rdy, this_dat, data_data_rsc_z, data_addr_rsc_z, data_rw_rsc_z,
      return_rsc_z, ccs_ccore_start_rsc_dat, ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  reg this_rdy;
  input [600:0] this_dat;
  output [511:0] data_data_rsc_z;
  output [23:0] data_addr_rsc_z;
  output data_rw_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations
  wire [511:0] nl_data_data_rsci_d;
  assign nl_data_data_rsci_d = this_dat[511:0];
  wire [23:0] nl_data_addr_rsci_d;
  assign nl_data_addr_rsci_d = this_dat[535:512];
  wire  nl_data_rw_rsci_d;
  assign nl_data_rw_rsci_d = this_dat[600];
  ActUnit_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd1),
  .width(32'sd512)) data_data_rsci (
      .d(nl_data_data_rsci_d[511:0]),
      .z(data_data_rsc_z)
    );
  ActUnit_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd2),
  .width(32'sd24)) data_addr_rsci (
      .d(nl_data_addr_rsci_d[23:0]),
      .z(data_addr_rsc_z)
    );
  ActUnit_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd4),
  .width(32'sd1)) data_rw_rsci (
      .d(nl_data_rw_rsci_d),
      .z(data_rw_rsc_z)
    );
  ActUnit_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd6),
  .width(32'sd1)) return_rsci (
      .d(this_vld),
      .z(return_rsc_z)
    );
  ActUnit_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1
      #(.rscid(32'sd58),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_rdy <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB
// ------------------------------------------------------------------


module ActUnit_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB
    (
  this_vld, this_rdy, this_dat, data_data_rsc_z, data_addr_rsc_z, data_rw_rsc_z,
      return_rsc_z, ccs_ccore_start_rsc_dat, ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  input [600:0] this_dat;
  output [511:0] data_data_rsc_z;
  output [23:0] data_addr_rsc_z;
  output data_rw_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  ActUnit_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_core
      Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .data_data_rsc_z(data_data_rsc_z),
      .data_addr_rsc_z(data_addr_rsc_z),
      .data_rw_rsc_z(data_rw_rsc_z),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./ActUnit_Connections_InBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ActUnit_Connections_InBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ./ActUnit_Connections_InBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ActUnit_Connections_InBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./ActUnit_Connections_InBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_PopNB.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   code@iron-06
//  Generated date: Mon Jan 26 19:49:30 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_spec_ActVectorType_Connections_SYN_PORT_PopNB_core
// ------------------------------------------------------------------


module ActUnit_Connections_InBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_spec_ActVectorType_Connections_SYN_PORT_PopNB_core
    (
  this_vld, this_rdy, this_dat, data_data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  reg this_rdy;
  input [511:0] this_dat;
  output [511:0] data_data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations
  ActUnit_Connections_InBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd7),
  .width(32'sd512)) data_data_rsci (
      .d(this_dat),
      .z(data_data_rsc_z)
    );
  ActUnit_Connections_InBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd9),
  .width(32'sd1)) return_rsci (
      .d(this_vld),
      .z(return_rsc_z)
    );
  ActUnit_Connections_InBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1
      #(.rscid(32'sd57),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_rdy <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_spec_ActVectorType_Connections_SYN_PORT_PopNB
// ------------------------------------------------------------------


module ActUnit_Connections_InBlocking_spec_ActVectorType_Connections_SYN_PORT_PopNB (
  this_vld, this_rdy, this_dat, data_data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  input [511:0] this_dat;
  output [511:0] data_data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  ActUnit_Connections_InBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_spec_ActVectorType_Connections_SYN_PORT_PopNB_core
      Connections_InBlocking_spec_ActVectorType_Connections_SYN_PORT_PopNB_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .data_data_rsc_z(data_data_rsc_z),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./ActUnit_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ActUnit_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./ActUnit_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module ActUnit_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./ActUnit_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   code@iron-06
//  Generated date: Mon Jan 26 19:49:27 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module ActUnit_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push_core
    (
  this_vld, this_rdy, this_dat, m_data_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  reg this_vld;
  input this_rdy;
  output [511:0] this_dat;
  reg [511:0] this_dat;
  input [511:0] m_data_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire [511:0] m_data_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  wire and_dcpl;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_4_cse;
  wire this_vld_mx0c1;


  // Interconnect Declarations for Component Instantiations
  wire  nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  ActUnit_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd11),
  .width(32'sd512)) m_data_rsci (
      .dat(m_data_rsc_dat),
      .idat(m_data_rsci_idat)
    );
  ActUnit_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd56),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  ActUnit_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1
      #(.rscid(32'sd61)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld)
    );
  assign or_4_cse = ccs_ccore_start_rsci_idat | and_dcpl;
  assign and_dcpl = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_rdy);
  assign this_vld_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_vld <= 1'b0;
    end
    else if ( or_4_cse | this_vld_mx0c1 ) begin
      this_vld <= ~ this_vld_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_dat <= 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~(and_dcpl | (~ ccs_ccore_start_rsci_idat)) ) begin
      this_dat <= m_data_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_4_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module ActUnit_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push
    (
  this_vld, this_rdy, this_dat, m_data_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  input this_rdy;
  output [511:0] this_dat;
  input [511:0] m_data_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  ActUnit_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push_core
      Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .m_data_rsc_dat(m_data_rsc_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./ActUnit_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ActUnit_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ./ActUnit_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ActUnit_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./ActUnit_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   code@iron-06
//  Generated date: Mon Jan 26 19:49:25 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_core
// ------------------------------------------------------------------


module ActUnit_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_core
    (
  this_vld, this_rdy, this_dat, data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  reg this_rdy;
  input this_dat;
  output data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations
  ActUnit_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd12),
  .width(32'sd1)) data_rsci (
      .d(this_dat),
      .z(data_rsc_z)
    );
  ActUnit_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd14),
  .width(32'sd1)) return_rsci (
      .d(this_vld),
      .z(return_rsc_z)
    );
  ActUnit_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1
      #(.rscid(32'sd55),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_rdy <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_bool_Connections_SYN_PORT_PopNB
// ------------------------------------------------------------------


module ActUnit_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB (
  this_vld, this_rdy, this_dat, data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  input this_dat;
  output data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  ActUnit_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_core
      Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_core_inst (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .data_rsc_z(data_rsc_z),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./ActUnit_Connections_OutBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ActUnit_Connections_OutBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./ActUnit_Connections_OutBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module ActUnit_Connections_OutBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./ActUnit_Connections_OutBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_Push.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   code@iron-06
//  Generated date: Mon Jan 26 19:49:23 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_spec_StreamType_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module ActUnit_Connections_OutBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_spec_StreamType_Connections_SYN_PORT_Push_core
    (
  this_vld, this_rdy, this_dat, m_data_data_rsc_dat, m_logical_addr_rsc_dat, ccs_ccore_start_rsc_dat,
      ccs_ccore_done_sync_vld, ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  reg this_vld;
  input this_rdy;
  output [521:0] this_dat;
  input [511:0] m_data_data_rsc_dat;
  input [7:0] m_logical_addr_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire [511:0] m_data_data_rsci_idat;
  wire [7:0] m_logical_addr_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  reg [7:0] m_logical_addr_buf_lpi_1_dfm;
  reg [511:0] m_data_data_buf_lpi_1_dfm;
  wire and_dcpl;
  wire or_dcpl_2;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_4_cse;
  wire this_vld_mx0c1;


  // Interconnect Declarations for Component Instantiations
  wire  nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  ActUnit_Connections_OutBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd15),
  .width(32'sd512)) m_data_data_rsci (
      .dat(m_data_data_rsc_dat),
      .idat(m_data_data_rsci_idat)
    );
  ActUnit_Connections_OutBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd17),
  .width(32'sd8)) m_logical_addr_rsci (
      .dat(m_logical_addr_rsc_dat),
      .idat(m_logical_addr_rsci_idat)
    );
  ActUnit_Connections_OutBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd54),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  ActUnit_Connections_OutBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1
      #(.rscid(32'sd60)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld)
    );
  assign this_dat = {m_logical_addr_buf_lpi_1_dfm , 2'b00 , m_data_data_buf_lpi_1_dfm};
  assign or_4_cse = ccs_ccore_start_rsci_idat | and_dcpl;
  assign and_dcpl = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_rdy);
  assign or_dcpl_2 = and_dcpl | (~ ccs_ccore_start_rsci_idat);
  assign this_vld_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_vld <= 1'b0;
    end
    else if ( or_4_cse | this_vld_mx0c1 ) begin
      this_vld <= ~ this_vld_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      m_logical_addr_buf_lpi_1_dfm <= 8'b00000000;
    end
    else if ( ~ or_dcpl_2 ) begin
      m_logical_addr_buf_lpi_1_dfm <= m_logical_addr_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      m_data_data_buf_lpi_1_dfm <= 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ or_dcpl_2 ) begin
      m_data_data_buf_lpi_1_dfm <= m_data_data_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_4_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_spec_StreamType_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module ActUnit_Connections_OutBlocking_spec_StreamType_Connections_SYN_PORT_Push (
  this_vld, this_rdy, this_dat, m_data_data_rsc_dat, m_logical_addr_rsc_dat, ccs_ccore_start_rsc_dat,
      ccs_ccore_done_sync_vld, ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  input this_rdy;
  output [521:0] this_dat;
  input [511:0] m_data_data_rsc_dat;
  input [7:0] m_logical_addr_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  ActUnit_Connections_OutBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_spec_StreamType_Connections_SYN_PORT_Push_core
      Connections_OutBlocking_spec_StreamType_Connections_SYN_PORT_Push_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .m_data_data_rsc_dat(m_data_data_rsc_dat),
      .m_logical_addr_rsc_dat(m_logical_addr_rsc_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./ActUnit_Connections_OutBlockingless_boolcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ActUnit_Connections_OutBlockingless_boolcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./ActUnit_Connections_OutBlockingless_boolcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module ActUnit_Connections_OutBlockingless_boolcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./ActUnit_Connections_OutBlockingless_boolcomma_Connections_SYN_PORTgreater_Push.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   code@iron-06
//  Generated date: Mon Jan 26 19:49:20 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlockingless_boolcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_bool_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module ActUnit_Connections_OutBlockingless_boolcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_bool_Connections_SYN_PORT_Push_core
    (
  this_vld, this_rdy, this_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  reg this_vld;
  input this_rdy;
  output this_dat;
  reg this_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_4_cse;
  wire this_vld_mx0c1;


  // Interconnect Declarations for Component Instantiations
  wire  nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  ActUnit_Connections_OutBlockingless_boolcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd53),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  ActUnit_Connections_OutBlockingless_boolcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1
      #(.rscid(32'sd59)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld)
    );
  assign or_4_cse = ccs_ccore_start_rsci_idat | (io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & (~ this_rdy));
  assign this_vld_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_vld <= 1'b0;
    end
    else if ( or_4_cse | this_vld_mx0c1 ) begin
      this_vld <= ~ this_vld_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_dat <= 1'b0;
    end
    else if ( (~((~ io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1) | this_rdy)) | ccs_ccore_start_rsci_idat
        ) begin
      this_dat <= 1'b1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_4_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_bool_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module ActUnit_Connections_OutBlocking_bool_Connections_SYN_PORT_Push (
  this_vld, this_rdy, this_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  input this_rdy;
  output this_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  ActUnit_Connections_OutBlockingless_boolcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_bool_Connections_SYN_PORT_Push_core
      Connections_OutBlocking_bool_Connections_SYN_PORT_Push_core_inst (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./ActUnit_mgc_mul_pipe_beh.v 
//
// File:      $Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_mul_pipe_beh.v
//
// BASELINE:  Catapult-C version 2006b.63
// MODIFIED:  2007-04-03, tnagler
//
// Note: this file uses Verilog2001 features;
//       please enable Verilog2001 in the flow!

module ActUnit_mgc_mul_pipe (a, b, clk, en, a_rst, s_rst, z);

    // Parameters:
    parameter integer width_a = 32'd4;  // input a bit width
    parameter         signd_a =  1'b1;  // input a type (1=signed, 0=unsigned)
    parameter integer width_b = 32'd4;  // input b bit width
    parameter         signd_b =  1'b1;  // input b type (1=signed, 0=unsigned)
    parameter integer width_z = 32'd8;  // result bit width (= width_a + width_b)
    parameter      clock_edge =  1'b0;  // clock polarity (1=posedge, 0=negedge)
    parameter   enable_active =  1'b0;  // enable polarity (1=posedge, 0=negedge)
    parameter    a_rst_active =  1'b1;  // unused
    parameter    s_rst_active =  1'b1;  // unused
    parameter integer  stages = 32'd2;  // number of output registers + 1 (careful!)
    parameter integer n_inreg = 32'd0;  // number of input registers

    localparam integer width_ab = width_a + width_b;  // multiplier result width
    localparam integer n_inreg_min = (n_inreg > 1) ? (n_inreg-1) : 0; // for Synopsys DC

    // I/O ports:
    input  [width_a-1:0] a;      // input A
    input  [width_b-1:0] b;      // input B
    input                clk;    // clock
    input                en;     // enable
    input                a_rst;  // spyglass disable SYNTH_5121,W240
    input                s_rst;  // spyglass disable SYNTH_5121,W240
    output [width_z-1:0] z;      // output


    // Input registers:

    wire [width_a-1:0] a_f;
    wire [width_b-1:0] b_f;

    integer i;

    generate
    if (clock_edge == 1'b0)
    begin: NEG_EDGE1
        case (n_inreg)
        32'd0: begin: B1
            assign a_f = a,
                   b_f = b;
        end
        default: begin: B2
            reg [width_a-1:0] a_reg [n_inreg_min:0];
            reg [width_b-1:0] b_reg [n_inreg_min:0];
            always @(negedge clk)
            if (en == enable_active)
            begin: B21
                a_reg[0] <= a;
                b_reg[0] <= b;
                for (i = 0; i < n_inreg_min; i = i + 1)
                begin: B3
                    a_reg[i+1] <= a_reg[i]; //spyglass disable FlopEConst
                    b_reg[i+1] <= b_reg[i]; //spyglass disable FlopEConst
                end
            end
            assign a_f = a_reg[n_inreg_min],
                   b_f = b_reg[n_inreg_min];
        end
        endcase
    end
    else
    begin: POS_EDGE1
        case (n_inreg)
        32'd0: begin: B1
            assign a_f = a,
                   b_f = b;
        end
        default: begin: B2
            reg [width_a-1:0] a_reg [n_inreg_min:0];
            reg [width_b-1:0] b_reg [n_inreg_min:0];
            always @(posedge clk)
            if (en == enable_active)
            begin: B21
                a_reg[0] <= a; //spyglass disable FlopEConst
                b_reg[0] <= b; //spyglass disable FlopEConst
                for (i = 0; i < n_inreg_min; i = i + 1)
                begin: B3
                    a_reg[i+1] <= a_reg[i]; //spyglass disable FlopEConst
                    b_reg[i+1] <= b_reg[i]; //spyglass disable FlopEConst
                end
            end
            assign a_f = a_reg[n_inreg_min],
                   b_f = b_reg[n_inreg_min];
        end
        endcase
    end
    endgenerate


    // Output:
    wire [width_z-1:0]  xz;

    function signed [width_z-1:0] conv_signed;
      input signed [width_ab-1:0] res;
      conv_signed = res[width_z-1:0];
    endfunction

    generate
      wire signed [width_ab-1:0] res;
      if ( (signd_a == 1'b1) && (signd_b == 1'b1) )
      begin: SIGNED_AB
              assign res = $signed(a_f) * $signed(b_f);
              assign xz = conv_signed(res);
      end
      else if ( (signd_a == 1'b1) && (signd_b == 1'b0) )
      begin: SIGNED_A
              assign res = $signed(a_f) * $signed({1'b0, b_f});
              assign xz = conv_signed(res);
      end
      else if ( (signd_a == 1'b0) && (signd_b == 1'b1) )
      begin: SIGNED_B
              assign res = $signed({1'b0,a_f}) * $signed(b_f);
              assign xz = conv_signed(res);
      end
      else
      begin: UNSIGNED_AB
              assign res = a_f * b_f;
	      assign xz = res[width_z-1:0];
      end
    endgenerate


    // Output registers:

    reg  [width_z-1:0] reg_array[stages-2:0];
    wire [width_z-1:0] z;

    generate
    if (clock_edge == 1'b0)
    begin: NEG_EDGE2
        always @(negedge clk)
        if (en == enable_active)
            for (i = stages-2; i >= 0; i = i-1)
                if (i == 0)
                    reg_array[i] <= xz; //spyglass disable FlopEConst
                else
                    reg_array[i] <= reg_array[i-1]; //spyglass disable FlopEConst
    end
    else
    begin: POS_EDGE2
        always @(posedge clk)
        if (en == enable_active)
            for (i = stages-2; i >= 0; i = i-1)
                if (i == 0)
                    reg_array[i] <= xz; //spyglass disable FlopEConst
                else
                    reg_array[i] <= reg_array[i-1]; //spyglass disable FlopEConst
    end
    endgenerate

    assign z = reg_array[stages-2];
endmodule

//------> ./ActUnit.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
// 
//  Generated by:   code@iron-06
//  Generated date: Thu Jan 29 12:29:03 2026
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_ActUnitRun_fsm
//  FSM Module
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_ActUnitRun_fsm (
  clk, rst, ActUnitRun_wen, fsm_output, while_C_0_tr0, ActUnit_RunInst_case_2_for_C_0_tr0,
      while_C_11_tr0, ActUnit_PushOutput_if_for_C_0_tr0, while_C_13_tr0, ActUnit_RunLoad_if_else_for_C_0_tr0
);
  input clk;
  input rst;
  input ActUnitRun_wen;
  output [4:0] fsm_output;
  reg [4:0] fsm_output;
  input while_C_0_tr0;
  input ActUnit_RunInst_case_2_for_C_0_tr0;
  input while_C_11_tr0;
  input ActUnit_PushOutput_if_for_C_0_tr0;
  input while_C_13_tr0;
  input ActUnit_RunLoad_if_else_for_C_0_tr0;


  // FSM State Type Declaration for ActUnit_ActUnit_ActUnitRun_ActUnitRun_fsm_1
  parameter
    ActUnitRun_rlp_C_0 = 5'd0,
    while_C_0 = 5'd1,
    ActUnit_RunInst_case_2_for_C_0 = 5'd2,
    while_C_1 = 5'd3,
    while_C_2 = 5'd4,
    while_C_3 = 5'd5,
    while_C_4 = 5'd6,
    while_C_5 = 5'd7,
    while_C_6 = 5'd8,
    while_C_7 = 5'd9,
    while_C_8 = 5'd10,
    while_C_9 = 5'd11,
    while_C_10 = 5'd12,
    while_C_11 = 5'd13,
    ActUnit_PushOutput_if_for_C_0 = 5'd14,
    while_C_12 = 5'd15,
    while_C_13 = 5'd16,
    ActUnit_RunLoad_if_else_for_C_0 = 5'd17,
    while_C_14 = 5'd18,
    while_C_15 = 5'd19;

  reg [4:0] state_var;
  reg [4:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : ActUnit_ActUnit_ActUnitRun_ActUnitRun_fsm_1
    case (state_var)
      while_C_0 : begin
        fsm_output = 5'b00001;
        if ( while_C_0_tr0 ) begin
          state_var_NS = while_C_1;
        end
        else begin
          state_var_NS = ActUnit_RunInst_case_2_for_C_0;
        end
      end
      ActUnit_RunInst_case_2_for_C_0 : begin
        fsm_output = 5'b00010;
        if ( ActUnit_RunInst_case_2_for_C_0_tr0 ) begin
          state_var_NS = while_C_1;
        end
        else begin
          state_var_NS = ActUnit_RunInst_case_2_for_C_0;
        end
      end
      while_C_1 : begin
        fsm_output = 5'b00011;
        state_var_NS = while_C_2;
      end
      while_C_2 : begin
        fsm_output = 5'b00100;
        state_var_NS = while_C_3;
      end
      while_C_3 : begin
        fsm_output = 5'b00101;
        state_var_NS = while_C_4;
      end
      while_C_4 : begin
        fsm_output = 5'b00110;
        state_var_NS = while_C_5;
      end
      while_C_5 : begin
        fsm_output = 5'b00111;
        state_var_NS = while_C_6;
      end
      while_C_6 : begin
        fsm_output = 5'b01000;
        state_var_NS = while_C_7;
      end
      while_C_7 : begin
        fsm_output = 5'b01001;
        state_var_NS = while_C_8;
      end
      while_C_8 : begin
        fsm_output = 5'b01010;
        state_var_NS = while_C_9;
      end
      while_C_9 : begin
        fsm_output = 5'b01011;
        state_var_NS = while_C_10;
      end
      while_C_10 : begin
        fsm_output = 5'b01100;
        state_var_NS = while_C_11;
      end
      while_C_11 : begin
        fsm_output = 5'b01101;
        if ( while_C_11_tr0 ) begin
          state_var_NS = while_C_12;
        end
        else begin
          state_var_NS = ActUnit_PushOutput_if_for_C_0;
        end
      end
      ActUnit_PushOutput_if_for_C_0 : begin
        fsm_output = 5'b01110;
        if ( ActUnit_PushOutput_if_for_C_0_tr0 ) begin
          state_var_NS = while_C_12;
        end
        else begin
          state_var_NS = ActUnit_PushOutput_if_for_C_0;
        end
      end
      while_C_12 : begin
        fsm_output = 5'b01111;
        state_var_NS = while_C_13;
      end
      while_C_13 : begin
        fsm_output = 5'b10000;
        if ( while_C_13_tr0 ) begin
          state_var_NS = while_C_14;
        end
        else begin
          state_var_NS = ActUnit_RunLoad_if_else_for_C_0;
        end
      end
      ActUnit_RunLoad_if_else_for_C_0 : begin
        fsm_output = 5'b10001;
        if ( ActUnit_RunLoad_if_else_for_C_0_tr0 ) begin
          state_var_NS = while_C_14;
        end
        else begin
          state_var_NS = ActUnit_RunLoad_if_else_for_C_0;
        end
      end
      while_C_14 : begin
        fsm_output = 5'b10010;
        state_var_NS = while_C_15;
      end
      while_C_15 : begin
        fsm_output = 5'b10011;
        state_var_NS = while_C_0;
      end
      // ActUnitRun_rlp_C_0
      default : begin
        fsm_output = 5'b00000;
        state_var_NS = while_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      state_var <= ActUnitRun_rlp_C_0;
    end
    else if ( ActUnitRun_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_staller
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_staller (
  clk, rst, ActUnitRun_wen, ActUnitRun_wten, rva_out_Push_mioi_wen_comp, output_port_Push_mioi_wen_comp,
      done_Push_mioi_wen_comp
);
  input clk;
  input rst;
  output ActUnitRun_wen;
  output ActUnitRun_wten;
  input rva_out_Push_mioi_wen_comp;
  input output_port_Push_mioi_wen_comp;
  input done_Push_mioi_wen_comp;


  // Interconnect Declarations
  reg ActUnitRun_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign ActUnitRun_wen = rva_out_Push_mioi_wen_comp & output_port_Push_mioi_wen_comp
      & done_Push_mioi_wen_comp;
  assign ActUnitRun_wten = ActUnitRun_wten_reg;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnitRun_wten_reg <= 1'b0;
    end
    else begin
      ActUnitRun_wten_reg <= ~ ActUnitRun_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_wait_dp
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_wait_dp (
  ActUnitRun_wen, Tanh_for_3_else_else_mul_1_cmp_cgo, Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg,
      Tanh_for_3_else_else_mul_1_cmp_en, Tanh_for_3_else_else_mul_1_cmp_cgo_1, Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_1,
      Tanh_for_3_else_else_mul_1_cmp_1_en, Tanh_for_3_else_else_mul_1_cmp_cgo_2,
      Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_2, Tanh_for_3_else_else_mul_1_cmp_2_en,
      Tanh_for_3_else_else_mul_1_cmp_cgo_3, Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_3,
      Tanh_for_3_else_else_mul_1_cmp_3_en, Tanh_for_3_else_else_mul_1_cmp_cgo_4,
      Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_4, Tanh_for_3_else_else_mul_1_cmp_4_en,
      Tanh_for_3_else_else_mul_1_cmp_cgo_5, Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_5,
      Tanh_for_3_else_else_mul_1_cmp_5_en, Tanh_for_3_else_else_mul_1_cmp_cgo_6,
      Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_6, Tanh_for_3_else_else_mul_1_cmp_6_en,
      Tanh_for_3_else_else_mul_1_cmp_cgo_7, Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_7,
      Tanh_for_3_else_else_mul_1_cmp_7_en, Tanh_for_3_else_else_mul_1_cmp_cgo_8,
      Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_8, Tanh_for_3_else_else_mul_1_cmp_8_en,
      Tanh_for_3_else_else_mul_1_cmp_cgo_9, Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_9,
      Tanh_for_3_else_else_mul_1_cmp_9_en, Tanh_for_3_else_else_mul_1_cmp_cgo_10,
      Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_10, Tanh_for_3_else_else_mul_1_cmp_10_en,
      Tanh_for_3_else_else_mul_1_cmp_cgo_11, Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_11,
      Tanh_for_3_else_else_mul_1_cmp_11_en, Tanh_for_3_else_else_mul_1_cmp_cgo_12,
      Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_12, Tanh_for_3_else_else_mul_1_cmp_12_en,
      Tanh_for_3_else_else_mul_1_cmp_cgo_13, Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_13,
      Tanh_for_3_else_else_mul_1_cmp_13_en, Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo,
      Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg, Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_en,
      Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_1, Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_1,
      Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_1_en, Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_2,
      Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_2, Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_2_en,
      Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_3, Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_3,
      Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_3_en, Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_4,
      Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_4, Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_4_en,
      Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_5, Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_5,
      Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_5_en, Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_6,
      Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_6, Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_6_en,
      Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_7, Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_7,
      Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_7_en, Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_8,
      Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_8, Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_8_en,
      Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_9, Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_9,
      Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_9_en, Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_10,
      Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_10, Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_10_en,
      Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_11, Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_11,
      Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_11_en, Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_12,
      Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_12, Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_12_en,
      Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_13, Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_13,
      Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_13_en, Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_14,
      Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_14, Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_14_en,
      Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_15, Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_15,
      Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_15_en, Tanh_for_1_else_else_mul_cmp_cgo,
      Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg, Tanh_for_1_else_else_mul_cmp_en,
      Tanh_for_1_else_else_mul_cmp_cgo_1, Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_1,
      Tanh_for_1_else_else_mul_cmp_1_en, Tanh_for_1_else_else_mul_cmp_cgo_2, Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_2,
      Tanh_for_1_else_else_mul_cmp_2_en, Tanh_for_1_else_else_mul_cmp_cgo_3, Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_3,
      Tanh_for_1_else_else_mul_cmp_3_en, Tanh_for_1_else_else_mul_cmp_cgo_4, Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_4,
      Tanh_for_1_else_else_mul_cmp_4_en, Tanh_for_1_else_else_mul_cmp_cgo_5, Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_5,
      Tanh_for_1_else_else_mul_cmp_5_en, Tanh_for_1_else_else_mul_cmp_cgo_6, Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_6,
      Tanh_for_1_else_else_mul_cmp_6_en, Tanh_for_1_else_else_mul_cmp_cgo_7, Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_7,
      Tanh_for_1_else_else_mul_cmp_7_en, Tanh_for_1_else_else_mul_cmp_cgo_8, Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_8,
      Tanh_for_1_else_else_mul_cmp_8_en, Tanh_for_1_else_else_mul_cmp_cgo_9, Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_9,
      Tanh_for_1_else_else_mul_cmp_9_en, Tanh_for_1_else_else_mul_cmp_cgo_10, Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_10,
      Tanh_for_1_else_else_mul_cmp_10_en, Tanh_for_1_else_else_mul_cmp_cgo_11, Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_11,
      Tanh_for_1_else_else_mul_cmp_11_en, Tanh_for_1_else_else_mul_cmp_cgo_12, Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_12,
      Tanh_for_1_else_else_mul_cmp_12_en, Tanh_for_1_else_else_mul_cmp_cgo_13, Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_13,
      Tanh_for_1_else_else_mul_cmp_13_en, Tanh_for_1_else_else_mul_cmp_cgo_14, Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_14,
      Tanh_for_1_else_else_mul_cmp_14_en, Tanh_for_1_else_else_mul_cmp_cgo_15, Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_15,
      Tanh_for_1_else_else_mul_cmp_15_en, Tanh_for_1_else_else_mul_1_cmp_cgo, Tanh_for_1_else_else_mul_1_cmp_cgo_ir_unreg,
      Tanh_for_1_else_else_mul_1_cmp_en, Tanh_for_1_else_else_mul_1_cmp_cgo_1, Tanh_for_1_else_else_mul_1_cmp_cgo_ir_unreg_1,
      Tanh_for_1_else_else_mul_1_cmp_1_en
);
  input ActUnitRun_wen;
  input Tanh_for_3_else_else_mul_1_cmp_cgo;
  input Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg;
  output Tanh_for_3_else_else_mul_1_cmp_en;
  input Tanh_for_3_else_else_mul_1_cmp_cgo_1;
  input Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_1;
  output Tanh_for_3_else_else_mul_1_cmp_1_en;
  input Tanh_for_3_else_else_mul_1_cmp_cgo_2;
  input Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_2;
  output Tanh_for_3_else_else_mul_1_cmp_2_en;
  input Tanh_for_3_else_else_mul_1_cmp_cgo_3;
  input Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_3;
  output Tanh_for_3_else_else_mul_1_cmp_3_en;
  input Tanh_for_3_else_else_mul_1_cmp_cgo_4;
  input Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_4;
  output Tanh_for_3_else_else_mul_1_cmp_4_en;
  input Tanh_for_3_else_else_mul_1_cmp_cgo_5;
  input Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_5;
  output Tanh_for_3_else_else_mul_1_cmp_5_en;
  input Tanh_for_3_else_else_mul_1_cmp_cgo_6;
  input Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_6;
  output Tanh_for_3_else_else_mul_1_cmp_6_en;
  input Tanh_for_3_else_else_mul_1_cmp_cgo_7;
  input Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_7;
  output Tanh_for_3_else_else_mul_1_cmp_7_en;
  input Tanh_for_3_else_else_mul_1_cmp_cgo_8;
  input Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_8;
  output Tanh_for_3_else_else_mul_1_cmp_8_en;
  input Tanh_for_3_else_else_mul_1_cmp_cgo_9;
  input Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_9;
  output Tanh_for_3_else_else_mul_1_cmp_9_en;
  input Tanh_for_3_else_else_mul_1_cmp_cgo_10;
  input Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_10;
  output Tanh_for_3_else_else_mul_1_cmp_10_en;
  input Tanh_for_3_else_else_mul_1_cmp_cgo_11;
  input Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_11;
  output Tanh_for_3_else_else_mul_1_cmp_11_en;
  input Tanh_for_3_else_else_mul_1_cmp_cgo_12;
  input Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_12;
  output Tanh_for_3_else_else_mul_1_cmp_12_en;
  input Tanh_for_3_else_else_mul_1_cmp_cgo_13;
  input Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_13;
  output Tanh_for_3_else_else_mul_1_cmp_13_en;
  input Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo;
  input Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg;
  output Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_en;
  input Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_1;
  input Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_1;
  output Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_1_en;
  input Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_2;
  input Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_2;
  output Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_2_en;
  input Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_3;
  input Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_3;
  output Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_3_en;
  input Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_4;
  input Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_4;
  output Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_4_en;
  input Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_5;
  input Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_5;
  output Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_5_en;
  input Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_6;
  input Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_6;
  output Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_6_en;
  input Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_7;
  input Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_7;
  output Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_7_en;
  input Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_8;
  input Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_8;
  output Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_8_en;
  input Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_9;
  input Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_9;
  output Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_9_en;
  input Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_10;
  input Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_10;
  output Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_10_en;
  input Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_11;
  input Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_11;
  output Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_11_en;
  input Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_12;
  input Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_12;
  output Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_12_en;
  input Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_13;
  input Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_13;
  output Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_13_en;
  input Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_14;
  input Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_14;
  output Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_14_en;
  input Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_15;
  input Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_15;
  output Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_15_en;
  input Tanh_for_1_else_else_mul_cmp_cgo;
  input Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg;
  output Tanh_for_1_else_else_mul_cmp_en;
  input Tanh_for_1_else_else_mul_cmp_cgo_1;
  input Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_1;
  output Tanh_for_1_else_else_mul_cmp_1_en;
  input Tanh_for_1_else_else_mul_cmp_cgo_2;
  input Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_2;
  output Tanh_for_1_else_else_mul_cmp_2_en;
  input Tanh_for_1_else_else_mul_cmp_cgo_3;
  input Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_3;
  output Tanh_for_1_else_else_mul_cmp_3_en;
  input Tanh_for_1_else_else_mul_cmp_cgo_4;
  input Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_4;
  output Tanh_for_1_else_else_mul_cmp_4_en;
  input Tanh_for_1_else_else_mul_cmp_cgo_5;
  input Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_5;
  output Tanh_for_1_else_else_mul_cmp_5_en;
  input Tanh_for_1_else_else_mul_cmp_cgo_6;
  input Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_6;
  output Tanh_for_1_else_else_mul_cmp_6_en;
  input Tanh_for_1_else_else_mul_cmp_cgo_7;
  input Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_7;
  output Tanh_for_1_else_else_mul_cmp_7_en;
  input Tanh_for_1_else_else_mul_cmp_cgo_8;
  input Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_8;
  output Tanh_for_1_else_else_mul_cmp_8_en;
  input Tanh_for_1_else_else_mul_cmp_cgo_9;
  input Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_9;
  output Tanh_for_1_else_else_mul_cmp_9_en;
  input Tanh_for_1_else_else_mul_cmp_cgo_10;
  input Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_10;
  output Tanh_for_1_else_else_mul_cmp_10_en;
  input Tanh_for_1_else_else_mul_cmp_cgo_11;
  input Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_11;
  output Tanh_for_1_else_else_mul_cmp_11_en;
  input Tanh_for_1_else_else_mul_cmp_cgo_12;
  input Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_12;
  output Tanh_for_1_else_else_mul_cmp_12_en;
  input Tanh_for_1_else_else_mul_cmp_cgo_13;
  input Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_13;
  output Tanh_for_1_else_else_mul_cmp_13_en;
  input Tanh_for_1_else_else_mul_cmp_cgo_14;
  input Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_14;
  output Tanh_for_1_else_else_mul_cmp_14_en;
  input Tanh_for_1_else_else_mul_cmp_cgo_15;
  input Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_15;
  output Tanh_for_1_else_else_mul_cmp_15_en;
  input Tanh_for_1_else_else_mul_1_cmp_cgo;
  input Tanh_for_1_else_else_mul_1_cmp_cgo_ir_unreg;
  output Tanh_for_1_else_else_mul_1_cmp_en;
  input Tanh_for_1_else_else_mul_1_cmp_cgo_1;
  input Tanh_for_1_else_else_mul_1_cmp_cgo_ir_unreg_1;
  output Tanh_for_1_else_else_mul_1_cmp_1_en;



  // Interconnect Declarations for Component Instantiations 
  assign Tanh_for_3_else_else_mul_1_cmp_en = ActUnitRun_wen & (Tanh_for_3_else_else_mul_1_cmp_cgo
      | Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg);
  assign Tanh_for_3_else_else_mul_1_cmp_1_en = ActUnitRun_wen & (Tanh_for_3_else_else_mul_1_cmp_cgo_1
      | Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_1);
  assign Tanh_for_3_else_else_mul_1_cmp_2_en = ActUnitRun_wen & (Tanh_for_3_else_else_mul_1_cmp_cgo_2
      | Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_2);
  assign Tanh_for_3_else_else_mul_1_cmp_3_en = ActUnitRun_wen & (Tanh_for_3_else_else_mul_1_cmp_cgo_3
      | Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_3);
  assign Tanh_for_3_else_else_mul_1_cmp_4_en = ActUnitRun_wen & (Tanh_for_3_else_else_mul_1_cmp_cgo_4
      | Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_4);
  assign Tanh_for_3_else_else_mul_1_cmp_5_en = ActUnitRun_wen & (Tanh_for_3_else_else_mul_1_cmp_cgo_5
      | Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_5);
  assign Tanh_for_3_else_else_mul_1_cmp_6_en = ActUnitRun_wen & (Tanh_for_3_else_else_mul_1_cmp_cgo_6
      | Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_6);
  assign Tanh_for_3_else_else_mul_1_cmp_7_en = ActUnitRun_wen & (Tanh_for_3_else_else_mul_1_cmp_cgo_7
      | Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_7);
  assign Tanh_for_3_else_else_mul_1_cmp_8_en = ActUnitRun_wen & (Tanh_for_3_else_else_mul_1_cmp_cgo_8
      | Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_8);
  assign Tanh_for_3_else_else_mul_1_cmp_9_en = ActUnitRun_wen & (Tanh_for_3_else_else_mul_1_cmp_cgo_9
      | Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_9);
  assign Tanh_for_3_else_else_mul_1_cmp_10_en = ActUnitRun_wen & (Tanh_for_3_else_else_mul_1_cmp_cgo_10
      | Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_10);
  assign Tanh_for_3_else_else_mul_1_cmp_11_en = ActUnitRun_wen & (Tanh_for_3_else_else_mul_1_cmp_cgo_11
      | Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_11);
  assign Tanh_for_3_else_else_mul_1_cmp_12_en = ActUnitRun_wen & (Tanh_for_3_else_else_mul_1_cmp_cgo_12
      | Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_12);
  assign Tanh_for_3_else_else_mul_1_cmp_13_en = ActUnitRun_wen & (Tanh_for_3_else_else_mul_1_cmp_cgo_13
      | Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_13);
  assign Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_en = ActUnitRun_wen & (Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo
      | Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg);
  assign Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_1_en = ActUnitRun_wen &
      (Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_1 | Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_1);
  assign Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_2_en = ActUnitRun_wen &
      (Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_2 | Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_2);
  assign Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_3_en = ActUnitRun_wen &
      (Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_3 | Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_3);
  assign Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_4_en = ActUnitRun_wen &
      (Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_4 | Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_4);
  assign Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_5_en = ActUnitRun_wen &
      (Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_5 | Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_5);
  assign Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_6_en = ActUnitRun_wen &
      (Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_6 | Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_6);
  assign Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_7_en = ActUnitRun_wen &
      (Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_7 | Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_7);
  assign Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_8_en = ActUnitRun_wen &
      (Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_8 | Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_8);
  assign Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_9_en = ActUnitRun_wen &
      (Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_9 | Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_9);
  assign Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_10_en = ActUnitRun_wen &
      (Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_10 | Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_10);
  assign Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_11_en = ActUnitRun_wen &
      (Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_11 | Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_11);
  assign Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_12_en = ActUnitRun_wen &
      (Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_12 | Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_12);
  assign Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_13_en = ActUnitRun_wen &
      (Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_13 | Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_13);
  assign Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_14_en = ActUnitRun_wen &
      (Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_14 | Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_14);
  assign Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_15_en = ActUnitRun_wen &
      (Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_15 | Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_15);
  assign Tanh_for_1_else_else_mul_cmp_en = ActUnitRun_wen & (Tanh_for_1_else_else_mul_cmp_cgo
      | Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg);
  assign Tanh_for_1_else_else_mul_cmp_1_en = ActUnitRun_wen & (Tanh_for_1_else_else_mul_cmp_cgo_1
      | Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_1);
  assign Tanh_for_1_else_else_mul_cmp_2_en = ActUnitRun_wen & (Tanh_for_1_else_else_mul_cmp_cgo_2
      | Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_2);
  assign Tanh_for_1_else_else_mul_cmp_3_en = ActUnitRun_wen & (Tanh_for_1_else_else_mul_cmp_cgo_3
      | Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_3);
  assign Tanh_for_1_else_else_mul_cmp_4_en = ActUnitRun_wen & (Tanh_for_1_else_else_mul_cmp_cgo_4
      | Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_4);
  assign Tanh_for_1_else_else_mul_cmp_5_en = ActUnitRun_wen & (Tanh_for_1_else_else_mul_cmp_cgo_5
      | Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_5);
  assign Tanh_for_1_else_else_mul_cmp_6_en = ActUnitRun_wen & (Tanh_for_1_else_else_mul_cmp_cgo_6
      | Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_6);
  assign Tanh_for_1_else_else_mul_cmp_7_en = ActUnitRun_wen & (Tanh_for_1_else_else_mul_cmp_cgo_7
      | Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_7);
  assign Tanh_for_1_else_else_mul_cmp_8_en = ActUnitRun_wen & (Tanh_for_1_else_else_mul_cmp_cgo_8
      | Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_8);
  assign Tanh_for_1_else_else_mul_cmp_9_en = ActUnitRun_wen & (Tanh_for_1_else_else_mul_cmp_cgo_9
      | Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_9);
  assign Tanh_for_1_else_else_mul_cmp_10_en = ActUnitRun_wen & (Tanh_for_1_else_else_mul_cmp_cgo_10
      | Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_10);
  assign Tanh_for_1_else_else_mul_cmp_11_en = ActUnitRun_wen & (Tanh_for_1_else_else_mul_cmp_cgo_11
      | Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_11);
  assign Tanh_for_1_else_else_mul_cmp_12_en = ActUnitRun_wen & (Tanh_for_1_else_else_mul_cmp_cgo_12
      | Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_12);
  assign Tanh_for_1_else_else_mul_cmp_13_en = ActUnitRun_wen & (Tanh_for_1_else_else_mul_cmp_cgo_13
      | Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_13);
  assign Tanh_for_1_else_else_mul_cmp_14_en = ActUnitRun_wen & (Tanh_for_1_else_else_mul_cmp_cgo_14
      | Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_14);
  assign Tanh_for_1_else_else_mul_cmp_15_en = ActUnitRun_wen & (Tanh_for_1_else_else_mul_cmp_cgo_15
      | Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_15);
  assign Tanh_for_1_else_else_mul_1_cmp_en = ActUnitRun_wen & (Tanh_for_1_else_else_mul_1_cmp_cgo
      | Tanh_for_1_else_else_mul_1_cmp_cgo_ir_unreg);
  assign Tanh_for_1_else_else_mul_1_cmp_1_en = ActUnitRun_wen & (Tanh_for_1_else_else_mul_1_cmp_cgo_1
      | Tanh_for_1_else_else_mul_1_cmp_cgo_ir_unreg_1);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_done_Push_mioi_done_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_done_Push_mioi_done_Push_mio_wait_ctrl (
  ActUnitRun_wten, done_Push_mioi_iswt0, done_Push_mioi_biwt, done_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct,
      done_Push_mioi_ccs_ccore_done_sync_vld, done_Push_mioi_iswt0_pff
);
  input ActUnitRun_wten;
  input done_Push_mioi_iswt0;
  output done_Push_mioi_biwt;
  output done_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct;
  input done_Push_mioi_ccs_ccore_done_sync_vld;
  input done_Push_mioi_iswt0_pff;



  // Interconnect Declarations for Component Instantiations 
  assign done_Push_mioi_biwt = done_Push_mioi_iswt0 & done_Push_mioi_ccs_ccore_done_sync_vld;
  assign done_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct = (~ ActUnitRun_wten)
      & done_Push_mioi_iswt0_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_output_port_Push_mioi_output_port_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_output_port_Push_mioi_output_port_Push_mio_wait_ctrl
    (
  ActUnitRun_wten, output_port_Push_mioi_iswt0, output_port_Push_mioi_biwt, output_port_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct,
      output_port_Push_mioi_ccs_ccore_done_sync_vld, output_port_Push_mioi_iswt0_pff
);
  input ActUnitRun_wten;
  input output_port_Push_mioi_iswt0;
  output output_port_Push_mioi_biwt;
  output output_port_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct;
  input output_port_Push_mioi_ccs_ccore_done_sync_vld;
  input output_port_Push_mioi_iswt0_pff;



  // Interconnect Declarations for Component Instantiations 
  assign output_port_Push_mioi_biwt = output_port_Push_mioi_iswt0 & output_port_Push_mioi_ccs_ccore_done_sync_vld;
  assign output_port_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct = (~ ActUnitRun_wten)
      & output_port_Push_mioi_iswt0_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_start_PopNB_mioi_start_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_start_PopNB_mioi_start_PopNB_mio_wait_dp (
  clk, rst, start_PopNB_mioi_data_rsc_z_mxwt, start_PopNB_mioi_return_rsc_z_mxwt,
      start_PopNB_mioi_biwt, start_PopNB_mioi_bdwt, start_PopNB_mioi_data_rsc_z,
      start_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output start_PopNB_mioi_data_rsc_z_mxwt;
  output start_PopNB_mioi_return_rsc_z_mxwt;
  input start_PopNB_mioi_biwt;
  input start_PopNB_mioi_bdwt;
  input start_PopNB_mioi_data_rsc_z;
  input start_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg start_PopNB_mioi_bcwt;
  reg start_PopNB_mioi_data_rsc_z_bfwt;
  reg start_PopNB_mioi_return_rsc_z_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign start_PopNB_mioi_data_rsc_z_mxwt = MUX_s_1_2_2(start_PopNB_mioi_data_rsc_z,
      start_PopNB_mioi_data_rsc_z_bfwt, start_PopNB_mioi_bcwt);
  assign start_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(start_PopNB_mioi_return_rsc_z,
      start_PopNB_mioi_return_rsc_z_bfwt, start_PopNB_mioi_bcwt);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      start_PopNB_mioi_bcwt <= 1'b0;
    end
    else begin
      start_PopNB_mioi_bcwt <= ~((~(start_PopNB_mioi_bcwt | start_PopNB_mioi_biwt))
          | start_PopNB_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      start_PopNB_mioi_data_rsc_z_bfwt <= 1'b0;
      start_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else if ( start_PopNB_mioi_biwt ) begin
      start_PopNB_mioi_data_rsc_z_bfwt <= start_PopNB_mioi_data_rsc_z;
      start_PopNB_mioi_return_rsc_z_bfwt <= start_PopNB_mioi_return_rsc_z;
    end
  end

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_start_PopNB_mioi_start_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_start_PopNB_mioi_start_PopNB_mio_wait_ctrl (
  ActUnitRun_wen, ActUnitRun_wten, start_PopNB_mioi_oswt, start_PopNB_mioi_biwt,
      start_PopNB_mioi_bdwt, start_PopNB_mioi_biwt_pff, start_PopNB_mioi_oswt_pff
);
  input ActUnitRun_wen;
  input ActUnitRun_wten;
  input start_PopNB_mioi_oswt;
  output start_PopNB_mioi_biwt;
  output start_PopNB_mioi_bdwt;
  output start_PopNB_mioi_biwt_pff;
  input start_PopNB_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign start_PopNB_mioi_bdwt = start_PopNB_mioi_oswt & ActUnitRun_wen;
  assign start_PopNB_mioi_biwt = (~ ActUnitRun_wten) & start_PopNB_mioi_oswt;
  assign start_PopNB_mioi_biwt_pff = ActUnitRun_wen & start_PopNB_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl (
  ActUnitRun_wten, rva_out_Push_mioi_iswt0, rva_out_Push_mioi_biwt, rva_out_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct,
      rva_out_Push_mioi_ccs_ccore_done_sync_vld, rva_out_Push_mioi_iswt0_pff
);
  input ActUnitRun_wten;
  input rva_out_Push_mioi_iswt0;
  output rva_out_Push_mioi_biwt;
  output rva_out_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct;
  input rva_out_Push_mioi_ccs_ccore_done_sync_vld;
  input rva_out_Push_mioi_iswt0_pff;



  // Interconnect Declarations for Component Instantiations 
  assign rva_out_Push_mioi_biwt = rva_out_Push_mioi_iswt0 & rva_out_Push_mioi_ccs_ccore_done_sync_vld;
  assign rva_out_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct = (~ ActUnitRun_wten)
      & rva_out_Push_mioi_iswt0_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_act_port_PopNB_mioi_act_port_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_act_port_PopNB_mioi_act_port_PopNB_mio_wait_dp
    (
  clk, rst, act_port_PopNB_mioi_data_data_rsc_z_mxwt, act_port_PopNB_mioi_return_rsc_z_mxwt,
      act_port_PopNB_mioi_biwt, act_port_PopNB_mioi_bdwt, act_port_PopNB_mioi_data_data_rsc_z,
      act_port_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output [511:0] act_port_PopNB_mioi_data_data_rsc_z_mxwt;
  output act_port_PopNB_mioi_return_rsc_z_mxwt;
  input act_port_PopNB_mioi_biwt;
  input act_port_PopNB_mioi_bdwt;
  input [511:0] act_port_PopNB_mioi_data_data_rsc_z;
  input act_port_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg act_port_PopNB_mioi_bcwt;
  reg [511:0] act_port_PopNB_mioi_data_data_rsc_z_bfwt;
  reg act_port_PopNB_mioi_return_rsc_z_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign act_port_PopNB_mioi_data_data_rsc_z_mxwt = MUX_v_512_2_2(act_port_PopNB_mioi_data_data_rsc_z,
      act_port_PopNB_mioi_data_data_rsc_z_bfwt, act_port_PopNB_mioi_bcwt);
  assign act_port_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(act_port_PopNB_mioi_return_rsc_z,
      act_port_PopNB_mioi_return_rsc_z_bfwt, act_port_PopNB_mioi_bcwt);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_PopNB_mioi_bcwt <= 1'b0;
    end
    else begin
      act_port_PopNB_mioi_bcwt <= ~((~(act_port_PopNB_mioi_bcwt | act_port_PopNB_mioi_biwt))
          | act_port_PopNB_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_PopNB_mioi_data_data_rsc_z_bfwt <= 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      act_port_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else if ( act_port_PopNB_mioi_biwt ) begin
      act_port_PopNB_mioi_data_data_rsc_z_bfwt <= act_port_PopNB_mioi_data_data_rsc_z;
      act_port_PopNB_mioi_return_rsc_z_bfwt <= act_port_PopNB_mioi_return_rsc_z;
    end
  end

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [511:0] MUX_v_512_2_2;
    input [511:0] input_0;
    input [511:0] input_1;
    input  sel;
    reg [511:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_512_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_act_port_PopNB_mioi_act_port_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_act_port_PopNB_mioi_act_port_PopNB_mio_wait_ctrl
    (
  ActUnitRun_wen, ActUnitRun_wten, act_port_PopNB_mioi_oswt, act_port_PopNB_mioi_biwt,
      act_port_PopNB_mioi_bdwt, act_port_PopNB_mioi_biwt_pff, act_port_PopNB_mioi_oswt_pff
);
  input ActUnitRun_wen;
  input ActUnitRun_wten;
  input act_port_PopNB_mioi_oswt;
  output act_port_PopNB_mioi_biwt;
  output act_port_PopNB_mioi_bdwt;
  output act_port_PopNB_mioi_biwt_pff;
  input act_port_PopNB_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign act_port_PopNB_mioi_bdwt = act_port_PopNB_mioi_oswt & ActUnitRun_wen;
  assign act_port_PopNB_mioi_biwt = (~ ActUnitRun_wten) & act_port_PopNB_mioi_oswt;
  assign act_port_PopNB_mioi_biwt_pff = ActUnitRun_wen & act_port_PopNB_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp (
  clk, rst, rva_in_PopNB_mioi_data_data_rsc_z_mxwt, rva_in_PopNB_mioi_data_addr_rsc_z_mxwt,
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt, rva_in_PopNB_mioi_return_rsc_z_mxwt,
      rva_in_PopNB_mioi_biwt, rva_in_PopNB_mioi_bdwt, rva_in_PopNB_mioi_data_data_rsc_z,
      rva_in_PopNB_mioi_data_addr_rsc_z, rva_in_PopNB_mioi_data_rw_rsc_z, rva_in_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output [511:0] rva_in_PopNB_mioi_data_data_rsc_z_mxwt;
  output [11:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt;
  output rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  output rva_in_PopNB_mioi_return_rsc_z_mxwt;
  input rva_in_PopNB_mioi_biwt;
  input rva_in_PopNB_mioi_bdwt;
  input [511:0] rva_in_PopNB_mioi_data_data_rsc_z;
  input [23:0] rva_in_PopNB_mioi_data_addr_rsc_z;
  input rva_in_PopNB_mioi_data_rw_rsc_z;
  input rva_in_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg rva_in_PopNB_mioi_bcwt;
  reg [511:0] rva_in_PopNB_mioi_data_data_rsc_z_bfwt;
  reg rva_in_PopNB_mioi_data_rw_rsc_z_bfwt;
  reg rva_in_PopNB_mioi_return_rsc_z_bfwt;
  reg [3:0] rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_23_20;
  reg [7:0] rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_11_4;

  wire[3:0] ActUnit_DecodeAxi_if_mux_3_nl;
  wire[7:0] ActUnit_DecodeAxi_if_mux_9_nl;

  // Interconnect Declarations for Component Instantiations 
  assign rva_in_PopNB_mioi_data_data_rsc_z_mxwt = MUX_v_512_2_2(rva_in_PopNB_mioi_data_data_rsc_z,
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt, rva_in_PopNB_mioi_bcwt);
  assign rva_in_PopNB_mioi_data_rw_rsc_z_mxwt = MUX_s_1_2_2(rva_in_PopNB_mioi_data_rw_rsc_z,
      rva_in_PopNB_mioi_data_rw_rsc_z_bfwt, rva_in_PopNB_mioi_bcwt);
  assign rva_in_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(rva_in_PopNB_mioi_return_rsc_z,
      rva_in_PopNB_mioi_return_rsc_z_bfwt, rva_in_PopNB_mioi_bcwt);
  assign ActUnit_DecodeAxi_if_mux_3_nl = MUX_v_4_2_2((rva_in_PopNB_mioi_data_addr_rsc_z[23:20]),
      rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_23_20, rva_in_PopNB_mioi_bcwt);
  assign ActUnit_DecodeAxi_if_mux_9_nl = MUX_v_8_2_2((rva_in_PopNB_mioi_data_addr_rsc_z[11:4]),
      rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_11_4, rva_in_PopNB_mioi_bcwt);
  assign rva_in_PopNB_mioi_data_addr_rsc_z_mxwt = {ActUnit_DecodeAxi_if_mux_3_nl
      , ActUnit_DecodeAxi_if_mux_9_nl};
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_PopNB_mioi_bcwt <= 1'b0;
    end
    else begin
      rva_in_PopNB_mioi_bcwt <= ~((~(rva_in_PopNB_mioi_bcwt | rva_in_PopNB_mioi_biwt))
          | rva_in_PopNB_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt <= 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_23_20 <= 4'b0000;
      rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_11_4 <= 8'b00000000;
      rva_in_PopNB_mioi_data_rw_rsc_z_bfwt <= 1'b0;
      rva_in_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else if ( rva_in_PopNB_mioi_biwt ) begin
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt <= rva_in_PopNB_mioi_data_data_rsc_z;
      rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_23_20 <= rva_in_PopNB_mioi_data_addr_rsc_z[23:20];
      rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_11_4 <= rva_in_PopNB_mioi_data_addr_rsc_z[11:4];
      rva_in_PopNB_mioi_data_rw_rsc_z_bfwt <= rva_in_PopNB_mioi_data_rw_rsc_z;
      rva_in_PopNB_mioi_return_rsc_z_bfwt <= rva_in_PopNB_mioi_return_rsc_z;
    end
  end

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input  sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [511:0] MUX_v_512_2_2;
    input [511:0] input_0;
    input [511:0] input_1;
    input  sel;
    reg [511:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_512_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl (
  ActUnitRun_wen, ActUnitRun_wten, rva_in_PopNB_mioi_oswt, rva_in_PopNB_mioi_biwt,
      rva_in_PopNB_mioi_bdwt, rva_in_PopNB_mioi_biwt_pff, rva_in_PopNB_mioi_oswt_pff
);
  input ActUnitRun_wen;
  input ActUnitRun_wten;
  input rva_in_PopNB_mioi_oswt;
  output rva_in_PopNB_mioi_biwt;
  output rva_in_PopNB_mioi_bdwt;
  output rva_in_PopNB_mioi_biwt_pff;
  input rva_in_PopNB_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign rva_in_PopNB_mioi_bdwt = rva_in_PopNB_mioi_oswt & ActUnitRun_wen;
  assign rva_in_PopNB_mioi_biwt = (~ ActUnitRun_wten) & rva_in_PopNB_mioi_oswt;
  assign rva_in_PopNB_mioi_biwt_pff = ActUnitRun_wen & rva_in_PopNB_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_done_Push_mioi
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_done_Push_mioi (
  clk, rst, done_vld, done_rdy, done_dat, ActUnitRun_wten, done_Push_mioi_oswt, done_Push_mioi_wen_comp,
      done_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output done_vld;
  input done_rdy;
  output done_dat;
  input ActUnitRun_wten;
  input done_Push_mioi_oswt;
  output done_Push_mioi_wen_comp;
  input done_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire done_Push_mioi_biwt;
  wire done_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct;
  wire done_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  ActUnit_Connections_OutBlocking_bool_Connections_SYN_PORT_Push  done_Push_mioi
      (
      .this_vld(done_vld),
      .this_rdy(done_rdy),
      .this_dat(done_dat),
      .ccs_ccore_start_rsc_dat(done_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct),
      .ccs_ccore_done_sync_vld(done_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  ActUnit_ActUnit_ActUnitRun_done_Push_mioi_done_Push_mio_wait_ctrl ActUnit_ActUnitRun_done_Push_mioi_done_Push_mio_wait_ctrl_inst
      (
      .ActUnitRun_wten(ActUnitRun_wten),
      .done_Push_mioi_iswt0(done_Push_mioi_oswt),
      .done_Push_mioi_biwt(done_Push_mioi_biwt),
      .done_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct(done_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct),
      .done_Push_mioi_ccs_ccore_done_sync_vld(done_Push_mioi_ccs_ccore_done_sync_vld),
      .done_Push_mioi_iswt0_pff(done_Push_mioi_oswt_pff)
    );
  assign done_Push_mioi_wen_comp = (~ done_Push_mioi_oswt) | done_Push_mioi_biwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_output_port_Push_mioi
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_output_port_Push_mioi (
  clk, rst, output_port_vld, output_port_rdy, output_port_dat, ActUnitRun_wten, output_port_Push_mioi_oswt,
      output_port_Push_mioi_wen_comp, output_port_Push_mioi_m_data_data_rsc_dat_ActUnitRun,
      output_port_Push_mioi_m_logical_addr_rsc_dat_ActUnitRun, output_port_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output output_port_vld;
  input output_port_rdy;
  output [521:0] output_port_dat;
  input ActUnitRun_wten;
  input output_port_Push_mioi_oswt;
  output output_port_Push_mioi_wen_comp;
  input [511:0] output_port_Push_mioi_m_data_data_rsc_dat_ActUnitRun;
  input [7:0] output_port_Push_mioi_m_logical_addr_rsc_dat_ActUnitRun;
  input output_port_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire output_port_Push_mioi_biwt;
  wire output_port_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct;
  wire output_port_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  ActUnit_Connections_OutBlocking_spec_StreamType_Connections_SYN_PORT_Push  output_port_Push_mioi
      (
      .this_vld(output_port_vld),
      .this_rdy(output_port_rdy),
      .this_dat(output_port_dat),
      .m_data_data_rsc_dat(output_port_Push_mioi_m_data_data_rsc_dat_ActUnitRun),
      .m_logical_addr_rsc_dat(output_port_Push_mioi_m_logical_addr_rsc_dat_ActUnitRun),
      .ccs_ccore_start_rsc_dat(output_port_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct),
      .ccs_ccore_done_sync_vld(output_port_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  ActUnit_ActUnit_ActUnitRun_output_port_Push_mioi_output_port_Push_mio_wait_ctrl
      ActUnit_ActUnitRun_output_port_Push_mioi_output_port_Push_mio_wait_ctrl_inst
      (
      .ActUnitRun_wten(ActUnitRun_wten),
      .output_port_Push_mioi_iswt0(output_port_Push_mioi_oswt),
      .output_port_Push_mioi_biwt(output_port_Push_mioi_biwt),
      .output_port_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct(output_port_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct),
      .output_port_Push_mioi_ccs_ccore_done_sync_vld(output_port_Push_mioi_ccs_ccore_done_sync_vld),
      .output_port_Push_mioi_iswt0_pff(output_port_Push_mioi_oswt_pff)
    );
  assign output_port_Push_mioi_wen_comp = (~ output_port_Push_mioi_oswt) | output_port_Push_mioi_biwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_start_PopNB_mioi
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_start_PopNB_mioi (
  clk, rst, start_vld, start_rdy, start_dat, ActUnitRun_wen, ActUnitRun_wten, start_PopNB_mioi_oswt,
      start_PopNB_mioi_data_rsc_z_mxwt, start_PopNB_mioi_return_rsc_z_mxwt, start_PopNB_mioi_oswt_pff
);
  input clk;
  input rst;
  input start_vld;
  output start_rdy;
  input start_dat;
  input ActUnitRun_wen;
  input ActUnitRun_wten;
  input start_PopNB_mioi_oswt;
  output start_PopNB_mioi_data_rsc_z_mxwt;
  output start_PopNB_mioi_return_rsc_z_mxwt;
  input start_PopNB_mioi_oswt_pff;


  // Interconnect Declarations
  wire start_PopNB_mioi_biwt;
  wire start_PopNB_mioi_bdwt;
  wire start_PopNB_mioi_data_rsc_z;
  wire start_PopNB_mioi_return_rsc_z;
  wire start_PopNB_mioi_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  ActUnit_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB  start_PopNB_mioi
      (
      .this_vld(start_vld),
      .this_rdy(start_rdy),
      .this_dat(start_dat),
      .data_rsc_z(start_PopNB_mioi_data_rsc_z),
      .return_rsc_z(start_PopNB_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(start_PopNB_mioi_biwt_iff),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  ActUnit_ActUnit_ActUnitRun_start_PopNB_mioi_start_PopNB_mio_wait_ctrl ActUnit_ActUnitRun_start_PopNB_mioi_start_PopNB_mio_wait_ctrl_inst
      (
      .ActUnitRun_wen(ActUnitRun_wen),
      .ActUnitRun_wten(ActUnitRun_wten),
      .start_PopNB_mioi_oswt(start_PopNB_mioi_oswt),
      .start_PopNB_mioi_biwt(start_PopNB_mioi_biwt),
      .start_PopNB_mioi_bdwt(start_PopNB_mioi_bdwt),
      .start_PopNB_mioi_biwt_pff(start_PopNB_mioi_biwt_iff),
      .start_PopNB_mioi_oswt_pff(start_PopNB_mioi_oswt_pff)
    );
  ActUnit_ActUnit_ActUnitRun_start_PopNB_mioi_start_PopNB_mio_wait_dp ActUnit_ActUnitRun_start_PopNB_mioi_start_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .start_PopNB_mioi_data_rsc_z_mxwt(start_PopNB_mioi_data_rsc_z_mxwt),
      .start_PopNB_mioi_return_rsc_z_mxwt(start_PopNB_mioi_return_rsc_z_mxwt),
      .start_PopNB_mioi_biwt(start_PopNB_mioi_biwt),
      .start_PopNB_mioi_bdwt(start_PopNB_mioi_bdwt),
      .start_PopNB_mioi_data_rsc_z(start_PopNB_mioi_data_rsc_z),
      .start_PopNB_mioi_return_rsc_z(start_PopNB_mioi_return_rsc_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_rva_out_Push_mioi
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_rva_out_Push_mioi (
  clk, rst, rva_out_vld, rva_out_rdy, rva_out_dat, ActUnitRun_wten, rva_out_Push_mioi_oswt,
      rva_out_Push_mioi_wen_comp, rva_out_Push_mioi_m_data_rsc_dat_ActUnitRun, rva_out_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output rva_out_vld;
  input rva_out_rdy;
  output [511:0] rva_out_dat;
  input ActUnitRun_wten;
  input rva_out_Push_mioi_oswt;
  output rva_out_Push_mioi_wen_comp;
  input [511:0] rva_out_Push_mioi_m_data_rsc_dat_ActUnitRun;
  input rva_out_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire rva_out_Push_mioi_biwt;
  wire rva_out_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct;
  wire rva_out_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  ActUnit_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push
      rva_out_Push_mioi (
      .this_vld(rva_out_vld),
      .this_rdy(rva_out_rdy),
      .this_dat(rva_out_dat),
      .m_data_rsc_dat(rva_out_Push_mioi_m_data_rsc_dat_ActUnitRun),
      .ccs_ccore_start_rsc_dat(rva_out_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct),
      .ccs_ccore_done_sync_vld(rva_out_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  ActUnit_ActUnit_ActUnitRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl ActUnit_ActUnitRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl_inst
      (
      .ActUnitRun_wten(ActUnitRun_wten),
      .rva_out_Push_mioi_iswt0(rva_out_Push_mioi_oswt),
      .rva_out_Push_mioi_biwt(rva_out_Push_mioi_biwt),
      .rva_out_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct(rva_out_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct),
      .rva_out_Push_mioi_ccs_ccore_done_sync_vld(rva_out_Push_mioi_ccs_ccore_done_sync_vld),
      .rva_out_Push_mioi_iswt0_pff(rva_out_Push_mioi_oswt_pff)
    );
  assign rva_out_Push_mioi_wen_comp = (~ rva_out_Push_mioi_oswt) | rva_out_Push_mioi_biwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_act_port_PopNB_mioi
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_act_port_PopNB_mioi (
  clk, rst, act_port_vld, act_port_rdy, act_port_dat, ActUnitRun_wen, ActUnitRun_wten,
      act_port_PopNB_mioi_oswt, act_port_PopNB_mioi_data_data_rsc_z_mxwt, act_port_PopNB_mioi_return_rsc_z_mxwt,
      act_port_PopNB_mioi_oswt_pff
);
  input clk;
  input rst;
  input act_port_vld;
  output act_port_rdy;
  input [511:0] act_port_dat;
  input ActUnitRun_wen;
  input ActUnitRun_wten;
  input act_port_PopNB_mioi_oswt;
  output [511:0] act_port_PopNB_mioi_data_data_rsc_z_mxwt;
  output act_port_PopNB_mioi_return_rsc_z_mxwt;
  input act_port_PopNB_mioi_oswt_pff;


  // Interconnect Declarations
  wire act_port_PopNB_mioi_biwt;
  wire act_port_PopNB_mioi_bdwt;
  wire [511:0] act_port_PopNB_mioi_data_data_rsc_z;
  wire act_port_PopNB_mioi_return_rsc_z;
  wire act_port_PopNB_mioi_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  ActUnit_Connections_InBlocking_spec_ActVectorType_Connections_SYN_PORT_PopNB  act_port_PopNB_mioi
      (
      .this_vld(act_port_vld),
      .this_rdy(act_port_rdy),
      .this_dat(act_port_dat),
      .data_data_rsc_z(act_port_PopNB_mioi_data_data_rsc_z),
      .return_rsc_z(act_port_PopNB_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(act_port_PopNB_mioi_biwt_iff),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  ActUnit_ActUnit_ActUnitRun_act_port_PopNB_mioi_act_port_PopNB_mio_wait_ctrl ActUnit_ActUnitRun_act_port_PopNB_mioi_act_port_PopNB_mio_wait_ctrl_inst
      (
      .ActUnitRun_wen(ActUnitRun_wen),
      .ActUnitRun_wten(ActUnitRun_wten),
      .act_port_PopNB_mioi_oswt(act_port_PopNB_mioi_oswt),
      .act_port_PopNB_mioi_biwt(act_port_PopNB_mioi_biwt),
      .act_port_PopNB_mioi_bdwt(act_port_PopNB_mioi_bdwt),
      .act_port_PopNB_mioi_biwt_pff(act_port_PopNB_mioi_biwt_iff),
      .act_port_PopNB_mioi_oswt_pff(act_port_PopNB_mioi_oswt_pff)
    );
  ActUnit_ActUnit_ActUnitRun_act_port_PopNB_mioi_act_port_PopNB_mio_wait_dp ActUnit_ActUnitRun_act_port_PopNB_mioi_act_port_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .act_port_PopNB_mioi_data_data_rsc_z_mxwt(act_port_PopNB_mioi_data_data_rsc_z_mxwt),
      .act_port_PopNB_mioi_return_rsc_z_mxwt(act_port_PopNB_mioi_return_rsc_z_mxwt),
      .act_port_PopNB_mioi_biwt(act_port_PopNB_mioi_biwt),
      .act_port_PopNB_mioi_bdwt(act_port_PopNB_mioi_bdwt),
      .act_port_PopNB_mioi_data_data_rsc_z(act_port_PopNB_mioi_data_data_rsc_z),
      .act_port_PopNB_mioi_return_rsc_z(act_port_PopNB_mioi_return_rsc_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_rva_in_PopNB_mioi
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_rva_in_PopNB_mioi (
  clk, rst, rva_in_vld, rva_in_rdy, rva_in_dat, ActUnitRun_wen, ActUnitRun_wten,
      rva_in_PopNB_mioi_oswt, rva_in_PopNB_mioi_data_data_rsc_z_mxwt, rva_in_PopNB_mioi_data_addr_rsc_z_mxwt,
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt, rva_in_PopNB_mioi_return_rsc_z_mxwt,
      rva_in_PopNB_mioi_oswt_pff
);
  input clk;
  input rst;
  input rva_in_vld;
  output rva_in_rdy;
  input [600:0] rva_in_dat;
  input ActUnitRun_wen;
  input ActUnitRun_wten;
  input rva_in_PopNB_mioi_oswt;
  output [511:0] rva_in_PopNB_mioi_data_data_rsc_z_mxwt;
  output [11:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt;
  output rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  output rva_in_PopNB_mioi_return_rsc_z_mxwt;
  input rva_in_PopNB_mioi_oswt_pff;


  // Interconnect Declarations
  wire rva_in_PopNB_mioi_biwt;
  wire rva_in_PopNB_mioi_bdwt;
  wire [511:0] rva_in_PopNB_mioi_data_data_rsc_z;
  wire [23:0] rva_in_PopNB_mioi_data_addr_rsc_z;
  wire rva_in_PopNB_mioi_data_rw_rsc_z;
  wire rva_in_PopNB_mioi_return_rsc_z;
  wire [11:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt_pconst;
  wire rva_in_PopNB_mioi_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  ActUnit_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB
      rva_in_PopNB_mioi (
      .this_vld(rva_in_vld),
      .this_rdy(rva_in_rdy),
      .this_dat(rva_in_dat),
      .data_data_rsc_z(rva_in_PopNB_mioi_data_data_rsc_z),
      .data_addr_rsc_z(rva_in_PopNB_mioi_data_addr_rsc_z),
      .data_rw_rsc_z(rva_in_PopNB_mioi_data_rw_rsc_z),
      .return_rsc_z(rva_in_PopNB_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(rva_in_PopNB_mioi_biwt_iff),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  ActUnit_ActUnit_ActUnitRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl ActUnit_ActUnitRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl_inst
      (
      .ActUnitRun_wen(ActUnitRun_wen),
      .ActUnitRun_wten(ActUnitRun_wten),
      .rva_in_PopNB_mioi_oswt(rva_in_PopNB_mioi_oswt),
      .rva_in_PopNB_mioi_biwt(rva_in_PopNB_mioi_biwt),
      .rva_in_PopNB_mioi_bdwt(rva_in_PopNB_mioi_bdwt),
      .rva_in_PopNB_mioi_biwt_pff(rva_in_PopNB_mioi_biwt_iff),
      .rva_in_PopNB_mioi_oswt_pff(rva_in_PopNB_mioi_oswt_pff)
    );
  ActUnit_ActUnit_ActUnitRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp ActUnit_ActUnitRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_in_PopNB_mioi_data_data_rsc_z_mxwt(rva_in_PopNB_mioi_data_data_rsc_z_mxwt),
      .rva_in_PopNB_mioi_data_addr_rsc_z_mxwt(rva_in_PopNB_mioi_data_addr_rsc_z_mxwt_pconst),
      .rva_in_PopNB_mioi_data_rw_rsc_z_mxwt(rva_in_PopNB_mioi_data_rw_rsc_z_mxwt),
      .rva_in_PopNB_mioi_return_rsc_z_mxwt(rva_in_PopNB_mioi_return_rsc_z_mxwt),
      .rva_in_PopNB_mioi_biwt(rva_in_PopNB_mioi_biwt),
      .rva_in_PopNB_mioi_bdwt(rva_in_PopNB_mioi_bdwt),
      .rva_in_PopNB_mioi_data_data_rsc_z(rva_in_PopNB_mioi_data_data_rsc_z),
      .rva_in_PopNB_mioi_data_addr_rsc_z(rva_in_PopNB_mioi_data_addr_rsc_z),
      .rva_in_PopNB_mioi_data_rw_rsc_z(rva_in_PopNB_mioi_data_rw_rsc_z),
      .rva_in_PopNB_mioi_return_rsc_z(rva_in_PopNB_mioi_return_rsc_z)
    );
  assign rva_in_PopNB_mioi_data_addr_rsc_z_mxwt = rva_in_PopNB_mioi_data_addr_rsc_z_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun (
  clk, rst, start_vld, start_rdy, start_dat, act_port_vld, act_port_rdy, act_port_dat,
      rva_in_vld, rva_in_rdy, rva_in_dat, rva_out_vld, rva_out_rdy, rva_out_dat,
      output_port_vld, output_port_rdy, output_port_dat, done_vld, done_rdy, done_dat
);
  input clk;
  input rst;
  input start_vld;
  output start_rdy;
  input start_dat;
  input act_port_vld;
  output act_port_rdy;
  input [511:0] act_port_dat;
  input rva_in_vld;
  output rva_in_rdy;
  input [600:0] rva_in_dat;
  output rva_out_vld;
  input rva_out_rdy;
  output [511:0] rva_out_dat;
  output output_port_vld;
  input output_port_rdy;
  output [521:0] output_port_dat;
  output done_vld;
  input done_rdy;
  output done_dat;


  // Interconnect Declarations
  wire ActUnitRun_wen;
  wire ActUnitRun_wten;
  wire [511:0] rva_in_PopNB_mioi_data_data_rsc_z_mxwt;
  wire [11:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt;
  wire rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  wire rva_in_PopNB_mioi_return_rsc_z_mxwt;
  wire [511:0] act_port_PopNB_mioi_data_data_rsc_z_mxwt;
  wire act_port_PopNB_mioi_return_rsc_z_mxwt;
  wire rva_out_Push_mioi_wen_comp;
  wire start_PopNB_mioi_data_rsc_z_mxwt;
  wire start_PopNB_mioi_return_rsc_z_mxwt;
  wire output_port_Push_mioi_wen_comp;
  wire done_Push_mioi_wen_comp;
  wire Tanh_for_3_else_else_mul_1_cmp_en;
  wire [48:0] Tanh_for_3_else_else_mul_1_cmp_z;
  wire Tanh_for_3_else_else_mul_1_cmp_1_en;
  wire [48:0] Tanh_for_3_else_else_mul_1_cmp_1_z;
  wire Tanh_for_3_else_else_mul_1_cmp_2_en;
  wire [48:0] Tanh_for_3_else_else_mul_1_cmp_2_z;
  wire Tanh_for_3_else_else_mul_1_cmp_3_en;
  wire [48:0] Tanh_for_3_else_else_mul_1_cmp_3_z;
  wire Tanh_for_3_else_else_mul_1_cmp_4_en;
  wire [48:0] Tanh_for_3_else_else_mul_1_cmp_4_z;
  wire Tanh_for_3_else_else_mul_1_cmp_5_en;
  wire [48:0] Tanh_for_3_else_else_mul_1_cmp_5_z;
  wire Tanh_for_3_else_else_mul_1_cmp_6_en;
  wire [48:0] Tanh_for_3_else_else_mul_1_cmp_6_z;
  wire Tanh_for_3_else_else_mul_1_cmp_7_en;
  wire [48:0] Tanh_for_3_else_else_mul_1_cmp_7_z;
  wire Tanh_for_3_else_else_mul_1_cmp_8_en;
  wire [48:0] Tanh_for_3_else_else_mul_1_cmp_8_z;
  wire Tanh_for_3_else_else_mul_1_cmp_9_en;
  wire [48:0] Tanh_for_3_else_else_mul_1_cmp_9_z;
  wire Tanh_for_3_else_else_mul_1_cmp_10_en;
  wire [48:0] Tanh_for_3_else_else_mul_1_cmp_10_z;
  wire Tanh_for_3_else_else_mul_1_cmp_11_en;
  wire [48:0] Tanh_for_3_else_else_mul_1_cmp_11_z;
  wire Tanh_for_3_else_else_mul_1_cmp_12_en;
  wire [48:0] Tanh_for_3_else_else_mul_1_cmp_12_z;
  wire Tanh_for_3_else_else_mul_1_cmp_13_en;
  wire [48:0] Tanh_for_3_else_else_mul_1_cmp_13_z;
  wire Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_en;
  wire [100:0] Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_z;
  wire Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_1_en;
  wire [100:0] Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_1_z;
  wire Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_2_en;
  wire [100:0] Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_2_z;
  wire Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_3_en;
  wire [100:0] Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_3_z;
  wire Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_4_en;
  wire [100:0] Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_4_z;
  wire Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_5_en;
  wire [100:0] Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_5_z;
  wire Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_6_en;
  wire [100:0] Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_6_z;
  wire Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_7_en;
  wire [100:0] Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_7_z;
  wire Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_8_en;
  wire [100:0] Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_8_z;
  wire Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_9_en;
  wire [100:0] Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_9_z;
  wire Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_10_en;
  wire [100:0] Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_10_z;
  wire Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_11_en;
  wire [100:0] Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_11_z;
  wire Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_12_en;
  wire [100:0] Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_12_z;
  wire Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_13_en;
  wire [100:0] Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_13_z;
  wire Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_14_en;
  wire [100:0] Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_14_z;
  wire Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_15_en;
  wire [100:0] Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_15_z;
  wire Tanh_for_1_else_else_mul_cmp_en;
  wire [74:0] Tanh_for_1_else_else_mul_cmp_z;
  wire Tanh_for_1_else_else_mul_cmp_1_en;
  wire [74:0] Tanh_for_1_else_else_mul_cmp_1_z;
  wire Tanh_for_1_else_else_mul_cmp_2_en;
  wire [74:0] Tanh_for_1_else_else_mul_cmp_2_z;
  wire Tanh_for_1_else_else_mul_cmp_3_en;
  wire [74:0] Tanh_for_1_else_else_mul_cmp_3_z;
  wire Tanh_for_1_else_else_mul_cmp_4_en;
  wire [74:0] Tanh_for_1_else_else_mul_cmp_4_z;
  wire Tanh_for_1_else_else_mul_cmp_5_en;
  wire [74:0] Tanh_for_1_else_else_mul_cmp_5_z;
  wire Tanh_for_1_else_else_mul_cmp_6_en;
  wire [74:0] Tanh_for_1_else_else_mul_cmp_6_z;
  wire Tanh_for_1_else_else_mul_cmp_7_en;
  wire [74:0] Tanh_for_1_else_else_mul_cmp_7_z;
  wire Tanh_for_1_else_else_mul_cmp_8_en;
  wire [74:0] Tanh_for_1_else_else_mul_cmp_8_z;
  wire Tanh_for_1_else_else_mul_cmp_9_en;
  wire [74:0] Tanh_for_1_else_else_mul_cmp_9_z;
  wire Tanh_for_1_else_else_mul_cmp_10_en;
  wire [74:0] Tanh_for_1_else_else_mul_cmp_10_z;
  wire Tanh_for_1_else_else_mul_cmp_11_en;
  wire [74:0] Tanh_for_1_else_else_mul_cmp_11_z;
  wire Tanh_for_1_else_else_mul_cmp_12_en;
  wire [74:0] Tanh_for_1_else_else_mul_cmp_12_z;
  wire Tanh_for_1_else_else_mul_cmp_13_en;
  wire [74:0] Tanh_for_1_else_else_mul_cmp_13_z;
  wire Tanh_for_1_else_else_mul_cmp_14_en;
  wire [74:0] Tanh_for_1_else_else_mul_cmp_14_z;
  wire Tanh_for_1_else_else_mul_cmp_15_en;
  wire [74:0] Tanh_for_1_else_else_mul_cmp_15_z;
  wire Tanh_for_1_else_else_mul_1_cmp_en;
  wire [53:0] Tanh_for_1_else_else_mul_1_cmp_z;
  wire Tanh_for_1_else_else_mul_1_cmp_1_en;
  wire [53:0] Tanh_for_1_else_else_mul_1_cmp_1_z;
  wire [4:0] fsm_output;
  wire act_config_InstIncr_if_act_config_InstIncr_if_if_nor_tmp;
  wire act_config_InstIncr_if_equal_1_tmp;
  wire [6:0] operator_6_false_acc_tmp;
  wire [7:0] nl_operator_6_false_acc_tmp;
  wire ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_2_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_less_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_less_1_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_less_2_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_less_3_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_less_4_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_less_5_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_less_6_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_less_7_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_less_8_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_less_9_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_less_10_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_less_11_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_less_12_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_less_13_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_1_less_14_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_less_14_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_1_less_15_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_less_15_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_less_tmp_1;
  wire operator_32_8_true_AC_TRN_AC_WRAP_3_less_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_less_1_tmp_1;
  wire operator_32_8_true_AC_TRN_AC_WRAP_3_less_1_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_less_2_tmp_1;
  wire operator_32_8_true_AC_TRN_AC_WRAP_3_less_2_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_less_3_tmp_1;
  wire operator_32_8_true_AC_TRN_AC_WRAP_3_less_3_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_less_4_tmp_1;
  wire operator_32_8_true_AC_TRN_AC_WRAP_3_less_4_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_less_5_tmp_1;
  wire operator_32_8_true_AC_TRN_AC_WRAP_3_less_5_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_less_6_tmp_1;
  wire operator_32_8_true_AC_TRN_AC_WRAP_3_less_6_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_less_7_tmp_1;
  wire operator_32_8_true_AC_TRN_AC_WRAP_3_less_7_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_less_8_tmp_1;
  wire operator_32_8_true_AC_TRN_AC_WRAP_3_less_8_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_less_9_tmp_1;
  wire operator_32_8_true_AC_TRN_AC_WRAP_3_less_9_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_less_10_tmp_1;
  wire operator_32_8_true_AC_TRN_AC_WRAP_3_less_10_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_less_11_tmp_1;
  wire operator_32_8_true_AC_TRN_AC_WRAP_3_less_11_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_less_12_tmp_1;
  wire operator_32_8_true_AC_TRN_AC_WRAP_3_less_12_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_less_13_tmp_1;
  wire operator_32_8_true_AC_TRN_AC_WRAP_3_less_13_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_less_14_tmp_1;
  wire operator_32_8_true_AC_TRN_AC_WRAP_3_less_14_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_less_15_tmp_1;
  wire operator_32_8_true_AC_TRN_AC_WRAP_3_less_15_tmp;
  wire [7:0] act_config_in_InstFetch_mux_tmp;
  wire [4:0] while_mux_55_tmp;
  wire while_and_1_tmp;
  wire and_dcpl_9;
  wire and_dcpl_13;
  wire and_dcpl_47;
  wire and_dcpl_51;
  wire and_dcpl_78;
  wire and_dcpl_162;
  wire and_dcpl_366;
  wire and_dcpl_368;
  wire and_dcpl_369;
  wire and_dcpl_370;
  wire or_tmp_68;
  wire mux_tmp_55;
  wire and_dcpl_374;
  wire and_dcpl_377;
  wire and_dcpl_379;
  wire or_tmp_111;
  wire and_dcpl_553;
  wire and_dcpl_554;
  wire and_dcpl_556;
  wire and_dcpl_557;
  wire and_dcpl_559;
  wire and_dcpl_560;
  wire and_dcpl_562;
  wire or_tmp_126;
  wire and_dcpl_563;
  wire and_dcpl_564;
  wire and_dcpl_565;
  wire and_dcpl_566;
  wire and_dcpl_568;
  wire and_dcpl_569;
  wire and_dcpl_570;
  wire and_dcpl_571;
  wire and_dcpl_572;
  wire and_dcpl_573;
  wire and_dcpl_574;
  wire and_dcpl_575;
  wire and_dcpl_576;
  wire and_dcpl_577;
  wire and_dcpl_578;
  wire and_dcpl_579;
  wire and_dcpl_581;
  wire and_dcpl_582;
  wire and_dcpl_583;
  wire and_dcpl_584;
  wire and_dcpl_585;
  wire and_dcpl_586;
  wire and_dcpl_587;
  wire or_tmp_131;
  wire or_tmp_133;
  wire or_tmp_134;
  wire or_tmp_135;
  wire or_tmp_136;
  wire and_tmp_9;
  wire or_tmp_139;
  wire or_tmp_140;
  wire and_tmp_11;
  wire not_tmp_248;
  wire nand_tmp_3;
  wire or_tmp_146;
  wire or_tmp_147;
  wire or_tmp_148;
  wire or_tmp_151;
  wire or_tmp_159;
  wire or_tmp_161;
  wire or_tmp_162;
  wire or_tmp_163;
  wire or_tmp_164;
  wire or_tmp_167;
  wire or_tmp_168;
  wire not_tmp_255;
  wire nand_tmp_9;
  wire or_tmp_174;
  wire or_tmp_175;
  wire or_tmp_176;
  wire or_tmp_179;
  wire and_dcpl_590;
  wire and_dcpl_591;
  wire and_dcpl_592;
  wire or_tmp_184;
  wire and_dcpl_596;
  wire and_dcpl_599;
  wire and_dcpl_600;
  wire not_tmp_262;
  wire or_tmp_198;
  wire and_dcpl_604;
  wire or_tmp_211;
  wire or_tmp_213;
  wire and_dcpl_609;
  wire and_dcpl_612;
  wire and_dcpl_613;
  wire and_dcpl_614;
  wire or_tmp_215;
  wire and_tmp_39;
  wire or_tmp_229;
  wire and_dcpl_616;
  wire and_dcpl_620;
  wire and_dcpl_621;
  wire or_tmp_237;
  wire mux_tmp_169;
  wire or_tmp_249;
  wire or_dcpl_290;
  wire and_dcpl_668;
  wire and_dcpl_746;
  wire and_dcpl_747;
  wire and_dcpl_748;
  wire not_tmp_311;
  wire and_dcpl_767;
  wire and_dcpl_768;
  wire and_dcpl_770;
  wire and_dcpl_774;
  wire and_dcpl_775;
  wire and_dcpl_786;
  wire and_dcpl_788;
  wire and_dcpl_789;
  wire and_dcpl_794;
  wire or_dcpl_296;
  wire or_dcpl_297;
  wire or_dcpl_299;
  wire or_dcpl_300;
  wire and_dcpl_797;
  wire or_dcpl_301;
  wire or_dcpl_303;
  wire or_dcpl_304;
  wire and_dcpl_798;
  wire and_dcpl_799;
  wire or_dcpl_310;
  wire or_dcpl_320;
  wire or_dcpl_322;
  wire and_dcpl_802;
  wire and_dcpl_803;
  wire and_dcpl_805;
  wire or_dcpl_328;
  wire or_dcpl_329;
  wire or_dcpl_330;
  wire or_dcpl_332;
  wire or_dcpl_333;
  wire or_dcpl_335;
  wire or_dcpl_338;
  wire or_dcpl_341;
  wire or_dcpl_342;
  wire or_dcpl_347;
  wire or_dcpl_348;
  wire or_dcpl_353;
  wire or_dcpl_358;
  wire or_dcpl_359;
  wire or_dcpl_364;
  wire or_dcpl_369;
  wire or_dcpl_370;
  wire or_dcpl_375;
  wire or_dcpl_380;
  wire or_dcpl_381;
  wire or_dcpl_386;
  wire or_dcpl_387;
  wire or_dcpl_392;
  wire or_dcpl_397;
  wire or_dcpl_402;
  wire or_dcpl_407;
  wire or_dcpl_412;
  wire or_dcpl_417;
  wire not_tmp_347;
  wire or_dcpl_423;
  wire and_dcpl_814;
  wire and_dcpl_829;
  wire or_tmp_315;
  wire mux_tmp_196;
  wire mux_tmp_197;
  wire nor_tmp_46;
  wire and_dcpl_831;
  wire and_dcpl_832;
  wire or_tmp_317;
  wire or_dcpl_440;
  wire or_dcpl_442;
  wire mux_tmp_203;
  wire and_dcpl_834;
  wire or_tmp_318;
  wire or_dcpl_443;
  wire and_dcpl_849;
  wire or_tmp_322;
  wire mux_tmp_214;
  wire and_dcpl_852;
  wire or_dcpl_447;
  wire or_dcpl_448;
  wire or_dcpl_449;
  wire and_dcpl_853;
  wire and_dcpl_854;
  wire and_dcpl_855;
  wire and_dcpl_856;
  wire and_dcpl_857;
  wire or_dcpl_450;
  wire or_dcpl_451;
  wire or_dcpl_452;
  wire or_dcpl_453;
  wire or_dcpl_455;
  wire or_dcpl_456;
  wire and_dcpl_860;
  wire and_dcpl_861;
  wire or_dcpl_457;
  wire or_dcpl_458;
  wire or_dcpl_460;
  wire or_dcpl_461;
  wire or_dcpl_462;
  wire and_dcpl_864;
  wire and_dcpl_865;
  wire and_dcpl_866;
  wire and_dcpl_867;
  wire or_dcpl_463;
  wire or_dcpl_464;
  wire or_dcpl_465;
  wire or_dcpl_466;
  wire or_dcpl_468;
  wire or_dcpl_469;
  wire and_dcpl_870;
  wire and_dcpl_871;
  wire or_dcpl_470;
  wire or_dcpl_471;
  wire or_dcpl_473;
  wire or_dcpl_474;
  wire and_dcpl_874;
  wire or_dcpl_475;
  wire or_dcpl_477;
  wire and_dcpl_877;
  wire or_dcpl_478;
  wire or_dcpl_480;
  wire or_dcpl_482;
  wire or_dcpl_484;
  wire or_dcpl_486;
  wire or_dcpl_487;
  wire or_dcpl_489;
  wire and_dcpl_888;
  wire or_dcpl_490;
  wire or_dcpl_492;
  wire and_dcpl_891;
  wire or_dcpl_493;
  wire or_dcpl_495;
  wire or_dcpl_497;
  wire or_dcpl_499;
  wire and_dcpl_900;
  wire or_tmp_323;
  wire and_dcpl_901;
  wire and_dcpl_903;
  wire and_dcpl_906;
  wire and_dcpl_908;
  wire and_dcpl_909;
  wire and_dcpl_916;
  wire or_dcpl_503;
  wire or_dcpl_504;
  wire or_dcpl_507;
  wire or_dcpl_508;
  wire and_dcpl_923;
  wire and_dcpl_924;
  wire or_dcpl_523;
  wire and_dcpl_929;
  wire or_dcpl_526;
  wire and_dcpl_958;
  wire and_dcpl_959;
  wire or_dcpl_541;
  wire and_dcpl_964;
  wire or_dcpl_544;
  wire and_dcpl_997;
  wire or_tmp_330;
  wire or_tmp_331;
  wire and_dcpl_1001;
  wire and_dcpl_1006;
  wire and_dcpl_1007;
  wire or_dcpl_561;
  wire or_dcpl_563;
  wire or_dcpl_566;
  wire or_dcpl_567;
  wire or_dcpl_582;
  wire or_dcpl_583;
  wire or_dcpl_586;
  wire or_dcpl_601;
  wire or_dcpl_602;
  wire or_dcpl_605;
  wire or_dcpl_620;
  wire or_dcpl_621;
  wire or_dcpl_624;
  wire act_config_InstIncr_act_config_InstIncr_if_and_svs_1;
  reg [7:0] act_config_output_counter_sva_dfm_3;
  wire [8:0] operator_8_false_acc_sdt_sva_1;
  wire [9:0] nl_operator_8_false_acc_sdt_sva_1;
  wire [4:0] ActUnit_RunInst_case_2_for_i_4_0_sva_2;
  wire [5:0] nl_ActUnit_RunInst_case_2_for_i_4_0_sva_2;
  reg ActUnit_RunInst_switch_lp_and_48_tmp;
  reg ActUnit_RunInst_switch_lp_equal_tmp_2;
  reg is_start_sva;
  reg while_nor_48_itm;
  reg Gelu_for_and_2_cse_sva;
  reg ActUnit_RunInst_switch_lp_equal_tmp_8;
  reg ActUnit_RunInst_switch_lp_equal_tmp_7;
  reg ActUnit_RunInst_switch_lp_equal_tmp_6;
  reg ActUnit_RunInst_switch_lp_equal_tmp_5;
  reg ActUnit_RunInst_switch_lp_equal_tmp_4;
  reg ActUnit_RunInst_switch_lp_and_32_tmp;
  reg while_nor_32_itm;
  reg ActUnit_RunInst_switch_lp_and_16_tmp;
  reg while_nor_16_itm;
  reg ActUnit_PushOutput_if_for_and_stg_2_7_sva;
  reg ActUnit_RunInst_switch_lp_and_tmp;
  reg while_nor_itm;
  reg Tanh_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  reg Tanh_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs;
  reg Tanh_for_15_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  reg Tanh_for_15_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs;
  reg Tanh_for_14_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  reg Tanh_for_14_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs;
  reg Tanh_for_13_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  reg Tanh_for_13_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs;
  reg Tanh_for_12_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  reg Tanh_for_12_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs;
  reg Tanh_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  reg Tanh_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs;
  reg Tanh_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  reg Tanh_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs;
  reg Tanh_for_9_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  reg Tanh_for_9_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs;
  reg Tanh_for_8_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  reg Tanh_for_8_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs;
  reg Tanh_for_7_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  reg Tanh_for_7_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs;
  reg Tanh_for_6_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  reg Tanh_for_6_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs;
  reg Tanh_for_5_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  reg Tanh_for_5_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs;
  reg Tanh_for_4_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  reg Tanh_for_4_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs;
  reg Tanh_for_3_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  reg Tanh_for_3_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs;
  reg Tanh_for_2_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  reg Tanh_for_2_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs;
  reg Tanh_for_1_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  reg Tanh_for_1_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs;
  wire act_config_ActConfigRead_unequal_tmp_1;
  wire ActUnit_DecodeAxi_if_or_7_tmp_1;
  wire while_and_88_tmp_1;
  wire ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_mx1;
  wire ActUnit_DecodeAxi_rva_in_reg_rw_sva_mx1;
  wire act_config_ActConfigRead_else_unequal_tmp_1;
  wire ActUnit_DecodeAxiRead_unequal_tmp_1;
  wire Tanh_for_nor_cse_sva_mx0w0;
  wire ActUnit_RunInst_switch_lp_nor_tmp_mx0;
  reg act_config_is_zero_first_sva_dfm_4;
  reg w_load_lpi_1_dfm_1;
  reg is_incr_lpi_1_dfm_1;
  reg ActUnit_CheckStart_start_reg_sva;
  reg act_config_is_valid_sva;
  reg ActUnit_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva;
  reg [7:0] act_config_inst_regs_16_sva_dfm_6;
  reg [7:0] act_config_inst_regs_17_sva_dfm_6;
  reg [7:0] act_config_inst_regs_18_sva_dfm_6;
  reg [7:0] act_config_inst_regs_19_sva_dfm_6;
  reg [7:0] act_config_inst_regs_20_sva_dfm_6;
  reg [7:0] act_config_inst_regs_21_sva_dfm_6;
  reg [7:0] act_config_inst_regs_22_sva_dfm_6;
  reg [7:0] act_config_inst_regs_23_sva_dfm_6;
  reg [7:0] act_config_inst_regs_24_sva_dfm_6;
  reg [7:0] act_config_inst_regs_25_sva_dfm_6;
  reg [7:0] act_config_inst_regs_26_sva_dfm_6;
  reg [7:0] act_config_inst_regs_27_sva_dfm_6;
  reg [7:0] act_config_inst_regs_28_sva_dfm_6;
  reg [7:0] act_config_inst_regs_29_sva_dfm_6;
  reg [7:0] act_config_inst_regs_30_sva_dfm_6;
  reg [7:0] act_config_inst_regs_31_sva_dfm_6;
  reg [4:0] act_config_inst_counter_sva_dfm_3;
  wire [7:0] ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_23_4_mx1_tmp_7_0;
  reg act_config_is_zero_first_sva;
  reg [5:0] act_config_in_InstFetch_return_sva_7_2;
  reg Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs;
  reg Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  reg Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs;
  reg Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  reg Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs;
  reg Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs;
  reg Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs;
  reg Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  reg Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs;
  reg Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  reg Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs;
  reg Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  reg Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs;
  reg Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  reg Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  reg Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs;
  reg Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs;
  reg Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  reg Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs;
  reg Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  reg Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs;
  reg Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  reg Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs;
  reg Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  reg Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs;
  reg Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  reg Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs;
  reg Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  reg Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs;
  reg Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  reg Gelu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs;
  reg Gelu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs;
  reg Gelu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs;
  reg Gelu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs;
  reg Gelu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs;
  reg Gelu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs;
  reg Gelu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs;
  reg Gelu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs;
  reg Gelu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs;
  reg Gelu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs;
  reg Gelu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs;
  reg Gelu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs;
  reg Gelu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs;
  reg Gelu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs;
  reg Gelu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs;
  reg Gelu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs;
  reg Gelu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs;
  reg Gelu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs;
  reg Gelu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs;
  reg Gelu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs;
  reg Gelu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs;
  reg Gelu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs;
  reg Gelu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs;
  reg Gelu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs;
  reg Gelu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs;
  reg Gelu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs;
  reg w_axi_rsp_lpi_1_dfm_1;
  reg act_read_req_valid_lpi_1_dfm_6;
  reg [3:0] ActUnit_PushOutput_if_for_i_4_0_sva_3_0;
  reg [1:0] nvhls_get_slc_2U_NVUINT8_return_3_sva;
  reg while_asn_262_itm;
  reg Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  reg Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  wire ActUnit_RunInst_switch_lp_equal_tmp_1_mx0w0;
  wire ActUnit_RunInst_switch_lp_equal_tmp_2_mx0w0;
  wire ActUnit_RunInst_switch_lp_equal_tmp_3_mx0w0;
  wire ActUnit_RunInst_switch_lp_equal_tmp_4_mx0w0;
  wire ActUnit_RunInst_switch_lp_equal_tmp_5_mx0w0;
  wire ActUnit_RunInst_switch_lp_equal_tmp_6_mx0w0;
  wire ActUnit_RunInst_switch_lp_equal_tmp_7_mx0w0;
  wire ActUnit_RunInst_switch_lp_equal_tmp_8_mx0w0;
  wire [1:0] nvhls_get_slc_2U_NVUINT8_return_3_sva_1;
  reg [7:0] act_config_inst_regs_0_sva_dfm_5;
  reg [7:0] act_config_inst_regs_1_sva_dfm_5;
  reg [7:0] act_config_inst_regs_2_sva_dfm_5;
  reg [7:0] act_config_inst_regs_3_sva_dfm_5;
  reg [7:0] act_config_inst_regs_4_sva_dfm_5;
  reg [7:0] act_config_inst_regs_5_sva_dfm_5;
  reg [7:0] act_config_inst_regs_6_sva_dfm_5;
  reg [7:0] act_config_inst_regs_7_sva_dfm_5;
  reg [7:0] act_config_inst_regs_8_sva_dfm_5;
  reg [7:0] act_config_inst_regs_9_sva_dfm_5;
  reg [7:0] act_config_inst_regs_10_sva_dfm_5;
  reg [7:0] act_config_inst_regs_11_sva_dfm_5;
  reg [7:0] act_config_inst_regs_12_sva_dfm_5;
  reg [7:0] act_config_inst_regs_13_sva_dfm_5;
  reg [7:0] act_config_inst_regs_14_sva_dfm_5;
  reg [7:0] act_config_inst_regs_15_sva_dfm_5;
  reg [25:0] reg_nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6;
  reg [25:0] reg_nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6;
  reg [25:0] reg_nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6;
  reg [25:0] reg_nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6;
  reg [25:0] reg_nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6;
  reg [25:0] reg_nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6;
  reg [25:0] reg_nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6;
  reg [25:0] reg_nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6;
  reg [25:0] reg_nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6;
  reg [25:0] reg_nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6;
  reg [25:0] reg_nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6;
  reg [25:0] reg_nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6;
  reg [25:0] reg_ActUnit_RunInst_case_11_nv_scvector_cctor_data_0_ftd_6;
  reg [7:0] reg_ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_23_4_ftd_12;
  wire act_mem_banks_write_if_for_if_mux_cse;
  wire act_mem_banks_write_if_for_if_mux_1_cse;
  wire act_mem_banks_read_for_mux_cse;
  wire act_mem_banks_read_for_mux_1_cse;
  reg reg_Tanh_for_1_else_else_mul_1_cmp_cgo_ir_1_cse;
  reg reg_Tanh_for_1_else_else_mul_1_cmp_cgo_ir_cse;
  reg reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_15_cse;
  reg reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_14_cse;
  reg reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_13_cse;
  reg reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_12_cse;
  reg reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_11_cse;
  reg reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_10_cse;
  reg reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_9_cse;
  reg reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_8_cse;
  reg reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_7_cse;
  reg reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_6_cse;
  reg reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_5_cse;
  reg reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_4_cse;
  reg reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_3_cse;
  reg reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_2_cse;
  reg reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_1_cse;
  reg reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_cse;
  reg reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_15_cse;
  reg reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_14_cse;
  reg reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_13_cse;
  reg reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_12_cse;
  reg reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_11_cse;
  reg reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_10_cse;
  reg reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_9_cse;
  reg reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_8_cse;
  reg reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_7_cse;
  reg reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_6_cse;
  reg reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_5_cse;
  reg reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_4_cse;
  reg reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_3_cse;
  reg reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_2_cse;
  reg reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_1_cse;
  reg reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_cse;
  reg reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_13_cse;
  reg reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_12_cse;
  reg reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_11_cse;
  reg reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_10_cse;
  reg reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_9_cse;
  reg reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_8_cse;
  reg reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_7_cse;
  reg reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_6_cse;
  reg reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_5_cse;
  reg reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_4_cse;
  reg reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_3_cse;
  reg reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_2_cse;
  reg reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_1_cse;
  reg reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_cse;
  reg reg_done_Push_mioi_iswt0_cse;
  reg reg_output_port_Push_mioi_iswt0_cse;
  reg reg_start_PopNB_mioi_iswt0_cse;
  reg reg_rva_out_Push_mioi_iswt0_cse;
  reg reg_act_port_PopNB_mioi_iswt0_cse;
  reg reg_rva_in_PopNB_mioi_iswt0_cse;
  wire act_config_num_inst_and_cse;
  wire rva_out_reg_data_and_cse;
  wire act_mem_banks_bank_a_and_cse;
  wire act_mem_banks_bank_a_and_1_cse;
  wire act_mem_banks_bank_a_and_2_cse;
  wire act_mem_banks_bank_a_and_3_cse;
  wire act_mem_banks_bank_a_and_4_cse;
  wire act_mem_banks_bank_a_and_5_cse;
  wire act_mem_banks_bank_a_and_6_cse;
  wire act_mem_banks_bank_a_and_7_cse;
  wire act_mem_banks_bank_a_and_8_cse;
  wire act_mem_banks_bank_a_and_9_cse;
  wire act_mem_banks_bank_a_and_10_cse;
  wire act_mem_banks_bank_a_and_11_cse;
  wire act_mem_banks_bank_a_and_12_cse;
  wire act_mem_banks_bank_a_and_13_cse;
  wire act_mem_banks_bank_a_and_14_cse;
  wire act_mem_banks_bank_a_and_15_cse;
  wire act_mem_banks_bank_a_and_16_cse;
  wire act_mem_banks_bank_a_and_17_cse;
  wire act_mem_banks_bank_a_and_18_cse;
  wire act_mem_banks_bank_a_and_19_cse;
  wire act_mem_banks_bank_a_and_20_cse;
  wire act_mem_banks_bank_a_and_21_cse;
  wire act_mem_banks_bank_a_and_22_cse;
  wire act_mem_banks_bank_a_and_23_cse;
  wire act_mem_banks_bank_a_and_24_cse;
  wire act_mem_banks_bank_a_and_25_cse;
  wire act_mem_banks_bank_a_and_26_cse;
  wire act_mem_banks_bank_a_and_27_cse;
  wire act_mem_banks_bank_a_and_28_cse;
  wire act_mem_banks_bank_a_and_29_cse;
  wire act_mem_banks_bank_a_and_30_cse;
  wire act_mem_banks_bank_a_and_31_cse;
  wire act_config_inst_regs_and_4_cse;
  wire act_config_inst_regs_and_20_cse;
  wire act_regs_data_and_cse;
  wire act_mem_banks_read_read_data_and_cse;
  wire act_port_read_out_data_and_cse;
  wire rva_out_reg_data_and_16_cse;
  wire ActUnit_RunInst_switch_lp_and_802_cse;
  wire ActUnit_RunInst_switch_lp_and_808_cse;
  wire ActUnit_RunInst_case_3_act_port_reg_data_and_cse;
  wire act_config_output_counter_and_1_cse;
  wire Gelu_for_else_else_and_1_cse;
  wire nor_333_cse;
  wire nor_28_cse;
  wire and_1101_cse;
  wire or_992_cse;
  wire and_1103_cse;
  wire and_1104_cse;
  wire nor_57_cse;
  wire nand_180_cse;
  wire nand_181_cse;
  wire nor_61_cse;
  wire nand_195_cse;
  wire nor_139_cse;
  reg ActUnit_RunInst_switch_lp_nor_tmp;
  wire Tanh_for_and_2_cse_sva_mx0w0;
  wire ActUnit_RunInst_switch_lp_and_48_tmp_mx0w0;
  wire Tanh_for_and_cse_sva_mx0w0;
  wire ActUnit_RunInst_switch_lp_and_32_tmp_mx0w1;
  wire Tanh_for_and_1_cse_sva_mx0w0;
  wire ActUnit_RunInst_switch_lp_and_16_tmp_mx0w1;
  wire ActUnit_RunInst_switch_lp_and_tmp_mx0w0;
  wire Tanh_for_and_85_m1c;
  wire while_and_203_cse;
  wire while_and_204_cse;
  reg reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_nor_cse;
  reg reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_2_cse;
  reg reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_1_cse;
  reg reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_cse;
  wire and_1046_cse;
  wire mux_51_cse;
  reg [46:0] Gelu_for_else_else_slc_Tanh_for_1_else_else_mul_cmp_z_46_0_itm;
  wire Tanh_for_else_else_or_1_cse;
  wire Tanh_for_or_cse;
  wire Tanh_for_and_87_cse;
  wire and_812_rmff;
  wire and_811_rmff;
  wire and_810_rmff;
  wire and_809_rmff;
  wire and_808_rmff;
  wire and_807_rmff;
  wire and_806_rmff;
  wire and_805_rmff;
  wire and_804_rmff;
  wire and_803_rmff;
  wire and_802_rmff;
  wire and_801_rmff;
  wire and_800_rmff;
  wire and_799_rmff;
  wire and_794_rmff;
  wire and_789_rmff;
  wire and_784_rmff;
  wire and_779_rmff;
  wire and_774_rmff;
  wire and_769_rmff;
  wire and_764_rmff;
  wire and_759_rmff;
  wire and_754_rmff;
  wire and_749_rmff;
  wire and_744_rmff;
  wire and_739_rmff;
  wire and_734_rmff;
  wire and_729_rmff;
  wire and_724_rmff;
  wire and_719_rmff;
  wire and_713_rmff;
  wire and_705_rmff;
  wire and_701_rmff;
  wire and_697_rmff;
  wire and_693_rmff;
  wire and_689_rmff;
  wire and_685_rmff;
  wire and_681_rmff;
  wire and_677_rmff;
  wire and_673_rmff;
  wire and_669_rmff;
  wire and_665_rmff;
  wire and_658_rmff;
  wire and_633_rmff;
  wire and_626_rmff;
  wire and_621_rmff;
  wire and_617_rmff;
  wire and_605_rmff;
  wire and_837_rmff;
  wire and_835_rmff;
  wire and_830_rmff;
  wire and_826_rmff;
  wire and_823_rmff;
  wire and_819_rmff;
  reg [7:0] act_config_output_addr_base_sva;
  reg [30:0] ActUnit_RunInst_case_15_nv_scvector_cctor_data_0_sva_30_0;
  reg [30:0] nv_scvector_cctor_nv_scvector_6_for_5_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0;
  reg [30:0] nv_scvector_cctor_nv_scvector_6_for_7_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0;
  reg [30:0] nv_scvector_cctor_nv_scvector_6_for_14_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0;
  reg [30:0] nv_scvector_cctor_nv_scvector_6_for_11_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0;
  reg [30:0] nv_scvector_cctor_nv_scvector_6_for_2_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0;
  reg [30:0] nv_scvector_cctor_nv_scvector_6_for_3_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0;
  reg [30:0] nv_scvector_cctor_nv_scvector_6_for_4_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0;
  reg [30:0] nv_scvector_cctor_nv_scvector_6_for_6_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0;
  reg [30:0] nv_scvector_cctor_nv_scvector_6_for_15_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0;
  reg [30:0] nv_scvector_cctor_nv_scvector_6_for_10_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0;
  reg [46:0] Gelu_for_else_else_slc_Tanh_for_1_else_else_mul_cmp_12_z_46_0_itm;
  reg [30:0] nv_scvector_cctor_nv_scvector_6_for_12_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0;
  reg [30:0] nv_scvector_cctor_nv_scvector_6_for_9_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0;
  reg [30:0] nv_scvector_cctor_nv_scvector_6_for_16_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0;
  reg [46:0] Gelu_for_else_else_slc_Tanh_for_1_else_else_mul_1_cmp_z_46_0_itm;
  reg [46:0] Gelu_for_else_else_slc_Tanh_for_1_else_else_mul_cmp_13_z_46_0_itm;
  reg [30:0] nv_scvector_cctor_nv_scvector_6_for_8_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0;
  reg [30:0] nv_scvector_cctor_nv_scvector_6_for_13_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0;
  reg [46:0] Gelu_for_else_else_slc_Tanh_for_1_else_else_mul_cmp_15_z_46_0_itm;
  reg [30:0] nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0;
  reg [30:0] nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0;
  reg [30:0] nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0;
  reg [30:0] nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0;
  reg [30:0] nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0;
  reg [30:0] nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0;
  reg [30:0] nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0;
  reg [30:0] nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0;
  reg [30:0] nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0;
  reg [30:0] nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0;
  reg [30:0] nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0;
  reg [30:0] nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0;
  reg [30:0] nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0;
  reg [30:0] nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0;
  reg [31:0] rva_out_reg_data_511_480_sva_dfm_3;
  wire [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_511_480_mx1;
  reg [31:0] rva_out_reg_data_479_448_sva_dfm_3;
  wire [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_479_448_mx1;
  reg [31:0] rva_out_reg_data_447_416_sva_dfm_3;
  wire [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_447_416_mx1;
  reg [31:0] rva_out_reg_data_415_384_sva_dfm_3;
  wire [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_415_384_mx1;
  reg [31:0] rva_out_reg_data_383_352_sva_dfm_3;
  wire [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_383_352_mx1;
  reg [31:0] rva_out_reg_data_351_320_sva_dfm_3;
  wire [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_351_320_mx1;
  reg [31:0] rva_out_reg_data_319_288_sva_dfm_3;
  wire [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_319_288_mx1;
  reg [31:0] rva_out_reg_data_287_256_sva_dfm_3;
  wire [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_287_256_mx1;
  reg [31:0] rva_out_reg_data_255_224_sva_dfm_3;
  wire [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_255_224_mx1;
  reg [31:0] rva_out_reg_data_223_192_sva_dfm_3;
  wire [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_223_192_mx1;
  reg [31:0] rva_out_reg_data_191_160_sva_dfm_3;
  wire [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_191_160_mx1;
  reg [31:0] rva_out_reg_data_159_128_sva_dfm_3;
  wire [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_159_128_mx1;
  reg [7:0] rva_out_reg_data_127_120_sva_dfm_3;
  wire [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_127_96_mx1;
  reg [7:0] rva_out_reg_data_119_112_sva_dfm_3;
  reg [7:0] rva_out_reg_data_111_104_sva_dfm_3;
  reg [7:0] rva_out_reg_data_103_96_sva_dfm_3;
  reg [7:0] rva_out_reg_data_95_88_sva_dfm_3;
  wire [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_95_64_mx1;
  reg [7:0] rva_out_reg_data_87_80_sva_dfm_3;
  reg [7:0] rva_out_reg_data_79_72_sva_dfm_3;
  reg [7:0] rva_out_reg_data_71_64_sva_dfm_3;
  reg [7:0] rva_out_reg_data_63_56_sva_dfm_3;
  wire [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_63_32_mx1;
  reg [2:0] rva_out_reg_data_55_53_sva_dfm_3;
  reg [4:0] rva_out_reg_data_52_48_sva_dfm_3;
  reg [7:0] rva_out_reg_data_47_40_sva_dfm_3;
  reg [7:0] rva_out_reg_data_39_32_sva_dfm_3;
  reg [1:0] rva_out_reg_data_31_30_sva_dfm_3;
  wire [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_31_0_mx1;
  reg [5:0] rva_out_reg_data_29_24_sva_dfm_3;
  reg [7:0] rva_out_reg_data_23_16_sva_dfm_3;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_3;
  reg rva_out_reg_data_8_sva_dfm_3;
  reg [6:0] rva_out_reg_data_7_1_sva_dfm_3;
  reg rva_out_reg_data_0_sva_dfm_3;
  wire or_dcpl_639;
  reg [511:0] ActUnit_RunInst_case_3_act_port_reg_data_sva;
  wire act_config_ActConfigRead_else_else_not_21;
  wire [4:0] act_read_addrs_sva_2_mx0w0;
  wire [5:0] nl_act_read_addrs_sva_2_mx0w0;
  reg [4:0] act_config_inst_counter_sva;
  reg [7:0] act_config_output_counter_sva;
  wire or_996_tmp;
  wire mux_205_itm;
  wire mux_215_itm;
  wire mux_229_itm;
  wire mux_231_itm;
  wire mux_234_itm;
  wire mux_235_itm;
  wire and_dcpl_1013;
  wire and_dcpl_1019;
  wire and_dcpl_1021;
  wire and_dcpl_1028;
  wire and_dcpl_1046;
  reg [5:0] act_config_num_inst_sva;
  reg [7:0] act_config_num_output_sva;
  reg [4:0] act_config_buffer_addr_base_sva;
  reg ActUnit_DecodeAxi_rva_in_reg_rw_sva;
  reg ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva;
  reg ActUnit_DecodeAxiWrite_else_unequal_tmp;
  reg ActUnit_DecodeAxiRead_else_unequal_tmp;
  reg [30:0] Relu_for_y_qr_30_0_1_lpi_1_dfm;
  reg [30:0] Relu_for_y_qr_30_0_2_lpi_1_dfm;
  reg [30:0] Relu_for_y_qr_30_0_3_lpi_1_dfm;
  reg [30:0] Relu_for_y_qr_30_0_4_lpi_1_dfm;
  reg [30:0] Relu_for_y_qr_30_0_5_lpi_1_dfm;
  reg [30:0] Relu_for_y_qr_30_0_6_lpi_1_dfm;
  reg [30:0] Relu_for_y_qr_30_0_7_lpi_1_dfm;
  reg [30:0] Relu_for_y_qr_30_0_8_lpi_1_dfm;
  reg [30:0] Relu_for_y_qr_30_0_9_lpi_1_dfm;
  reg [30:0] Relu_for_y_qr_30_0_10_lpi_1_dfm;
  reg [30:0] Relu_for_y_qr_30_0_11_lpi_1_dfm;
  reg [30:0] Relu_for_y_qr_30_0_12_lpi_1_dfm;
  reg [30:0] Relu_for_y_qr_30_0_13_lpi_1_dfm;
  reg [30:0] Relu_for_y_qr_30_0_14_lpi_1_dfm;
  reg [30:0] Relu_for_y_qr_30_0_15_lpi_1_dfm;
  reg [30:0] Relu_for_y_qr_30_0_lpi_1_dfm;
  reg [4:0] act_write_addrs_lpi_1_dfm_5;
  reg [31:0] act_mem_banks_bank_a_0_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_0_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_0_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_0_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_0_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_0_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_0_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_0_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_0_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_0_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_0_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_0_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_0_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_0_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_0_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_0_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_1_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_1_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_1_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_1_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_1_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_1_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_1_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_1_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_1_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_1_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_1_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_1_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_1_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_1_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_1_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_1_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_2_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_2_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_2_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_2_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_2_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_2_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_2_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_2_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_2_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_2_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_2_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_2_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_2_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_2_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_2_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_2_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_3_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_3_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_3_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_3_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_3_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_3_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_3_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_3_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_3_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_3_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_3_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_3_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_3_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_3_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_3_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_3_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_4_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_4_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_4_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_4_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_4_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_4_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_4_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_4_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_4_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_4_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_4_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_4_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_4_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_4_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_4_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_4_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_5_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_5_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_5_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_5_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_5_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_5_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_5_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_5_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_5_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_5_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_5_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_5_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_5_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_5_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_5_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_5_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_6_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_6_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_6_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_6_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_6_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_6_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_6_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_6_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_6_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_6_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_6_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_6_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_6_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_6_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_6_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_6_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_7_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_7_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_7_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_7_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_7_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_7_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_7_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_7_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_7_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_7_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_7_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_7_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_7_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_7_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_7_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_7_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_8_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_8_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_8_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_8_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_8_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_8_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_8_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_8_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_8_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_8_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_8_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_8_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_8_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_8_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_8_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_8_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_9_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_9_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_9_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_9_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_9_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_9_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_9_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_9_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_9_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_9_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_9_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_9_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_9_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_9_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_9_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_9_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_10_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_10_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_10_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_10_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_10_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_10_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_10_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_10_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_10_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_10_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_10_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_10_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_10_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_10_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_10_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_10_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_11_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_11_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_11_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_11_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_11_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_11_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_11_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_11_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_11_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_11_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_11_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_11_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_11_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_11_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_11_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_11_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_12_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_12_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_12_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_12_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_12_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_12_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_12_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_12_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_12_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_12_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_12_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_12_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_12_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_12_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_12_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_12_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_13_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_13_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_13_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_13_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_13_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_13_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_13_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_13_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_13_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_13_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_13_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_13_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_13_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_13_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_13_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_13_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_14_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_14_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_14_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_14_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_14_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_14_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_14_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_14_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_14_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_14_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_14_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_14_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_14_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_14_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_14_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_14_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_15_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_15_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_15_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_15_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_15_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_15_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_15_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_15_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_15_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_15_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_15_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_15_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_15_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_15_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_15_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_15_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_16_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_16_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_16_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_16_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_16_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_16_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_16_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_16_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_16_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_16_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_16_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_16_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_16_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_16_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_16_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_16_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_17_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_17_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_17_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_17_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_17_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_17_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_17_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_17_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_17_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_17_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_17_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_17_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_17_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_17_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_17_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_17_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_18_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_18_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_18_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_18_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_18_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_18_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_18_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_18_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_18_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_18_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_18_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_18_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_18_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_18_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_18_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_18_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_19_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_19_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_19_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_19_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_19_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_19_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_19_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_19_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_19_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_19_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_19_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_19_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_19_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_19_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_19_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_19_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_20_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_20_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_20_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_20_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_20_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_20_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_20_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_20_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_20_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_20_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_20_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_20_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_20_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_20_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_20_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_20_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_21_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_21_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_21_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_21_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_21_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_21_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_21_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_21_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_21_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_21_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_21_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_21_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_21_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_21_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_21_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_21_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_22_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_22_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_22_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_22_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_22_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_22_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_22_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_22_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_22_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_22_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_22_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_22_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_22_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_22_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_22_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_22_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_23_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_23_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_23_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_23_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_23_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_23_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_23_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_23_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_23_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_23_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_23_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_23_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_23_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_23_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_23_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_23_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_24_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_24_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_24_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_24_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_24_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_24_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_24_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_24_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_24_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_24_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_24_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_24_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_24_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_24_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_24_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_24_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_25_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_25_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_25_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_25_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_25_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_25_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_25_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_25_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_25_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_25_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_25_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_25_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_25_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_25_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_25_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_25_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_26_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_26_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_26_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_26_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_26_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_26_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_26_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_26_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_26_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_26_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_26_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_26_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_26_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_26_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_26_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_26_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_27_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_27_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_27_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_27_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_27_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_27_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_27_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_27_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_27_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_27_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_27_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_27_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_27_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_27_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_27_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_27_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_28_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_28_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_28_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_28_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_28_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_28_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_28_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_28_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_28_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_28_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_28_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_28_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_28_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_28_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_28_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_28_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_29_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_29_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_29_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_29_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_29_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_29_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_29_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_29_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_29_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_29_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_29_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_29_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_29_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_29_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_29_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_29_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_30_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_30_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_30_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_30_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_30_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_30_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_30_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_30_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_30_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_30_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_30_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_30_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_30_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_30_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_30_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_30_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_31_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_31_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_31_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_31_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_31_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_31_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_31_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_31_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_31_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_31_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_31_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_31_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_31_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_31_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_31_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_31_31_0_sva_dfm;
  reg [31:0] act_port_read_out_data_0_0_sva_dfm;
  reg [31:0] act_port_read_out_data_0_1_sva_dfm;
  reg [31:0] act_port_read_out_data_0_2_sva_dfm;
  reg [31:0] act_port_read_out_data_0_3_sva_dfm;
  reg [31:0] act_port_read_out_data_0_4_sva_dfm;
  reg [31:0] act_port_read_out_data_0_5_sva_dfm;
  reg [31:0] act_port_read_out_data_0_6_sva_dfm;
  reg [31:0] act_port_read_out_data_0_7_sva_dfm;
  reg [31:0] act_port_read_out_data_0_8_sva_dfm;
  reg [31:0] act_port_read_out_data_0_9_sva_dfm;
  reg [31:0] act_port_read_out_data_0_10_sva_dfm;
  reg [31:0] act_port_read_out_data_0_11_sva_dfm;
  reg [31:0] act_port_read_out_data_0_12_sva_dfm;
  reg [31:0] act_port_read_out_data_0_13_sva_dfm;
  reg [31:0] act_port_read_out_data_0_14_sva_dfm;
  reg [31:0] act_port_read_out_data_0_15_sva_dfm;
  reg [1:0] nvhls_get_slc_2U_NVUINT8_return_2_sva;
  reg act_config_InstIncr_if_act_config_InstIncr_if_if_nor_mdf_sva;
  reg [7:0] rva_out_reg_data_71_64_sva_dfm_6;
  reg [4:0] rva_out_reg_data_52_48_sva_dfm_6;
  reg [7:0] rva_out_reg_data_39_32_sva_dfm_6;
  reg [5:0] rva_out_reg_data_29_24_sva_dfm_6;
  reg [31:0] act_mem_banks_read_for_mux_itm;
  reg [31:0] act_mem_banks_read_for_mux_1_itm;
  reg [31:0] act_mem_banks_read_for_mux_2_itm;
  reg [31:0] act_mem_banks_read_for_mux_3_itm;
  reg [31:0] act_mem_banks_read_for_mux_4_itm;
  reg [31:0] act_mem_banks_read_for_mux_5_itm;
  reg [31:0] act_mem_banks_read_for_mux_6_itm;
  reg [31:0] act_mem_banks_read_for_mux_7_itm;
  reg [31:0] act_mem_banks_read_for_mux_8_itm;
  reg [31:0] act_mem_banks_read_for_mux_9_itm;
  reg [31:0] act_mem_banks_read_for_mux_10_itm;
  reg [31:0] act_mem_banks_read_for_mux_11_itm;
  reg [31:0] act_mem_banks_read_for_mux_12_itm;
  reg [31:0] act_mem_banks_read_for_mux_13_itm;
  reg [31:0] act_mem_banks_read_for_mux_14_itm;
  reg [31:0] act_mem_banks_read_for_mux_15_itm;
  reg while_else_1_mux_1_itm;
  reg [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_511_480;
  reg [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_479_448;
  reg [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_447_416;
  reg [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_415_384;
  reg [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_383_352;
  reg [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_351_320;
  reg [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_319_288;
  reg [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_287_256;
  reg [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_255_224;
  reg [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_223_192;
  reg [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_191_160;
  reg [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_159_128;
  reg [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_127_96;
  reg [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_95_64;
  reg [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_63_32;
  reg [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_31_0;
  reg act_config_inst_regs_16_sva_0;
  reg act_config_inst_regs_17_sva_0;
  reg act_config_inst_regs_1_sva_0;
  reg act_config_inst_regs_0_sva_0;
  wire ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0;
  wire act_config_output_counter_sva_mx0c1;
  wire act_config_inst_counter_sva_mx0c1;
  wire [4:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_2_mx0w2;
  wire ActUnit_PushOutput_if_for_and_stg_2_7_sva_1;
  wire ActUnit_RunInst_switch_lp_equal_tmp_9;
  wire ActUnit_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva_mx0c2;
  wire ActUnit_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva_mx0c3;
  wire ActUnit_CheckStart_if_ActUnit_CheckStart_if_and_itm_1;
  wire ActUnit_PushOutput_if_for_i_4_0_sva_3_0_mx0c0;
  wire act_regs_data_0_0_sva_8_mx3c1;
  wire act_regs_data_0_1_sva_8_mx3c1;
  wire act_regs_data_0_10_sva_8_mx3c1;
  wire act_regs_data_0_11_sva_8_mx3c1;
  wire act_regs_data_0_12_sva_8_mx3c1;
  wire act_regs_data_0_13_sva_8_mx3c1;
  wire act_regs_data_0_14_sva_8_mx3c1;
  wire act_regs_data_0_15_sva_8_mx3c1;
  wire act_regs_data_0_2_sva_8_mx3c1;
  wire act_regs_data_0_3_sva_8_mx3c1;
  wire act_regs_data_0_4_sva_8_mx3c1;
  wire act_regs_data_0_5_sva_8_mx3c1;
  wire act_regs_data_0_6_sva_8_mx3c1;
  wire act_regs_data_0_7_sva_8_mx3c1;
  wire act_regs_data_0_8_sva_8_mx3c1;
  wire [4:0] while_mux_53_ssc_mx0;
  wire [4:0] act_read_addrs_lpi_1_dfm_7;
  wire act_regs_data_3_0_sva_8_mx2c1;
  wire act_regs_data_2_15_sva_8_mx2c1;
  wire act_regs_data_2_14_sva_8_mx2c1;
  wire act_regs_data_2_13_sva_8_mx2c1;
  wire act_regs_data_2_12_sva_8_mx2c1;
  wire act_regs_data_2_11_sva_8_mx2c1;
  wire act_regs_data_2_10_sva_8_mx2c1;
  wire act_regs_data_2_9_sva_8_mx2c1;
  wire act_regs_data_2_8_sva_8_mx2c1;
  wire act_regs_data_2_7_sva_8_mx2c1;
  wire act_regs_data_2_6_sva_8_mx2c1;
  wire act_regs_data_2_5_sva_8_mx2c1;
  wire act_regs_data_2_4_sva_8_mx2c1;
  wire act_regs_data_2_3_sva_8_mx2c1;
  wire act_regs_data_2_2_sva_8_mx2c1;
  wire act_regs_data_2_1_sva_8_mx2c1;
  wire act_regs_data_2_0_sva_8_mx2c1;
  wire act_regs_data_1_15_sva_8_mx2c1;
  wire act_regs_data_1_14_sva_8_mx2c1;
  wire act_regs_data_1_13_sva_8_mx2c1;
  wire act_regs_data_1_12_sva_8_mx2c1;
  wire act_regs_data_1_11_sva_8_mx2c1;
  wire act_regs_data_1_10_sva_8_mx2c1;
  wire act_regs_data_1_9_sva_8_mx2c1;
  wire act_regs_data_1_8_sva_8_mx2c1;
  wire act_regs_data_1_7_sva_8_mx2c1;
  wire act_regs_data_1_6_sva_8_mx2c1;
  wire act_regs_data_1_5_sva_8_mx2c1;
  wire act_regs_data_1_4_sva_8_mx2c1;
  wire act_regs_data_1_3_sva_8_mx2c1;
  wire act_regs_data_1_2_sva_8_mx2c1;
  wire act_regs_data_1_1_sva_8_mx2c1;
  wire act_regs_data_1_0_sva_8_mx2c1;
  wire act_regs_data_0_9_sva_8_mx2c1;
  wire [31:0] act_write_data_data_0_0_lpi_1_dfm_7;
  wire [31:0] act_write_data_data_0_1_lpi_1_dfm_7;
  wire [31:0] act_write_data_data_0_2_lpi_1_dfm_7;
  wire [31:0] act_write_data_data_0_3_lpi_1_dfm_7;
  wire [31:0] act_write_data_data_0_4_lpi_1_dfm_7;
  wire [31:0] act_write_data_data_0_5_lpi_1_dfm_7;
  wire [31:0] act_write_data_data_0_6_lpi_1_dfm_7;
  wire [31:0] act_write_data_data_0_7_lpi_1_dfm_7;
  wire [31:0] act_write_data_data_0_8_lpi_1_dfm_7;
  wire [31:0] act_write_data_data_0_9_lpi_1_dfm_7;
  wire [31:0] act_write_data_data_0_10_lpi_1_dfm_7;
  wire [31:0] act_write_data_data_0_11_lpi_1_dfm_7;
  wire [31:0] act_write_data_data_0_12_lpi_1_dfm_7;
  wire [31:0] act_write_data_data_0_13_lpi_1_dfm_7;
  wire [31:0] act_write_data_data_0_14_lpi_1_dfm_7;
  wire [31:0] act_write_data_data_0_15_lpi_1_dfm_7;
  wire while_asn_1331;
  wire while_asn_1333;
  wire while_asn_1335;
  wire while_asn_1341;
  wire while_asn_1343;
  wire while_asn_1345;
  wire while_asn_1347;
  wire while_asn_1349;
  wire while_asn_1351;
  wire while_asn_1353;
  wire while_asn_1355;
  wire while_asn_1357;
  wire while_asn_1359;
  wire while_asn_1361;
  wire while_asn_1363;
  wire while_asn_1365;
  wire while_asn_1367;
  wire while_asn_1369;
  wire while_asn_1371;
  wire while_asn_1373;
  wire while_asn_1375;
  wire while_asn_1377;
  wire while_asn_1379;
  wire while_asn_1381;
  wire while_asn_1383;
  wire while_asn_1385;
  wire while_asn_1387;
  wire while_asn_1389;
  wire while_asn_1391;
  wire while_asn_1393;
  wire while_asn_1395;
  wire [31:0] ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1;
  wire while_asn_1397;
  wire while_asn_1399;
  wire while_asn_1401;
  reg [30:0] ActUnit_RunInst_case_14_nv_scvector_cctor_data_0_sva_30_0;
  reg [30:0] nv_scvector_cctor_nv_scvector_5_for_2_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_65_0;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_67_0;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_69_0;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_71_0;
  wire [30:0] Tanh_for_16_exs_5_30_0;
  wire [30:0] Tanh_for_15_exs_5_30_0;
  wire [30:0] Tanh_for_14_exs_5_30_0;
  wire [30:0] Tanh_for_13_exs_5_30_0;
  wire [30:0] Tanh_for_12_exs_5_30_0;
  wire [30:0] Tanh_for_11_exs_5_30_0;
  wire [30:0] Tanh_for_10_exs_5_30_0;
  wire [30:0] Tanh_for_9_exs_5_30_0;
  wire [30:0] Tanh_for_8_exs_5_30_0;
  wire [30:0] Tanh_for_7_exs_5_30_0;
  wire [30:0] Tanh_for_6_exs_5_30_0;
  wire [30:0] Tanh_for_5_exs_5_30_0;
  wire [30:0] Tanh_for_4_exs_5_30_0;
  wire [30:0] Tanh_for_3_exs_5_30_0;
  wire [30:0] Tanh_for_2_exs_5_30_0;
  wire [30:0] Tanh_for_1_exs_5_30_0;
  wire Gelu_for_y_lpi_1_dfm_2_31;
  wire [30:0] Gelu_for_y_lpi_1_dfm_2_30_0;
  wire Gelu_for_y_11_lpi_1_dfm_2_31;
  wire [30:0] Gelu_for_y_11_lpi_1_dfm_2_30_0;
  wire Gelu_for_y_10_lpi_1_dfm_2_31;
  wire [30:0] Gelu_for_y_10_lpi_1_dfm_2_30_0;
  wire ActUnit_PushOutput_if_for_and_28_cse;
  wire Silu_for_y_and_7_cse;
  wire and_1152_cse;
  wire and_1156_cse;
  wire and_1158_cse;
  wire and_1161_cse;
  wire and_1154_cse;
  wire and_1181_cse;
  wire and_1183_cse;
  wire and_1185_cse;
  wire and_1190_cse;
  wire and_1191_cse;
  wire nv_scvector_cctor_nv_scvector_5_for_and_cse;
  wire ActUnit_RunInst_switch_lp_and_812_cse;
  wire nv_scvector_cctor_nv_scvector_5_for_and_3_cse;
  wire nv_scvector_cctor_nv_scvector_5_for_and_5_cse;
  wire nv_scvector_cctor_nv_scvector_5_for_and_7_cse;
  wire nv_scvector_cctor_nv_scvector_5_for_and_9_cse;
  wire nv_scvector_cctor_nv_scvector_5_for_and_11_cse;
  wire nv_scvector_cctor_nv_scvector_5_for_and_13_cse;
  wire nv_scvector_cctor_nv_scvector_6_for_and_7_cse;
  reg ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_31;
  reg [30:0] ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_30_0;
  reg ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_31;
  reg [30:0] ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_30_0;
  reg ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_31;
  reg [30:0] ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_30_0;
  reg ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_31;
  reg [30:0] ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_30_0;
  reg ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_31;
  reg [30:0] ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_30_0;
  reg ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_31;
  reg [30:0] ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_30_0;
  reg ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_31;
  reg [30:0] ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_30_0;
  reg ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_31;
  reg [30:0] ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_30_0;
  reg ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_31;
  reg [30:0] ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_30_0;
  reg ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_31;
  reg [30:0] ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_30_0;
  reg ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_31;
  reg [30:0] ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_30_0;
  reg ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_31;
  reg [30:0] ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_30_0;
  reg ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_31;
  reg [30:0] ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_30_0;
  reg ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_31;
  reg [30:0] ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_30_0;
  reg ActUnit_PushOutput_if_output_port_reg_data_data_1_sva_31;
  reg [30:0] ActUnit_PushOutput_if_output_port_reg_data_data_1_sva_30_0;
  wire ActUnit_RunInst_case_2_for_and_27_seb;
  reg ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_31;
  reg [30:0] ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_30_0;
  wire Silu_for_y_and_ssc;
  reg Silu_for_y_2_lpi_1_dfm_1_31;
  reg [30:0] Silu_for_y_2_lpi_1_dfm_1_30_0;
  reg Silu_for_y_3_lpi_1_dfm_1_31;
  reg [30:0] Silu_for_y_3_lpi_1_dfm_1_30_0;
  wire Silu_for_y_and_13_ssc;
  reg Silu_for_y_4_lpi_1_dfm_1_31;
  reg [30:0] Silu_for_y_4_lpi_1_dfm_1_30_0;
  reg Silu_for_y_5_lpi_1_dfm_1_31;
  reg [30:0] Silu_for_y_5_lpi_1_dfm_1_30_0;
  wire Silu_for_y_and_15_ssc;
  reg Silu_for_y_6_lpi_1_dfm_1_31;
  reg [30:0] Silu_for_y_6_lpi_1_dfm_1_30_0;
  reg Silu_for_y_7_lpi_1_dfm_1_31;
  reg [30:0] Silu_for_y_7_lpi_1_dfm_1_30_0;
  wire Silu_for_y_and_17_ssc;
  reg Silu_for_y_8_lpi_1_dfm_1_31;
  reg [30:0] Silu_for_y_8_lpi_1_dfm_1_30_0;
  wire Silu_for_y_and_19_ssc;
  reg Silu_for_y_9_lpi_1_dfm_1_31;
  reg [30:0] Silu_for_y_9_lpi_1_dfm_1_30_0;
  wire Silu_for_y_and_8_ssc;
  reg Silu_for_y_12_lpi_1_dfm_1_31;
  reg [30:0] Silu_for_y_12_lpi_1_dfm_1_30_0;
  reg Silu_for_y_13_lpi_1_dfm_1_31;
  reg [30:0] Silu_for_y_13_lpi_1_dfm_1_30_0;
  wire Silu_for_y_and_20_ssc;
  reg Silu_for_y_14_lpi_1_dfm_1_31;
  reg [30:0] Silu_for_y_14_lpi_1_dfm_1_30_0;
  reg Silu_for_y_15_lpi_1_dfm_1_31;
  reg [30:0] Silu_for_y_15_lpi_1_dfm_1_30_0;
  wire Silu_for_y_and_22_ssc;
  reg Silu_for_y_lpi_1_dfm_1_31;
  reg [30:0] Silu_for_y_lpi_1_dfm_1_30_0;
  reg act_regs_data_0_15_sva_31;
  reg [30:0] act_regs_data_0_15_sva_30_0;
  reg act_regs_data_0_14_sva_31;
  reg [30:0] act_regs_data_0_14_sva_30_0;
  reg act_regs_data_0_13_sva_31;
  reg [30:0] act_regs_data_0_13_sva_30_0;
  reg act_regs_data_0_12_sva_31;
  reg [30:0] act_regs_data_0_12_sva_30_0;
  reg act_regs_data_0_11_sva_31;
  reg [30:0] act_regs_data_0_11_sva_30_0;
  reg act_regs_data_0_10_sva_31;
  reg [30:0] act_regs_data_0_10_sva_30_0;
  reg act_regs_data_0_8_sva_31;
  reg [30:0] act_regs_data_0_8_sva_30_0;
  reg act_regs_data_0_7_sva_31;
  reg [30:0] act_regs_data_0_7_sva_30_0;
  reg act_regs_data_0_6_sva_31;
  reg [30:0] act_regs_data_0_6_sva_30_0;
  reg act_regs_data_0_5_sva_31;
  reg [30:0] act_regs_data_0_5_sva_30_0;
  reg act_regs_data_0_4_sva_31;
  reg [30:0] act_regs_data_0_4_sva_30_0;
  reg act_regs_data_0_3_sva_31;
  reg [30:0] act_regs_data_0_3_sva_30_0;
  reg act_regs_data_0_2_sva_31;
  reg [30:0] act_regs_data_0_2_sva_30_0;
  reg act_regs_data_0_1_sva_31;
  reg [30:0] act_regs_data_0_1_sva_30_0;
  reg act_regs_data_0_0_sva_31;
  reg [30:0] act_regs_data_0_0_sva_30_0;
  reg act_regs_data_0_0_sva_dfm_2_31;
  reg [30:0] act_regs_data_0_0_sva_dfm_2_30_0;
  reg act_regs_data_0_1_sva_dfm_2_31;
  reg [30:0] act_regs_data_0_1_sva_dfm_2_30_0;
  reg act_regs_data_0_2_sva_dfm_2_31;
  reg [30:0] act_regs_data_0_2_sva_dfm_2_30_0;
  reg act_regs_data_0_3_sva_dfm_2_31;
  reg [30:0] act_regs_data_0_3_sva_dfm_2_30_0;
  reg act_regs_data_0_4_sva_dfm_2_31;
  reg [30:0] act_regs_data_0_4_sva_dfm_2_30_0;
  reg act_regs_data_0_5_sva_dfm_2_31;
  reg [30:0] act_regs_data_0_5_sva_dfm_2_30_0;
  reg act_regs_data_0_6_sva_dfm_2_31;
  reg [30:0] act_regs_data_0_6_sva_dfm_2_30_0;
  reg act_regs_data_0_7_sva_dfm_2_31;
  reg [30:0] act_regs_data_0_7_sva_dfm_2_30_0;
  reg act_regs_data_0_8_sva_dfm_2_31;
  reg [30:0] act_regs_data_0_8_sva_dfm_2_30_0;
  reg act_regs_data_0_10_sva_dfm_2_31;
  reg [30:0] act_regs_data_0_10_sva_dfm_2_30_0;
  reg act_regs_data_0_11_sva_dfm_2_31;
  reg [30:0] act_regs_data_0_11_sva_dfm_2_30_0;
  reg act_regs_data_0_12_sva_dfm_2_31;
  reg [30:0] act_regs_data_0_12_sva_dfm_2_30_0;
  reg act_regs_data_0_13_sva_dfm_2_31;
  reg [30:0] act_regs_data_0_13_sva_dfm_2_30_0;
  reg act_regs_data_0_14_sva_dfm_2_31;
  reg [30:0] act_regs_data_0_14_sva_dfm_2_30_0;
  reg act_regs_data_0_15_sva_dfm_2_31;
  reg [30:0] act_regs_data_0_15_sva_dfm_2_30_0;
  wire Tanh_for_else_else_and_2_cse;
  wire Tanh_for_else_else_and_3_cse;
  wire Tanh_for_else_else_or_cse;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31;
  reg [30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31;
  reg [30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31;
  reg [30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31;
  reg [30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31;
  reg [30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31;
  reg [30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31;
  reg [30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31;
  reg [30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31;
  reg [30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31;
  reg [30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31;
  reg [30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31;
  reg [30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31;
  reg [30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31;
  reg [30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31;
  reg [30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0;
  wire act_regs_data_and_418_ssc;
  wire act_regs_data_and_419_ssc;
  wire act_regs_data_and_71_ssc;
  reg act_regs_data_0_15_sva_8_31;
  reg [30:0] act_regs_data_0_15_sva_8_30_0;
  wire act_regs_data_and_416_ssc;
  wire act_regs_data_and_417_ssc;
  wire act_regs_data_and_70_ssc;
  reg act_regs_data_0_14_sva_8_31;
  reg [30:0] act_regs_data_0_14_sva_8_30_0;
  wire act_regs_data_and_414_ssc;
  wire act_regs_data_and_415_ssc;
  wire act_regs_data_and_69_ssc;
  reg act_regs_data_0_13_sva_8_31;
  reg [30:0] act_regs_data_0_13_sva_8_30_0;
  wire act_regs_data_and_412_ssc;
  wire act_regs_data_and_413_ssc;
  wire act_regs_data_and_68_ssc;
  reg act_regs_data_0_12_sva_8_31;
  reg [30:0] act_regs_data_0_12_sva_8_30_0;
  wire act_regs_data_and_410_ssc;
  wire act_regs_data_and_411_ssc;
  wire act_regs_data_and_67_ssc;
  reg act_regs_data_0_11_sva_8_31;
  reg [30:0] act_regs_data_0_11_sva_8_30_0;
  wire act_regs_data_and_408_ssc;
  wire act_regs_data_and_409_ssc;
  wire act_regs_data_and_66_ssc;
  reg act_regs_data_0_10_sva_8_31;
  reg [30:0] act_regs_data_0_10_sva_8_30_0;
  wire act_regs_data_and_432_ssc;
  wire act_regs_data_and_433_ssc;
  wire act_regs_data_and_78_ssc;
  reg act_regs_data_0_8_sva_8_31;
  reg [30:0] act_regs_data_0_8_sva_8_30_0;
  wire act_regs_data_and_430_ssc;
  wire act_regs_data_and_431_ssc;
  wire act_regs_data_and_77_ssc;
  reg act_regs_data_0_7_sva_8_31;
  reg [30:0] act_regs_data_0_7_sva_8_30_0;
  wire act_regs_data_and_428_ssc;
  wire act_regs_data_and_429_ssc;
  wire act_regs_data_and_76_ssc;
  reg act_regs_data_0_6_sva_8_31;
  reg [30:0] act_regs_data_0_6_sva_8_30_0;
  wire act_regs_data_and_426_ssc;
  wire act_regs_data_and_427_ssc;
  wire act_regs_data_and_75_ssc;
  reg act_regs_data_0_5_sva_8_31;
  reg [30:0] act_regs_data_0_5_sva_8_30_0;
  wire act_regs_data_and_424_ssc;
  wire act_regs_data_and_425_ssc;
  wire act_regs_data_and_74_ssc;
  reg act_regs_data_0_4_sva_8_31;
  reg [30:0] act_regs_data_0_4_sva_8_30_0;
  wire act_regs_data_and_422_ssc;
  wire act_regs_data_and_423_ssc;
  wire act_regs_data_and_73_ssc;
  reg act_regs_data_0_3_sva_8_31;
  reg [30:0] act_regs_data_0_3_sva_8_30_0;
  wire act_regs_data_and_420_ssc;
  wire act_regs_data_and_421_ssc;
  wire act_regs_data_and_72_ssc;
  reg act_regs_data_0_2_sva_8_31;
  reg [30:0] act_regs_data_0_2_sva_8_30_0;
  wire act_regs_data_and_406_ssc;
  wire act_regs_data_and_407_ssc;
  wire act_regs_data_and_65_ssc;
  reg act_regs_data_0_1_sva_8_31;
  reg [30:0] act_regs_data_0_1_sva_8_30_0;
  wire act_regs_data_and_404_ssc;
  wire act_regs_data_and_405_ssc;
  wire act_regs_data_and_64_ssc;
  reg act_regs_data_0_0_sva_8_31;
  reg [30:0] act_regs_data_0_0_sva_8_30_0;
  wire ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_31;
  wire [30:0] ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_30_0;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_2_31;
  wire [30:0] ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_2_30_0;
  reg act_regs_data_1_15_sva_31;
  reg [30:0] act_regs_data_1_15_sva_30_0;
  reg act_regs_data_1_14_sva_31;
  reg [30:0] act_regs_data_1_14_sva_30_0;
  reg act_regs_data_1_13_sva_31;
  reg [30:0] act_regs_data_1_13_sva_30_0;
  reg act_regs_data_1_12_sva_31;
  reg [30:0] act_regs_data_1_12_sva_30_0;
  reg act_regs_data_1_11_sva_31;
  reg [30:0] act_regs_data_1_11_sva_30_0;
  reg act_regs_data_1_10_sva_31;
  reg [30:0] act_regs_data_1_10_sva_30_0;
  reg act_regs_data_1_7_sva_31;
  reg [30:0] act_regs_data_1_7_sva_30_0;
  reg act_regs_data_1_6_sva_31;
  reg [30:0] act_regs_data_1_6_sva_30_0;
  reg act_regs_data_1_5_sva_31;
  reg [30:0] act_regs_data_1_5_sva_30_0;
  reg act_regs_data_1_4_sva_31;
  reg [30:0] act_regs_data_1_4_sva_30_0;
  reg act_regs_data_1_3_sva_31;
  reg [30:0] act_regs_data_1_3_sva_30_0;
  reg act_regs_data_1_2_sva_31;
  reg [30:0] act_regs_data_1_2_sva_30_0;
  reg act_regs_data_1_1_sva_31;
  reg [30:0] act_regs_data_1_1_sva_30_0;
  reg act_regs_data_1_0_sva_31;
  reg [30:0] act_regs_data_1_0_sva_30_0;
  reg act_regs_data_0_9_sva_31;
  reg [30:0] act_regs_data_0_9_sva_30_0;
  reg act_regs_data_0_9_sva_dfm_2_31;
  reg [30:0] act_regs_data_0_9_sva_dfm_2_30_0;
  reg act_regs_data_1_0_sva_dfm_2_31;
  reg [30:0] act_regs_data_1_0_sva_dfm_2_30_0;
  reg act_regs_data_1_1_sva_dfm_2_31;
  reg [30:0] act_regs_data_1_1_sva_dfm_2_30_0;
  reg act_regs_data_1_2_sva_dfm_2_31;
  reg [30:0] act_regs_data_1_2_sva_dfm_2_30_0;
  reg act_regs_data_1_3_sva_dfm_2_31;
  reg [30:0] act_regs_data_1_3_sva_dfm_2_30_0;
  reg act_regs_data_1_4_sva_dfm_2_31;
  reg [30:0] act_regs_data_1_4_sva_dfm_2_30_0;
  reg act_regs_data_1_5_sva_dfm_2_31;
  reg [30:0] act_regs_data_1_5_sva_dfm_2_30_0;
  reg act_regs_data_1_6_sva_dfm_2_31;
  reg [30:0] act_regs_data_1_6_sva_dfm_2_30_0;
  reg act_regs_data_1_7_sva_dfm_2_31;
  reg [30:0] act_regs_data_1_7_sva_dfm_2_30_0;
  reg act_regs_data_1_8_sva_dfm_2_31;
  reg [30:0] act_regs_data_1_8_sva_dfm_2_30_0;
  reg act_regs_data_1_9_sva_dfm_2_31;
  reg [30:0] act_regs_data_1_9_sva_dfm_2_30_0;
  reg act_regs_data_1_10_sva_dfm_2_31;
  reg [30:0] act_regs_data_1_10_sva_dfm_2_30_0;
  reg act_regs_data_1_11_sva_dfm_2_31;
  reg [30:0] act_regs_data_1_11_sva_dfm_2_30_0;
  reg act_regs_data_1_12_sva_dfm_2_31;
  reg [30:0] act_regs_data_1_12_sva_dfm_2_30_0;
  reg act_regs_data_1_13_sva_dfm_2_31;
  reg [30:0] act_regs_data_1_13_sva_dfm_2_30_0;
  reg act_regs_data_1_14_sva_dfm_2_31;
  reg [30:0] act_regs_data_1_14_sva_dfm_2_30_0;
  reg act_regs_data_1_15_sva_dfm_2_31;
  reg [30:0] act_regs_data_1_15_sva_dfm_2_30_0;
  reg act_regs_data_2_0_sva_dfm_2_31;
  reg [30:0] act_regs_data_2_0_sva_dfm_2_30_0;
  reg act_regs_data_2_1_sva_dfm_2_31;
  reg [30:0] act_regs_data_2_1_sva_dfm_2_30_0;
  reg act_regs_data_2_2_sva_dfm_2_31;
  reg [30:0] act_regs_data_2_2_sva_dfm_2_30_0;
  reg act_regs_data_2_3_sva_dfm_2_31;
  reg [30:0] act_regs_data_2_3_sva_dfm_2_30_0;
  reg act_regs_data_2_4_sva_dfm_2_31;
  reg [30:0] act_regs_data_2_4_sva_dfm_2_30_0;
  reg act_regs_data_2_5_sva_dfm_2_31;
  reg [30:0] act_regs_data_2_5_sva_dfm_2_30_0;
  reg act_regs_data_2_6_sva_dfm_2_31;
  reg [30:0] act_regs_data_2_6_sva_dfm_2_30_0;
  reg act_regs_data_2_7_sva_dfm_2_31;
  reg [30:0] act_regs_data_2_7_sva_dfm_2_30_0;
  reg act_regs_data_2_8_sva_dfm_2_31;
  reg [30:0] act_regs_data_2_8_sva_dfm_2_30_0;
  reg act_regs_data_2_9_sva_dfm_2_31;
  reg [30:0] act_regs_data_2_9_sva_dfm_2_30_0;
  reg act_regs_data_2_10_sva_dfm_2_31;
  reg [30:0] act_regs_data_2_10_sva_dfm_2_30_0;
  reg act_regs_data_2_11_sva_dfm_2_31;
  reg [30:0] act_regs_data_2_11_sva_dfm_2_30_0;
  reg act_regs_data_2_12_sva_dfm_2_31;
  reg [30:0] act_regs_data_2_12_sva_dfm_2_30_0;
  reg act_regs_data_2_13_sva_dfm_2_31;
  reg [30:0] act_regs_data_2_13_sva_dfm_2_30_0;
  reg act_regs_data_2_14_sva_dfm_2_31;
  reg [30:0] act_regs_data_2_14_sva_dfm_2_30_0;
  reg act_regs_data_2_15_sva_dfm_2_31;
  reg [30:0] act_regs_data_2_15_sva_dfm_2_30_0;
  reg act_regs_data_3_0_sva_dfm_2_31;
  reg [30:0] act_regs_data_3_0_sva_dfm_2_30_0;
  reg act_regs_data_3_1_sva_dfm_2_31;
  reg [30:0] act_regs_data_3_1_sva_dfm_2_30_0;
  reg act_regs_data_3_2_sva_dfm_2_31;
  reg [30:0] act_regs_data_3_2_sva_dfm_2_30_0;
  reg act_regs_data_3_3_sva_dfm_2_31;
  reg [30:0] act_regs_data_3_3_sva_dfm_2_30_0;
  reg act_regs_data_3_4_sva_dfm_2_31;
  reg [30:0] act_regs_data_3_4_sva_dfm_2_30_0;
  reg act_regs_data_3_5_sva_dfm_2_31;
  reg [30:0] act_regs_data_3_5_sva_dfm_2_30_0;
  reg act_regs_data_3_6_sva_dfm_2_31;
  reg [30:0] act_regs_data_3_6_sva_dfm_2_30_0;
  reg act_regs_data_3_7_sva_dfm_2_31;
  reg [30:0] act_regs_data_3_7_sva_dfm_2_30_0;
  reg act_regs_data_3_8_sva_dfm_2_31;
  reg [30:0] act_regs_data_3_8_sva_dfm_2_30_0;
  reg act_regs_data_3_9_sva_dfm_2_31;
  reg [30:0] act_regs_data_3_9_sva_dfm_2_30_0;
  reg act_regs_data_3_10_sva_dfm_2_31;
  reg [30:0] act_regs_data_3_10_sva_dfm_2_30_0;
  reg act_regs_data_3_11_sva_dfm_2_31;
  reg [30:0] act_regs_data_3_11_sva_dfm_2_30_0;
  reg act_regs_data_3_12_sva_dfm_2_31;
  reg [30:0] act_regs_data_3_12_sva_dfm_2_30_0;
  reg act_regs_data_3_13_sva_dfm_2_31;
  reg [30:0] act_regs_data_3_13_sva_dfm_2_30_0;
  reg act_regs_data_3_14_sva_dfm_2_31;
  reg [30:0] act_regs_data_3_14_sva_dfm_2_30_0;
  reg act_regs_data_3_15_sva_dfm_2_31;
  reg [30:0] act_regs_data_3_15_sva_dfm_2_30_0;
  wire ActUnit_DecodeAxi_if_and_37_cse;
  wire act_config_inst_regs_and_36_cse;
  wire Relu_for_y_qelse_and_cse;
  wire operator_32_8_true_AC_TRN_AC_WRAP_and_cse;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_and_cse;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_and_17_cse;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_and_19_cse;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_and_21_cse;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_and_23_cse;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_and_25_cse;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_and_27_cse;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_and_29_cse;
  wire act_mem_banks_read_for_and_cse;
  wire rva_out_reg_data_and_62_cse;
  wire act_regs_data_and_284_cse;
  wire nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31;
  wire [30:0] nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
  wire nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31;
  wire [30:0] nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
  wire nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31;
  wire [30:0] nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
  wire nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31;
  wire [30:0] nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
  wire nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31;
  wire [30:0] nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
  wire nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31;
  wire [30:0] nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
  wire nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31;
  wire [30:0] nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
  wire nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31;
  wire [30:0] nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
  wire nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31;
  wire [30:0] nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
  wire nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31;
  wire [30:0] nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
  wire nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31;
  wire [30:0] nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
  wire nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31;
  wire [30:0] nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
  wire nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31;
  wire [30:0] nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
  wire ActUnit_RunInst_case_11_nv_scvector_cctor_data_0_sva_1_31;
  wire [30:0] ActUnit_RunInst_case_11_nv_scvector_cctor_data_0_sva_1_30_0;
  reg act_regs_data_2_0_sva_31;
  reg [30:0] act_regs_data_2_0_sva_30_0;
  reg act_regs_data_2_1_sva_31;
  reg [30:0] act_regs_data_2_1_sva_30_0;
  reg act_regs_data_2_2_sva_31;
  reg [30:0] act_regs_data_2_2_sva_30_0;
  reg act_regs_data_2_3_sva_31;
  reg [30:0] act_regs_data_2_3_sva_30_0;
  reg act_regs_data_2_4_sva_31;
  reg [30:0] act_regs_data_2_4_sva_30_0;
  reg act_regs_data_2_5_sva_31;
  reg [30:0] act_regs_data_2_5_sva_30_0;
  reg act_regs_data_1_9_sva_31;
  reg [30:0] act_regs_data_1_9_sva_30_0;
  reg act_regs_data_2_6_sva_31;
  reg [30:0] act_regs_data_2_6_sva_30_0;
  reg act_regs_data_1_8_sva_31;
  reg [30:0] act_regs_data_1_8_sva_30_0;
  reg act_regs_data_2_7_sva_31;
  reg [30:0] act_regs_data_2_7_sva_30_0;
  reg act_regs_data_2_8_sva_31;
  reg [30:0] act_regs_data_2_8_sva_30_0;
  reg act_regs_data_2_9_sva_31;
  reg [30:0] act_regs_data_2_9_sva_30_0;
  reg act_regs_data_2_10_sva_31;
  reg [30:0] act_regs_data_2_10_sva_30_0;
  reg act_regs_data_2_11_sva_31;
  reg [30:0] act_regs_data_2_11_sva_30_0;
  reg act_regs_data_2_12_sva_31;
  reg [30:0] act_regs_data_2_12_sva_30_0;
  reg act_regs_data_2_13_sva_31;
  reg [30:0] act_regs_data_2_13_sva_30_0;
  reg act_regs_data_2_14_sva_31;
  reg [30:0] act_regs_data_2_14_sva_30_0;
  reg act_regs_data_2_15_sva_31;
  reg [30:0] act_regs_data_2_15_sva_30_0;
  reg act_regs_data_3_0_sva_31;
  reg [30:0] act_regs_data_3_0_sva_30_0;
  reg act_regs_data_3_1_sva_31;
  reg [30:0] act_regs_data_3_1_sva_30_0;
  reg act_regs_data_3_2_sva_31;
  reg [30:0] act_regs_data_3_2_sva_30_0;
  reg act_regs_data_3_3_sva_31;
  reg [30:0] act_regs_data_3_3_sva_30_0;
  reg act_regs_data_3_4_sva_31;
  reg [30:0] act_regs_data_3_4_sva_30_0;
  reg act_regs_data_3_5_sva_31;
  reg [30:0] act_regs_data_3_5_sva_30_0;
  reg act_regs_data_3_6_sva_31;
  reg [30:0] act_regs_data_3_6_sva_30_0;
  reg act_regs_data_3_7_sva_31;
  reg [30:0] act_regs_data_3_7_sva_30_0;
  reg act_regs_data_3_8_sva_31;
  reg [30:0] act_regs_data_3_8_sva_30_0;
  reg act_regs_data_3_9_sva_31;
  reg [30:0] act_regs_data_3_9_sva_30_0;
  reg act_regs_data_3_10_sva_31;
  reg [30:0] act_regs_data_3_10_sva_30_0;
  reg act_regs_data_3_11_sva_31;
  reg [30:0] act_regs_data_3_11_sva_30_0;
  reg act_regs_data_3_12_sva_31;
  reg [30:0] act_regs_data_3_12_sva_30_0;
  reg act_regs_data_3_13_sva_31;
  reg [30:0] act_regs_data_3_13_sva_30_0;
  reg act_regs_data_3_14_sva_31;
  reg [30:0] act_regs_data_3_14_sva_30_0;
  reg act_regs_data_3_15_sva_31;
  reg [30:0] act_regs_data_3_15_sva_30_0;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31;
  reg [30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0;
  wire act_regs_data_and_468_ssc;
  wire act_regs_data_and_469_ssc;
  wire act_regs_data_and_111_ssc;
  reg act_regs_data_1_15_sva_8_31;
  reg [30:0] act_regs_data_1_15_sva_8_30_0;
  wire act_regs_data_and_466_ssc;
  wire act_regs_data_and_467_ssc;
  wire act_regs_data_and_110_ssc;
  reg act_regs_data_2_0_sva_8_31;
  reg [30:0] act_regs_data_2_0_sva_8_30_0;
  wire act_regs_data_and_470_ssc;
  wire act_regs_data_and_471_ssc;
  wire act_regs_data_and_112_ssc;
  reg act_regs_data_1_14_sva_8_31;
  reg [30:0] act_regs_data_1_14_sva_8_30_0;
  wire act_regs_data_and_464_ssc;
  wire act_regs_data_and_465_ssc;
  wire act_regs_data_and_109_ssc;
  reg act_regs_data_2_1_sva_8_31;
  reg [30:0] act_regs_data_2_1_sva_8_30_0;
  wire act_regs_data_and_472_ssc;
  wire act_regs_data_and_473_ssc;
  wire act_regs_data_and_113_ssc;
  reg act_regs_data_1_13_sva_8_31;
  reg [30:0] act_regs_data_1_13_sva_8_30_0;
  wire act_regs_data_and_462_ssc;
  wire act_regs_data_and_463_ssc;
  wire act_regs_data_and_108_ssc;
  reg act_regs_data_2_2_sva_8_31;
  reg [30:0] act_regs_data_2_2_sva_8_30_0;
  wire act_regs_data_and_474_ssc;
  wire act_regs_data_and_475_ssc;
  wire act_regs_data_and_114_ssc;
  reg act_regs_data_1_12_sva_8_31;
  reg [30:0] act_regs_data_1_12_sva_8_30_0;
  wire act_regs_data_and_460_ssc;
  wire act_regs_data_and_461_ssc;
  wire act_regs_data_and_107_ssc;
  reg act_regs_data_2_3_sva_8_31;
  reg [30:0] act_regs_data_2_3_sva_8_30_0;
  wire act_regs_data_and_476_ssc;
  wire act_regs_data_and_477_ssc;
  wire act_regs_data_and_115_ssc;
  reg act_regs_data_1_11_sva_8_31;
  reg [30:0] act_regs_data_1_11_sva_8_30_0;
  wire act_regs_data_and_458_ssc;
  wire act_regs_data_and_459_ssc;
  wire act_regs_data_and_106_ssc;
  reg act_regs_data_2_4_sva_8_31;
  reg [30:0] act_regs_data_2_4_sva_8_30_0;
  wire act_regs_data_and_478_ssc;
  wire act_regs_data_and_479_ssc;
  wire act_regs_data_and_116_ssc;
  reg act_regs_data_1_10_sva_8_31;
  reg [30:0] act_regs_data_1_10_sva_8_30_0;
  wire act_regs_data_and_456_ssc;
  wire act_regs_data_and_457_ssc;
  wire act_regs_data_and_105_ssc;
  reg act_regs_data_2_5_sva_8_31;
  reg [30:0] act_regs_data_2_5_sva_8_30_0;
  wire act_regs_data_and_480_ssc;
  wire act_regs_data_and_481_ssc;
  wire act_regs_data_and_117_ssc;
  reg act_regs_data_1_9_sva_8_31;
  reg [30:0] act_regs_data_1_9_sva_8_30_0;
  wire act_regs_data_and_454_ssc;
  wire act_regs_data_and_455_ssc;
  wire act_regs_data_and_104_ssc;
  reg act_regs_data_2_6_sva_8_31;
  reg [30:0] act_regs_data_2_6_sva_8_30_0;
  wire act_regs_data_and_482_ssc;
  wire act_regs_data_and_483_ssc;
  wire act_regs_data_and_118_ssc;
  reg act_regs_data_1_8_sva_8_31;
  reg [30:0] act_regs_data_1_8_sva_8_30_0;
  wire act_regs_data_and_452_ssc;
  wire act_regs_data_and_453_ssc;
  wire act_regs_data_and_103_ssc;
  reg act_regs_data_2_7_sva_8_31;
  reg [30:0] act_regs_data_2_7_sva_8_30_0;
  wire act_regs_data_and_484_ssc;
  wire act_regs_data_and_485_ssc;
  wire act_regs_data_and_119_ssc;
  reg act_regs_data_1_7_sva_8_31;
  reg [30:0] act_regs_data_1_7_sva_8_30_0;
  wire act_regs_data_and_450_ssc;
  wire act_regs_data_and_451_ssc;
  wire act_regs_data_and_102_ssc;
  reg act_regs_data_2_8_sva_8_31;
  reg [30:0] act_regs_data_2_8_sva_8_30_0;
  wire act_regs_data_and_486_ssc;
  wire act_regs_data_and_487_ssc;
  wire act_regs_data_and_120_ssc;
  reg act_regs_data_1_6_sva_8_31;
  reg [30:0] act_regs_data_1_6_sva_8_30_0;
  wire act_regs_data_and_448_ssc;
  wire act_regs_data_and_449_ssc;
  wire act_regs_data_and_101_ssc;
  reg act_regs_data_2_9_sva_8_31;
  reg [30:0] act_regs_data_2_9_sva_8_30_0;
  wire act_regs_data_and_488_ssc;
  wire act_regs_data_and_489_ssc;
  wire act_regs_data_and_121_ssc;
  reg act_regs_data_1_5_sva_8_31;
  reg [30:0] act_regs_data_1_5_sva_8_30_0;
  wire act_regs_data_and_446_ssc;
  wire act_regs_data_and_447_ssc;
  wire act_regs_data_and_100_ssc;
  reg act_regs_data_2_10_sva_8_31;
  reg [30:0] act_regs_data_2_10_sva_8_30_0;
  wire act_regs_data_and_490_ssc;
  wire act_regs_data_and_491_ssc;
  wire act_regs_data_and_122_ssc;
  reg act_regs_data_1_4_sva_8_31;
  reg [30:0] act_regs_data_1_4_sva_8_30_0;
  wire act_regs_data_and_444_ssc;
  wire act_regs_data_and_445_ssc;
  wire act_regs_data_and_99_ssc;
  reg act_regs_data_2_11_sva_8_31;
  reg [30:0] act_regs_data_2_11_sva_8_30_0;
  wire act_regs_data_and_492_ssc;
  wire act_regs_data_and_493_ssc;
  wire act_regs_data_and_123_ssc;
  reg act_regs_data_1_3_sva_8_31;
  reg [30:0] act_regs_data_1_3_sva_8_30_0;
  wire act_regs_data_and_442_ssc;
  wire act_regs_data_and_443_ssc;
  wire act_regs_data_and_98_ssc;
  reg act_regs_data_2_12_sva_8_31;
  reg [30:0] act_regs_data_2_12_sva_8_30_0;
  wire act_regs_data_and_494_ssc;
  wire act_regs_data_and_495_ssc;
  wire act_regs_data_and_124_ssc;
  reg act_regs_data_1_2_sva_8_31;
  reg [30:0] act_regs_data_1_2_sva_8_30_0;
  wire act_regs_data_and_440_ssc;
  wire act_regs_data_and_441_ssc;
  wire act_regs_data_and_97_ssc;
  reg act_regs_data_2_13_sva_8_31;
  reg [30:0] act_regs_data_2_13_sva_8_30_0;
  wire act_regs_data_and_496_ssc;
  wire act_regs_data_and_497_ssc;
  wire act_regs_data_and_125_ssc;
  reg act_regs_data_1_1_sva_8_31;
  reg [30:0] act_regs_data_1_1_sva_8_30_0;
  wire act_regs_data_and_438_ssc;
  wire act_regs_data_and_439_ssc;
  wire act_regs_data_and_96_ssc;
  reg act_regs_data_2_14_sva_8_31;
  reg [30:0] act_regs_data_2_14_sva_8_30_0;
  wire act_regs_data_and_498_ssc;
  wire act_regs_data_and_499_ssc;
  wire act_regs_data_and_126_ssc;
  reg act_regs_data_1_0_sva_8_31;
  reg [30:0] act_regs_data_1_0_sva_8_30_0;
  wire act_regs_data_and_436_ssc;
  wire act_regs_data_and_437_ssc;
  wire act_regs_data_and_95_ssc;
  reg act_regs_data_2_15_sva_8_31;
  reg [30:0] act_regs_data_2_15_sva_8_30_0;
  wire act_regs_data_and_434_ssc;
  wire act_regs_data_and_435_ssc;
  wire act_regs_data_and_94_ssc;
  reg act_regs_data_3_0_sva_8_31;
  reg [30:0] act_regs_data_3_0_sva_8_30_0;
  wire or_848_ssc;
  reg act_regs_data_3_1_sva_8_31;
  reg [30:0] act_regs_data_3_1_sva_8_30_0;
  wire or_847_ssc;
  reg act_regs_data_3_2_sva_8_31;
  reg [30:0] act_regs_data_3_2_sva_8_30_0;
  wire or_846_ssc;
  reg act_regs_data_3_3_sva_8_31;
  reg [30:0] act_regs_data_3_3_sva_8_30_0;
  wire or_845_ssc;
  reg act_regs_data_3_4_sva_8_31;
  reg [30:0] act_regs_data_3_4_sva_8_30_0;
  wire or_844_ssc;
  reg act_regs_data_3_5_sva_8_31;
  reg [30:0] act_regs_data_3_5_sva_8_30_0;
  wire act_regs_data_and_500_ssc;
  wire act_regs_data_and_501_ssc;
  wire act_regs_data_and_127_ssc;
  reg act_regs_data_0_9_sva_8_31;
  reg [30:0] act_regs_data_0_9_sva_8_30_0;
  wire or_843_ssc;
  reg act_regs_data_3_6_sva_8_31;
  reg [30:0] act_regs_data_3_6_sva_8_30_0;
  wire or_842_ssc;
  reg act_regs_data_3_7_sva_8_31;
  reg [30:0] act_regs_data_3_7_sva_8_30_0;
  wire or_841_ssc;
  reg act_regs_data_3_8_sva_8_31;
  reg [30:0] act_regs_data_3_8_sva_8_30_0;
  wire or_840_ssc;
  reg act_regs_data_3_9_sva_8_31;
  reg [30:0] act_regs_data_3_9_sva_8_30_0;
  wire or_839_ssc;
  reg act_regs_data_3_10_sva_8_31;
  reg [30:0] act_regs_data_3_10_sva_8_30_0;
  wire or_838_ssc;
  reg act_regs_data_3_11_sva_8_31;
  reg [30:0] act_regs_data_3_11_sva_8_30_0;
  wire or_837_ssc;
  reg act_regs_data_3_12_sva_8_31;
  reg [30:0] act_regs_data_3_12_sva_8_30_0;
  wire or_836_ssc;
  reg act_regs_data_3_13_sva_8_31;
  reg [30:0] act_regs_data_3_13_sva_8_30_0;
  wire or_833_ssc;
  reg act_regs_data_3_14_sva_8_31;
  reg [30:0] act_regs_data_3_14_sva_8_30_0;
  wire or_832_ssc;
  reg act_regs_data_3_15_sva_8_31;
  reg [30:0] act_regs_data_3_15_sva_8_30_0;
  wire nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31;
  wire [30:0] nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
  wire nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31;
  wire [30:0] nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
  wire act_regs_data_and_299_cse;
  wire act_regs_data_and_300_cse;
  wire act_regs_data_and_301_cse;
  wire act_regs_data_and_302_cse;
  wire act_regs_data_and_303_cse;
  wire act_regs_data_and_304_cse;
  wire act_regs_data_and_305_cse;
  wire act_regs_data_and_523_cse;
  wire act_regs_data_and_524_cse;
  wire act_regs_data_and_525_cse;
  wire act_regs_data_and_526_cse;
  wire act_regs_data_and_527_cse;
  wire act_regs_data_and_528_cse;
  wire act_regs_data_and_529_cse;
  wire act_regs_data_and_635_cse;
  wire act_regs_data_and_636_cse;
  wire act_regs_data_and_637_cse;
  wire act_regs_data_and_638_cse;
  wire act_regs_data_and_639_cse;
  wire act_regs_data_and_640_cse;
  wire act_regs_data_and_641_cse;
  wire act_regs_data_and_747_cse;
  wire act_regs_data_and_748_cse;
  wire act_regs_data_and_749_cse;
  wire act_regs_data_and_750_cse;
  wire act_regs_data_and_751_cse;
  wire act_regs_data_and_752_cse;
  wire act_regs_data_and_753_cse;
  wire or_tmp_421;
  wire nand_tmp_13;
  wire or_tmp_446;
  wire or_tmp_517;
  wire or_tmp_518;
  wire or_tmp_547;
  wire nand_tmp_45;
  wire or_tmp_654;
  wire or_tmp_726;
  wire or_tmp_755;
  wire and_1211_cse;
  wire mux_330_cse;
  wire and_1451_cse;
  wire mux_336_cse;
  wire mux_329_cse;
  wire or_1077_cse;
  wire and_1108_cse;
  wire nand_297_cse;
  wire or_1097_cse;
  wire and_1485_cse;
  wire and_1488_cse;
  wire nor_734_cse;
  wire or_1033_cse;
  wire or_1071_cse;
  wire or_1488_cse;
  wire mux_328_cse;
  wire mux_337_cse;
  wire mux_342_cse;
  wire mux_344_cse;
  wire and_1249_cse;
  wire mux_350_cse;
  wire mux_355_cse;
  wire nor_736_cse;
  wire mux_411_cse;
  wire nor_744_cse;
  wire mux_467_cse;
  wire nor_752_cse;
  wire mux_523_cse;
  wire nor_760_cse;
  wire nand_298_cse;
  wire nand_338_cse;
  wire nand_378_cse;
  wire nand_418_cse;
  wire or_dcpl_652;
  wire and_dcpl_1229;
  wire or_dcpl_655;
  wire and_1876_cse;
  reg reg_act_regs_data_3_15_3_enexo;
  reg reg_act_regs_data_2_2_3_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo;
  reg reg_is_start_enexo;
  reg reg_act_regs_data_3_15_sva_dfm_2_1_enexo;
  reg reg_act_regs_data_2_15_3_enexo;
  reg reg_act_regs_data_3_14_3_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_1;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_1;
  reg reg_is_start_enexo_1;
  reg reg_act_regs_data_3_14_sva_dfm_2_1_enexo;
  reg reg_act_regs_data_2_14_3_enexo;
  reg reg_act_regs_data_3_13_3_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_2;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_2;
  reg reg_is_start_enexo_2;
  reg reg_act_regs_data_3_13_sva_dfm_2_1_enexo;
  reg reg_act_regs_data_3_12_3_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_3;
  reg reg_act_regs_data_2_13_3_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_3;
  reg reg_is_start_enexo_3;
  reg reg_act_regs_data_3_12_sva_dfm_2_1_enexo;
  reg reg_act_regs_data_3_11_3_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_4;
  reg reg_act_regs_data_2_12_3_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_4;
  reg reg_is_start_enexo_4;
  reg reg_act_regs_data_3_11_sva_dfm_2_1_enexo;
  reg reg_act_regs_data_3_10_3_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_5;
  reg reg_act_regs_data_2_11_3_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_5;
  reg reg_is_start_enexo_5;
  reg reg_act_regs_data_3_10_sva_dfm_2_1_enexo;
  reg reg_act_regs_data_3_0_3_enexo;
  reg reg_act_regs_data_3_9_3_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_6;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_6;
  reg reg_is_start_enexo_6;
  reg reg_act_regs_data_3_9_sva_dfm_2_1_enexo;
  reg reg_act_regs_data_3_8_3_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_7;
  reg reg_act_regs_data_2_9_3_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_7;
  reg reg_is_start_enexo_7;
  reg reg_act_regs_data_3_8_sva_dfm_2_1_enexo;
  reg reg_act_regs_data_3_7_3_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_8;
  reg reg_act_regs_data_2_8_3_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_8;
  reg reg_is_start_enexo_8;
  reg reg_act_regs_data_3_7_sva_dfm_2_1_enexo;
  reg reg_act_regs_data_3_6_3_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_9;
  reg reg_act_regs_data_2_7_3_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_9;
  reg reg_is_start_enexo_9;
  reg reg_act_regs_data_3_6_sva_dfm_2_1_enexo;
  reg reg_act_regs_data_3_5_3_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_10;
  reg reg_act_regs_data_2_6_3_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_10;
  reg reg_is_start_enexo_10;
  reg reg_act_regs_data_3_5_sva_dfm_2_1_enexo;
  reg reg_act_regs_data_3_4_3_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_11;
  reg reg_act_regs_data_2_5_3_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_11;
  reg reg_is_start_enexo_11;
  reg reg_act_regs_data_3_4_sva_dfm_2_1_enexo;
  reg reg_act_regs_data_3_3_3_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_12;
  reg reg_act_regs_data_2_4_3_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_12;
  reg reg_is_start_enexo_12;
  reg reg_act_regs_data_3_3_sva_dfm_2_1_enexo;
  reg reg_act_regs_data_3_2_3_enexo;
  reg reg_act_regs_data_2_3_3_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_13;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_13;
  reg reg_is_start_enexo_13;
  reg reg_act_regs_data_3_2_sva_dfm_2_1_enexo;
  reg reg_act_regs_data_3_1_3_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_14;
  reg reg_act_regs_data_2_10_3_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_14;
  reg reg_is_start_enexo_14;
  reg reg_act_regs_data_3_1_sva_dfm_2_1_enexo;
  reg reg_act_regs_data_3_0_3_enexo_1;
  reg reg_act_regs_data_2_1_3_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_15;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_15;
  reg reg_is_start_enexo_15;
  reg reg_act_regs_data_3_0_sva_dfm_2_1_enexo;
  reg reg_act_regs_data_2_15_3_enexo_1;
  reg reg_w_load_lpi_1_dfm_1_enexo_16;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_16;
  reg reg_act_regs_data_1_2_3_enexo;
  reg reg_is_start_enexo_16;
  reg reg_act_regs_data_2_15_sva_dfm_2_1_enexo;
  reg reg_act_regs_data_2_14_3_enexo_1;
  reg reg_act_regs_data_1_15_3_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_17;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_17;
  reg reg_is_start_enexo_17;
  reg reg_act_regs_data_2_14_sva_dfm_2_1_enexo;
  reg reg_act_regs_data_1_14_3_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_18;
  reg reg_act_regs_data_2_13_3_enexo_1;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_18;
  reg reg_is_start_enexo_18;
  reg reg_act_regs_data_2_13_sva_dfm_2_1_enexo;
  reg reg_act_regs_data_1_13_3_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_19;
  reg reg_act_regs_data_2_12_3_enexo_1;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_19;
  reg reg_is_start_enexo_19;
  reg reg_act_regs_data_2_12_sva_dfm_2_1_enexo;
  reg reg_act_regs_data_1_12_3_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_20;
  reg reg_act_regs_data_2_11_3_enexo_1;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_20;
  reg reg_is_start_enexo_20;
  reg reg_act_regs_data_2_11_sva_dfm_2_1_enexo;
  reg reg_act_regs_data_1_11_3_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_21;
  reg reg_act_regs_data_2_10_3_enexo_1;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_21;
  reg reg_is_start_enexo_21;
  reg reg_act_regs_data_2_10_sva_dfm_2_1_enexo;
  reg reg_act_regs_data_2_0_3_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_22;
  reg reg_act_regs_data_2_9_3_enexo_1;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_22;
  reg reg_is_start_enexo_22;
  reg reg_act_regs_data_2_9_sva_dfm_2_1_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_23;
  reg reg_act_regs_data_2_8_3_enexo_1;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_23;
  reg reg_act_regs_data_1_9_3_enexo;
  reg reg_is_start_enexo_23;
  reg reg_act_regs_data_2_8_sva_dfm_2_1_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_24;
  reg reg_act_regs_data_2_7_3_enexo_1;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_24;
  reg reg_act_regs_data_1_8_3_enexo;
  reg reg_is_start_enexo_24;
  reg reg_act_regs_data_2_7_sva_dfm_2_1_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_25;
  reg reg_act_regs_data_2_6_3_enexo_1;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_25;
  reg reg_act_regs_data_1_7_3_enexo;
  reg reg_is_start_enexo_25;
  reg reg_act_regs_data_2_6_sva_dfm_2_1_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_26;
  reg reg_act_regs_data_2_5_3_enexo_1;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_26;
  reg reg_act_regs_data_1_6_3_enexo;
  reg reg_is_start_enexo_26;
  reg reg_act_regs_data_2_5_sva_dfm_2_1_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_27;
  reg reg_act_regs_data_2_4_3_enexo_1;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_27;
  reg reg_act_regs_data_1_5_3_enexo;
  reg reg_is_start_enexo_27;
  reg reg_act_regs_data_2_4_sva_dfm_2_1_enexo;
  reg reg_act_regs_data_2_3_3_enexo_1;
  reg reg_w_load_lpi_1_dfm_1_enexo_28;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_28;
  reg reg_act_regs_data_1_4_3_enexo;
  reg reg_is_start_enexo_28;
  reg reg_act_regs_data_2_3_sva_dfm_2_1_enexo;
  reg reg_act_regs_data_2_2_3_enexo_1;
  reg reg_w_load_lpi_1_dfm_1_enexo_29;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_29;
  reg reg_act_regs_data_1_3_3_enexo;
  reg reg_is_start_enexo_29;
  reg reg_act_regs_data_2_2_sva_dfm_2_1_enexo;
  reg reg_act_regs_data_2_1_3_enexo_1;
  reg reg_act_regs_data_1_10_3_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_30;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_30;
  reg reg_is_start_enexo_30;
  reg reg_act_regs_data_2_1_sva_dfm_2_1_enexo;
  reg reg_act_regs_data_2_0_3_enexo_1;
  reg reg_w_load_lpi_1_dfm_1_enexo_31;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_31;
  reg reg_act_regs_data_1_1_3_enexo;
  reg reg_is_start_enexo_31;
  reg reg_act_regs_data_2_0_sva_dfm_2_1_enexo;
  reg reg_act_regs_data_1_15_3_enexo_1;
  reg reg_w_load_lpi_1_dfm_1_enexo_32;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_32;
  reg reg_act_regs_data_0_2_3_enexo;
  reg reg_is_start_enexo_32;
  reg reg_act_regs_data_1_15_sva_dfm_2_1_enexo;
  reg reg_act_regs_data_1_14_3_enexo_1;
  reg reg_w_load_lpi_1_dfm_1_enexo_33;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_33;
  reg reg_is_start_enexo_33;
  reg reg_act_regs_data_1_14_sva_dfm_2_1_enexo;
  reg reg_act_regs_data_0_15_3_enexo;
  reg reg_act_regs_data_1_13_3_enexo_1;
  reg reg_w_load_lpi_1_dfm_1_enexo_34;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_34;
  reg reg_is_start_enexo_34;
  reg reg_act_regs_data_1_13_sva_dfm_2_1_enexo;
  reg reg_act_regs_data_0_14_3_enexo;
  reg reg_act_regs_data_1_12_3_enexo_1;
  reg reg_w_load_lpi_1_dfm_1_enexo_35;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_35;
  reg reg_is_start_enexo_35;
  reg reg_act_regs_data_0_13_3_enexo;
  reg reg_act_regs_data_1_12_sva_dfm_2_1_enexo;
  reg reg_act_regs_data_1_11_3_enexo_1;
  reg reg_w_load_lpi_1_dfm_1_enexo_36;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_36;
  reg reg_is_start_enexo_36;
  reg reg_act_regs_data_0_12_3_enexo;
  reg reg_act_regs_data_1_11_sva_dfm_2_1_enexo;
  reg reg_act_regs_data_1_10_3_enexo_1;
  reg reg_w_load_lpi_1_dfm_1_enexo_37;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_37;
  reg reg_is_start_enexo_37;
  reg reg_act_regs_data_0_11_3_enexo;
  reg reg_act_regs_data_1_10_sva_dfm_2_1_enexo;
  reg reg_act_regs_data_1_0_3_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_38;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_38;
  reg reg_act_regs_data_1_9_3_enexo_1;
  reg reg_is_start_enexo_38;
  reg reg_act_regs_data_1_9_sva_dfm_2_1_enexo;
  reg reg_act_regs_data_0_9_3_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_39;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_39;
  reg reg_act_regs_data_1_8_3_enexo_1;
  reg reg_is_start_enexo_39;
  reg reg_act_regs_data_1_8_sva_dfm_2_1_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_40;
  reg reg_act_regs_data_0_8_3_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_40;
  reg reg_act_regs_data_1_7_3_enexo_1;
  reg reg_is_start_enexo_40;
  reg reg_act_regs_data_1_7_sva_dfm_2_1_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_41;
  reg reg_act_regs_data_0_7_3_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_41;
  reg reg_act_regs_data_1_6_3_enexo_1;
  reg reg_is_start_enexo_41;
  reg reg_act_regs_data_1_6_sva_dfm_2_1_enexo;
  reg reg_act_regs_data_0_6_3_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_42;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_42;
  reg reg_act_regs_data_1_5_3_enexo_1;
  reg reg_is_start_enexo_42;
  reg reg_act_regs_data_1_5_sva_dfm_2_1_enexo;
  reg reg_act_regs_data_0_5_3_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_43;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_43;
  reg reg_act_regs_data_1_4_3_enexo_1;
  reg reg_is_start_enexo_43;
  reg reg_act_regs_data_1_4_sva_dfm_2_1_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_44;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_44;
  reg reg_act_regs_data_0_4_3_enexo;
  reg reg_act_regs_data_1_3_3_enexo_1;
  reg reg_is_start_enexo_44;
  reg reg_act_regs_data_1_3_sva_dfm_2_1_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_45;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_45;
  reg reg_act_regs_data_0_3_3_enexo;
  reg reg_act_regs_data_1_2_3_enexo_1;
  reg reg_is_start_enexo_45;
  reg reg_act_regs_data_1_2_sva_dfm_2_1_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_46;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_46;
  reg reg_act_regs_data_1_1_3_enexo_1;
  reg reg_is_start_enexo_46;
  reg reg_act_regs_data_0_10_3_enexo;
  reg reg_act_regs_data_1_1_sva_dfm_2_1_enexo;
  reg reg_act_regs_data_1_0_3_enexo_1;
  reg reg_w_load_lpi_1_dfm_1_enexo_47;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_47;
  reg reg_act_regs_data_0_1_3_enexo;
  reg reg_is_start_enexo_47;
  reg reg_act_regs_data_1_0_sva_dfm_2_1_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_48;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_48;
  reg reg_ActUnit_PushOutput_if_output_port_reg_data_data_2_1_enexo;
  reg reg_is_start_enexo_48;
  reg reg_act_regs_data_0_15_sva_dfm_2_1_enexo;
  reg reg_act_regs_data_0_15_3_enexo_1;
  reg reg_w_load_lpi_1_dfm_1_enexo_49;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_49;
  reg reg_ActUnit_PushOutput_if_output_port_reg_data_data_14_1_enexo;
  reg reg_is_start_enexo_49;
  reg reg_act_regs_data_0_14_sva_dfm_2_1_enexo;
  reg reg_act_regs_data_0_14_3_enexo_1;
  reg reg_w_load_lpi_1_dfm_1_enexo_50;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_50;
  reg reg_is_start_enexo_50;
  reg reg_ActUnit_PushOutput_if_output_port_reg_data_data_13_1_enexo;
  reg reg_act_regs_data_0_13_3_enexo_1;
  reg reg_act_regs_data_0_13_sva_dfm_2_1_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_51;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_51;
  reg reg_ActUnit_PushOutput_if_output_port_reg_data_data_12_1_enexo;
  reg reg_is_start_enexo_51;
  reg reg_act_regs_data_0_12_3_enexo_1;
  reg reg_act_regs_data_0_12_sva_dfm_2_1_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_52;
  reg reg_ActUnit_PushOutput_if_output_port_reg_data_data_11_1_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_52;
  reg reg_is_start_enexo_52;
  reg reg_act_regs_data_0_11_3_enexo_1;
  reg reg_act_regs_data_0_11_sva_dfm_2_1_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_53;
  reg reg_ActUnit_PushOutput_if_output_port_reg_data_data_10_1_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_53;
  reg reg_is_start_enexo_53;
  reg reg_act_regs_data_0_10_3_enexo_1;
  reg reg_act_regs_data_0_10_sva_dfm_2_1_enexo;
  reg reg_act_regs_data_0_9_3_enexo_1;
  reg reg_w_load_lpi_1_dfm_1_enexo_54;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_54;
  reg reg_act_regs_data_0_0_3_enexo;
  reg reg_is_start_enexo_54;
  reg reg_act_regs_data_0_9_sva_dfm_2_1_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_55;
  reg reg_act_regs_data_0_8_3_enexo_1;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_55;
  reg reg_is_start_enexo_55;
  reg reg_ActUnit_PushOutput_if_output_port_reg_data_data_9_1_enexo;
  reg reg_act_regs_data_0_8_sva_dfm_2_1_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_56;
  reg reg_act_regs_data_0_7_3_enexo_1;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_56;
  reg reg_ActUnit_PushOutput_if_output_port_reg_data_data_8_1_enexo;
  reg reg_is_start_enexo_56;
  reg reg_act_regs_data_0_7_sva_dfm_2_1_enexo;
  reg reg_ActUnit_PushOutput_if_output_port_reg_data_data_7_1_enexo;
  reg reg_act_regs_data_0_6_3_enexo_1;
  reg reg_w_load_lpi_1_dfm_1_enexo_57;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_57;
  reg reg_is_start_enexo_57;
  reg reg_act_regs_data_0_6_sva_dfm_2_1_enexo;
  reg reg_act_regs_data_0_5_3_enexo_1;
  reg reg_w_load_lpi_1_dfm_1_enexo_58;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_58;
  reg reg_is_start_enexo_58;
  reg reg_ActUnit_PushOutput_if_output_port_reg_data_data_6_1_enexo;
  reg reg_act_regs_data_0_5_sva_dfm_2_1_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_59;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_59;
  reg reg_act_regs_data_0_4_3_enexo_1;
  reg reg_is_start_enexo_59;
  reg reg_ActUnit_PushOutput_if_output_port_reg_data_data_5_1_enexo;
  reg reg_act_regs_data_0_4_sva_dfm_2_1_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_60;
  reg reg_ActUnit_PushOutput_if_output_port_reg_data_data_4_1_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_60;
  reg reg_act_regs_data_0_3_3_enexo_1;
  reg reg_is_start_enexo_60;
  reg reg_act_regs_data_0_3_sva_dfm_2_1_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_61;
  reg reg_ActUnit_PushOutput_if_output_port_reg_data_data_3_1_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_61;
  reg reg_act_regs_data_0_2_3_enexo_1;
  reg reg_is_start_enexo_61;
  reg reg_act_regs_data_0_2_sva_dfm_2_1_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_62;
  reg reg_ActUnit_PushOutput_if_output_port_reg_data_data_1_1_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_62;
  reg reg_act_regs_data_0_1_3_enexo_1;
  reg reg_is_start_enexo_62;
  reg reg_act_regs_data_0_1_sva_dfm_2_1_enexo;
  reg reg_ActUnit_PushOutput_if_output_port_reg_data_data_0_1_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_63;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_63;
  reg reg_act_regs_data_0_0_3_enexo_1;
  reg reg_is_start_enexo_63;
  reg reg_act_regs_data_0_0_sva_dfm_2_1_enexo;
  reg reg_act_mem_banks_read_for_mux_15_enexo;
  reg reg_act_mem_banks_read_for_mux_14_enexo;
  reg reg_act_mem_banks_read_for_mux_13_enexo;
  reg reg_act_mem_banks_read_for_mux_12_enexo;
  reg reg_act_mem_banks_read_for_mux_11_enexo;
  reg reg_act_mem_banks_read_for_mux_10_enexo;
  reg reg_act_mem_banks_read_for_mux_9_enexo;
  reg reg_act_mem_banks_read_for_mux_8_enexo;
  reg reg_act_mem_banks_read_for_mux_7_enexo;
  reg reg_act_mem_banks_read_for_mux_6_enexo;
  reg reg_act_mem_banks_read_for_mux_5_enexo;
  reg reg_act_mem_banks_read_for_mux_4_enexo;
  reg reg_act_mem_banks_read_for_mux_3_enexo;
  reg reg_act_mem_banks_read_for_mux_2_enexo;
  reg reg_act_mem_banks_read_for_mux_1_enexo;
  reg reg_act_mem_banks_read_for_mux_enexo;
  reg reg_act_mem_banks_read_for_mux_15_enexo_1;
  reg reg_act_mem_banks_read_read_data_lpi_1_dfm_1_31_0_enexo;
  reg reg_ActUnit_CheckStart_start_reg_enexo;
  reg reg_act_mem_banks_read_read_data_lpi_1_dfm_1_63_32_enexo;
  reg reg_ActUnit_CheckStart_start_reg_enexo_1;
  reg reg_act_mem_banks_read_for_mux_14_enexo_1;
  reg reg_act_mem_banks_read_read_data_lpi_1_dfm_1_95_64_enexo;
  reg reg_ActUnit_CheckStart_start_reg_enexo_2;
  reg reg_act_mem_banks_read_for_mux_13_enexo_1;
  reg reg_ActUnit_CheckStart_start_reg_enexo_3;
  reg reg_act_mem_banks_read_for_mux_12_enexo_1;
  reg reg_act_mem_banks_read_read_data_lpi_1_dfm_1_127_96_enexo;
  reg reg_act_mem_banks_read_for_mux_11_enexo_1;
  reg reg_ActUnit_CheckStart_start_reg_enexo_4;
  reg reg_act_mem_banks_read_read_data_lpi_1_dfm_1_159_128_enexo;
  reg reg_act_mem_banks_read_for_mux_10_enexo_1;
  reg reg_act_mem_banks_read_read_data_lpi_1_dfm_1_191_160_enexo;
  reg reg_ActUnit_CheckStart_start_reg_enexo_5;
  reg reg_act_mem_banks_read_for_mux_9_enexo_1;
  reg reg_act_mem_banks_read_read_data_lpi_1_dfm_1_223_192_enexo;
  reg reg_ActUnit_CheckStart_start_reg_enexo_6;
  reg reg_act_mem_banks_read_for_mux_8_enexo_1;
  reg reg_ActUnit_CheckStart_start_reg_enexo_7;
  reg reg_act_mem_banks_read_read_data_lpi_1_dfm_1_255_224_enexo;
  reg reg_act_mem_banks_read_read_data_lpi_1_dfm_1_287_256_enexo;
  reg reg_act_mem_banks_read_for_mux_7_enexo_1;
  reg reg_ActUnit_CheckStart_start_reg_enexo_8;
  reg reg_act_mem_banks_read_for_mux_6_enexo_1;
  reg reg_act_mem_banks_read_read_data_lpi_1_dfm_1_319_288_enexo;
  reg reg_ActUnit_CheckStart_start_reg_enexo_9;
  reg reg_act_mem_banks_read_for_mux_5_enexo_1;
  reg reg_ActUnit_CheckStart_start_reg_enexo_10;
  reg reg_act_mem_banks_read_read_data_lpi_1_dfm_1_351_320_enexo;
  reg reg_act_mem_banks_read_for_mux_4_enexo_1;
  reg reg_act_mem_banks_read_read_data_lpi_1_dfm_1_383_352_enexo;
  reg reg_ActUnit_CheckStart_start_reg_enexo_11;
  reg reg_act_mem_banks_read_read_data_lpi_1_dfm_1_415_384_enexo;
  reg reg_act_mem_banks_read_for_mux_3_enexo_1;
  reg reg_ActUnit_CheckStart_start_reg_enexo_12;
  reg reg_act_mem_banks_read_read_data_lpi_1_dfm_1_447_416_enexo;
  reg reg_act_mem_banks_read_for_mux_2_enexo_1;
  reg reg_ActUnit_CheckStart_start_reg_enexo_13;
  reg reg_act_mem_banks_read_read_data_lpi_1_dfm_1_479_448_enexo;
  reg reg_act_mem_banks_read_for_mux_1_enexo_1;
  reg reg_ActUnit_CheckStart_start_reg_enexo_14;
  reg reg_act_mem_banks_read_for_mux_enexo_1;
  reg reg_ActUnit_CheckStart_start_reg_enexo_15;
  reg reg_act_mem_banks_read_read_data_lpi_1_dfm_1_511_480_enexo;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo;
  reg reg_act_regs_data_1_15_2_enexo;
  reg reg_act_regs_data_2_15_2_enexo;
  reg reg_act_regs_data_0_15_2_enexo;
  reg reg_act_config_inst_counter_enexo;
  reg reg_act_regs_data_3_15_2_enexo;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_1;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_1;
  reg reg_act_regs_data_3_14_2_enexo;
  reg reg_act_regs_data_0_14_2_enexo;
  reg reg_act_regs_data_1_14_2_enexo;
  reg reg_act_regs_data_2_14_2_enexo;
  reg reg_act_config_inst_counter_enexo_1;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_2;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_2;
  reg reg_act_regs_data_1_13_2_enexo;
  reg reg_act_regs_data_0_13_2_enexo;
  reg reg_act_regs_data_3_13_2_enexo;
  reg reg_act_regs_data_2_13_2_enexo;
  reg reg_act_config_inst_counter_enexo_2;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_3;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_3;
  reg reg_act_regs_data_1_12_2_enexo;
  reg reg_act_regs_data_2_12_2_enexo;
  reg reg_act_regs_data_0_12_2_enexo;
  reg reg_act_regs_data_3_12_2_enexo;
  reg reg_act_config_inst_counter_enexo_3;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_4;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_4;
  reg reg_act_regs_data_2_11_2_enexo;
  reg reg_act_regs_data_3_11_2_enexo;
  reg reg_act_regs_data_1_11_2_enexo;
  reg reg_act_regs_data_0_11_2_enexo;
  reg reg_act_config_inst_counter_enexo_4;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_5;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_5;
  reg reg_act_regs_data_0_10_2_enexo;
  reg reg_act_regs_data_1_10_2_enexo;
  reg reg_act_regs_data_2_10_2_enexo;
  reg reg_act_regs_data_3_10_2_enexo;
  reg reg_act_config_inst_counter_enexo_5;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_6;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_6;
  reg reg_act_regs_data_1_9_2_enexo;
  reg reg_act_regs_data_0_9_2_enexo;
  reg reg_act_regs_data_2_9_2_enexo;
  reg reg_act_regs_data_3_9_2_enexo;
  reg reg_act_config_inst_counter_enexo_6;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_7;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_7;
  reg reg_act_regs_data_3_8_2_enexo;
  reg reg_act_regs_data_1_8_2_enexo;
  reg reg_act_regs_data_0_8_2_enexo;
  reg reg_act_regs_data_2_8_2_enexo;
  reg reg_act_config_inst_counter_enexo_7;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_8;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_8;
  reg reg_act_regs_data_2_7_2_enexo;
  reg reg_act_regs_data_1_7_2_enexo;
  reg reg_act_regs_data_0_7_2_enexo;
  reg reg_act_regs_data_3_7_2_enexo;
  reg reg_act_config_inst_counter_enexo_8;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_9;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_9;
  reg reg_act_regs_data_3_6_2_enexo;
  reg reg_act_regs_data_1_6_2_enexo;
  reg reg_act_regs_data_0_6_2_enexo;
  reg reg_act_regs_data_2_6_2_enexo;
  reg reg_act_config_inst_counter_enexo_9;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_10;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_10;
  reg reg_act_regs_data_0_5_2_enexo;
  reg reg_act_regs_data_2_5_2_enexo;
  reg reg_act_regs_data_3_5_2_enexo;
  reg reg_act_regs_data_1_5_2_enexo;
  reg reg_act_config_inst_counter_enexo_10;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_11;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_11;
  reg reg_act_regs_data_2_4_2_enexo;
  reg reg_act_regs_data_3_4_2_enexo;
  reg reg_act_regs_data_1_4_2_enexo;
  reg reg_act_regs_data_0_4_2_enexo;
  reg reg_act_config_inst_counter_enexo_11;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_12;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_12;
  reg reg_act_regs_data_2_3_2_enexo;
  reg reg_act_regs_data_3_3_2_enexo;
  reg reg_act_regs_data_1_3_2_enexo;
  reg reg_act_regs_data_0_3_2_enexo;
  reg reg_act_config_inst_counter_enexo_12;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_13;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_13;
  reg reg_act_regs_data_0_2_2_enexo;
  reg reg_act_regs_data_2_2_2_enexo;
  reg reg_act_regs_data_1_2_2_enexo;
  reg reg_act_regs_data_3_2_2_enexo;
  reg reg_act_config_inst_counter_enexo_13;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_14;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_14;
  reg reg_act_regs_data_1_1_2_enexo;
  reg reg_act_regs_data_3_1_2_enexo;
  reg reg_act_regs_data_0_1_2_enexo;
  reg reg_act_regs_data_2_1_2_enexo;
  reg reg_act_config_inst_counter_enexo_14;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_15;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_15;
  reg reg_act_regs_data_2_0_2_enexo;
  reg reg_act_regs_data_3_0_2_enexo;
  reg reg_act_regs_data_1_0_2_enexo;
  reg reg_act_regs_data_0_0_2_enexo;
  reg reg_act_config_inst_counter_enexo_15;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_16;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_16;
  reg reg_act_regs_data_3_15_enexo;
  reg reg_act_regs_data_1_15_2_enexo_1;
  reg reg_act_regs_data_2_15_2_enexo_1;
  reg reg_act_regs_data_0_15_2_enexo_1;
  reg reg_act_config_inst_counter_enexo_16;
  reg reg_act_regs_data_3_15_2_enexo_1;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_17;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_17;
  reg reg_act_regs_data_1_14_enexo;
  reg reg_act_regs_data_3_14_2_enexo_1;
  reg reg_act_regs_data_0_14_2_enexo_1;
  reg reg_act_regs_data_1_14_2_enexo_1;
  reg reg_act_regs_data_2_14_2_enexo_1;
  reg reg_act_config_inst_counter_enexo_17;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_18;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_18;
  reg reg_act_regs_data_1_13_2_enexo_1;
  reg reg_act_regs_data_1_13_enexo;
  reg reg_act_regs_data_0_13_2_enexo_1;
  reg reg_act_regs_data_3_13_2_enexo_1;
  reg reg_act_regs_data_2_13_2_enexo_1;
  reg reg_act_config_inst_counter_enexo_18;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_19;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_19;
  reg reg_act_regs_data_1_12_enexo;
  reg reg_act_regs_data_1_12_2_enexo_1;
  reg reg_act_regs_data_2_12_2_enexo_1;
  reg reg_act_regs_data_0_12_2_enexo_1;
  reg reg_act_regs_data_3_12_2_enexo_1;
  reg reg_act_config_inst_counter_enexo_19;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_20;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_20;
  reg reg_act_regs_data_1_11_enexo;
  reg reg_act_regs_data_2_11_2_enexo_1;
  reg reg_act_regs_data_3_11_2_enexo_1;
  reg reg_act_regs_data_1_11_2_enexo_1;
  reg reg_act_regs_data_0_11_2_enexo_1;
  reg reg_act_config_inst_counter_enexo_20;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_21;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_21;
  reg reg_act_regs_data_0_10_2_enexo_1;
  reg reg_act_regs_data_2_10_enexo;
  reg reg_act_regs_data_1_10_2_enexo_1;
  reg reg_act_regs_data_2_10_2_enexo_1;
  reg reg_act_regs_data_3_10_2_enexo_1;
  reg reg_act_config_inst_counter_enexo_21;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_22;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_22;
  reg reg_act_regs_data_0_9_enexo;
  reg reg_act_regs_data_1_9_2_enexo_1;
  reg reg_act_regs_data_0_9_2_enexo_1;
  reg reg_act_regs_data_2_9_2_enexo_1;
  reg reg_act_regs_data_3_9_2_enexo_1;
  reg reg_act_config_inst_counter_enexo_22;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_23;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_23;
  reg reg_act_regs_data_0_8_enexo;
  reg reg_act_regs_data_3_8_2_enexo_1;
  reg reg_act_regs_data_1_8_2_enexo_1;
  reg reg_act_regs_data_0_8_2_enexo_1;
  reg reg_act_regs_data_2_8_2_enexo_1;
  reg reg_act_config_inst_counter_enexo_23;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_24;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_24;
  reg reg_act_regs_data_2_7_2_enexo_1;
  reg reg_act_regs_data_1_7_enexo;
  reg reg_act_regs_data_1_7_2_enexo_1;
  reg reg_act_regs_data_0_7_2_enexo_1;
  reg reg_act_regs_data_3_7_2_enexo_1;
  reg reg_act_config_inst_counter_enexo_24;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_25;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_25;
  reg reg_act_regs_data_2_6_enexo;
  reg reg_act_regs_data_3_6_2_enexo_1;
  reg reg_act_regs_data_1_6_2_enexo_1;
  reg reg_act_regs_data_0_6_2_enexo_1;
  reg reg_act_regs_data_2_6_2_enexo_1;
  reg reg_act_config_inst_counter_enexo_25;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_26;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_26;
  reg reg_act_regs_data_0_5_2_enexo_1;
  reg reg_act_regs_data_2_5_2_enexo_1;
  reg reg_act_regs_data_3_5_enexo;
  reg reg_act_regs_data_3_5_2_enexo_1;
  reg reg_act_regs_data_1_5_2_enexo_1;
  reg reg_act_config_inst_counter_enexo_26;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_27;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_27;
  reg reg_act_regs_data_1_4_enexo;
  reg reg_act_regs_data_2_4_2_enexo_1;
  reg reg_act_regs_data_3_4_2_enexo_1;
  reg reg_act_regs_data_1_4_2_enexo_1;
  reg reg_act_regs_data_0_4_2_enexo_1;
  reg reg_act_config_inst_counter_enexo_27;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_28;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_28;
  reg reg_act_regs_data_0_3_enexo;
  reg reg_act_regs_data_2_3_2_enexo_1;
  reg reg_act_regs_data_3_3_2_enexo_1;
  reg reg_act_regs_data_1_3_2_enexo_1;
  reg reg_act_regs_data_0_3_2_enexo_1;
  reg reg_act_config_inst_counter_enexo_28;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_29;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_29;
  reg reg_act_regs_data_1_2_enexo;
  reg reg_act_regs_data_0_2_2_enexo_1;
  reg reg_act_regs_data_2_2_2_enexo_1;
  reg reg_act_regs_data_1_2_2_enexo_1;
  reg reg_act_regs_data_3_2_2_enexo_1;
  reg reg_act_config_inst_counter_enexo_29;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_30;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_30;
  reg reg_act_regs_data_0_1_enexo;
  reg reg_act_regs_data_1_1_2_enexo_1;
  reg reg_act_regs_data_3_1_2_enexo_1;
  reg reg_act_regs_data_0_1_2_enexo_1;
  reg reg_act_regs_data_2_1_2_enexo_1;
  reg reg_act_config_inst_counter_enexo_30;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_31;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_31;
  reg reg_act_regs_data_2_0_enexo;
  reg reg_act_regs_data_2_0_2_enexo_1;
  reg reg_act_regs_data_3_0_2_enexo_1;
  reg reg_act_regs_data_1_0_2_enexo_1;
  reg reg_act_regs_data_0_0_2_enexo_1;
  reg reg_act_config_inst_counter_enexo_31;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_32;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_32;
  reg reg_act_regs_data_0_2_2_enexo_2;
  reg reg_act_regs_data_2_2_2_enexo_2;
  reg reg_act_regs_data_1_2_2_enexo_2;
  reg reg_act_regs_data_3_2_2_enexo_2;
  reg reg_act_config_inst_counter_enexo_32;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_33;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_33;
  reg reg_act_regs_data_2_3_2_enexo_2;
  reg reg_act_regs_data_3_3_2_enexo_2;
  reg reg_act_regs_data_1_3_2_enexo_2;
  reg reg_act_regs_data_0_3_2_enexo_2;
  reg reg_act_config_inst_counter_enexo_33;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_34;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_34;
  reg reg_act_regs_data_2_0_2_enexo_2;
  reg reg_act_regs_data_3_0_2_enexo_2;
  reg reg_act_regs_data_1_0_2_enexo_2;
  reg reg_act_regs_data_0_0_2_enexo_2;
  reg reg_act_config_inst_counter_enexo_34;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_35;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_35;
  reg reg_act_regs_data_1_1_2_enexo_2;
  reg reg_act_regs_data_3_1_2_enexo_2;
  reg reg_act_regs_data_0_1_2_enexo_2;
  reg reg_act_regs_data_2_1_2_enexo_2;
  reg reg_act_config_inst_counter_enexo_35;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_36;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_36;
  reg reg_act_regs_data_2_4_2_enexo_2;
  reg reg_act_regs_data_3_4_2_enexo_2;
  reg reg_act_regs_data_1_4_2_enexo_2;
  reg reg_act_regs_data_0_4_2_enexo_2;
  reg reg_act_config_inst_counter_enexo_36;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_37;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_37;
  reg reg_act_regs_data_0_5_2_enexo_2;
  reg reg_act_regs_data_2_5_2_enexo_2;
  reg reg_act_regs_data_3_5_2_enexo_2;
  reg reg_act_regs_data_1_5_2_enexo_2;
  reg reg_act_config_inst_counter_enexo_37;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_38;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_38;
  reg reg_act_regs_data_3_6_2_enexo_2;
  reg reg_act_regs_data_1_6_2_enexo_2;
  reg reg_act_regs_data_0_6_2_enexo_2;
  reg reg_act_regs_data_2_6_2_enexo_2;
  reg reg_act_config_inst_counter_enexo_38;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_39;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_39;
  reg reg_act_regs_data_2_7_2_enexo_2;
  reg reg_act_regs_data_1_7_2_enexo_2;
  reg reg_act_regs_data_0_7_2_enexo_2;
  reg reg_act_regs_data_3_7_2_enexo_2;
  reg reg_act_config_inst_counter_enexo_39;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_40;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_40;
  reg reg_act_regs_data_3_8_2_enexo_2;
  reg reg_act_regs_data_1_8_2_enexo_2;
  reg reg_act_regs_data_0_8_2_enexo_2;
  reg reg_act_regs_data_2_8_2_enexo_2;
  reg reg_act_config_inst_counter_enexo_40;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_41;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_41;
  reg reg_act_regs_data_1_9_2_enexo_2;
  reg reg_act_regs_data_0_9_2_enexo_2;
  reg reg_act_regs_data_2_9_2_enexo_2;
  reg reg_act_regs_data_3_9_2_enexo_2;
  reg reg_act_config_inst_counter_enexo_41;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_42;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_42;
  reg reg_act_regs_data_0_10_2_enexo_2;
  reg reg_act_regs_data_1_10_2_enexo_2;
  reg reg_act_regs_data_2_10_2_enexo_2;
  reg reg_act_regs_data_3_10_2_enexo_2;
  reg reg_act_config_inst_counter_enexo_42;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_43;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_43;
  reg reg_act_regs_data_2_11_2_enexo_2;
  reg reg_act_regs_data_3_11_2_enexo_2;
  reg reg_act_regs_data_1_11_2_enexo_2;
  reg reg_act_regs_data_0_11_2_enexo_2;
  reg reg_act_config_inst_counter_enexo_43;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_44;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_44;
  reg reg_act_regs_data_1_12_2_enexo_2;
  reg reg_act_regs_data_2_12_2_enexo_2;
  reg reg_act_regs_data_0_12_2_enexo_2;
  reg reg_act_regs_data_3_12_2_enexo_2;
  reg reg_act_config_inst_counter_enexo_44;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_45;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_45;
  reg reg_act_regs_data_1_13_2_enexo_2;
  reg reg_act_regs_data_0_13_2_enexo_2;
  reg reg_act_regs_data_3_13_2_enexo_2;
  reg reg_act_regs_data_2_13_2_enexo_2;
  reg reg_act_config_inst_counter_enexo_45;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_46;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_46;
  reg reg_act_regs_data_3_14_2_enexo_2;
  reg reg_act_regs_data_0_14_2_enexo_2;
  reg reg_act_regs_data_1_14_2_enexo_2;
  reg reg_act_regs_data_2_14_2_enexo_2;
  reg reg_act_config_inst_counter_enexo_46;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_47;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_47;
  reg reg_act_regs_data_1_15_2_enexo_2;
  reg reg_act_regs_data_2_15_2_enexo_2;
  reg reg_act_regs_data_0_15_2_enexo_2;
  reg reg_act_config_inst_counter_enexo_47;
  reg reg_act_regs_data_3_15_2_enexo_2;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_48;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_48;
  reg reg_act_regs_data_0_2_2_enexo_3;
  reg reg_act_regs_data_2_2_2_enexo_3;
  reg reg_act_regs_data_1_2_2_enexo_3;
  reg reg_act_regs_data_3_2_2_enexo_3;
  reg reg_act_config_inst_counter_enexo_48;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_49;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_49;
  reg reg_act_regs_data_2_11_2_enexo_3;
  reg reg_act_regs_data_3_11_2_enexo_3;
  reg reg_act_regs_data_1_11_2_enexo_3;
  reg reg_act_regs_data_0_11_2_enexo_3;
  reg reg_act_config_inst_counter_enexo_49;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_50;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_50;
  reg reg_act_regs_data_2_0_2_enexo_3;
  reg reg_act_regs_data_3_0_2_enexo_3;
  reg reg_act_regs_data_1_0_2_enexo_3;
  reg reg_act_regs_data_0_0_2_enexo_3;
  reg reg_act_config_inst_counter_enexo_50;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_51;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_51;
  reg reg_act_regs_data_1_1_2_enexo_3;
  reg reg_act_regs_data_3_1_2_enexo_3;
  reg reg_act_regs_data_0_1_2_enexo_3;
  reg reg_act_regs_data_2_1_2_enexo_3;
  reg reg_act_config_inst_counter_enexo_51;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_52;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_52;
  reg reg_act_regs_data_2_3_2_enexo_3;
  reg reg_act_regs_data_3_3_2_enexo_3;
  reg reg_act_regs_data_1_3_2_enexo_3;
  reg reg_act_regs_data_0_3_2_enexo_3;
  reg reg_act_config_inst_counter_enexo_52;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_53;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_53;
  reg reg_act_regs_data_2_4_2_enexo_3;
  reg reg_act_regs_data_3_4_2_enexo_3;
  reg reg_act_regs_data_1_4_2_enexo_3;
  reg reg_act_regs_data_0_4_2_enexo_3;
  reg reg_act_config_inst_counter_enexo_53;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_54;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_54;
  reg reg_act_regs_data_0_5_2_enexo_3;
  reg reg_act_regs_data_2_5_2_enexo_3;
  reg reg_act_regs_data_3_5_2_enexo_3;
  reg reg_act_regs_data_1_5_2_enexo_3;
  reg reg_act_config_inst_counter_enexo_54;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_55;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_55;
  reg reg_act_regs_data_3_6_2_enexo_3;
  reg reg_act_regs_data_1_6_2_enexo_3;
  reg reg_act_regs_data_0_6_2_enexo_3;
  reg reg_act_regs_data_2_6_2_enexo_3;
  reg reg_act_config_inst_counter_enexo_55;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_56;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_56;
  reg reg_act_regs_data_2_7_2_enexo_3;
  reg reg_act_regs_data_1_7_2_enexo_3;
  reg reg_act_regs_data_0_7_2_enexo_3;
  reg reg_act_regs_data_3_7_2_enexo_3;
  reg reg_act_config_inst_counter_enexo_56;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_57;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_57;
  reg reg_act_regs_data_3_8_2_enexo_3;
  reg reg_act_regs_data_1_8_2_enexo_3;
  reg reg_act_regs_data_0_8_2_enexo_3;
  reg reg_act_regs_data_2_8_2_enexo_3;
  reg reg_act_config_inst_counter_enexo_57;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_58;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_58;
  reg reg_act_regs_data_1_9_2_enexo_3;
  reg reg_act_regs_data_0_9_2_enexo_3;
  reg reg_act_regs_data_2_9_2_enexo_3;
  reg reg_act_regs_data_3_9_2_enexo_3;
  reg reg_act_config_inst_counter_enexo_58;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_59;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_59;
  reg reg_act_regs_data_0_10_2_enexo_3;
  reg reg_act_regs_data_1_10_2_enexo_3;
  reg reg_act_regs_data_2_10_2_enexo_3;
  reg reg_act_regs_data_3_10_2_enexo_3;
  reg reg_act_config_inst_counter_enexo_59;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_60;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_60;
  reg reg_act_regs_data_1_12_2_enexo_3;
  reg reg_act_regs_data_2_12_2_enexo_3;
  reg reg_act_regs_data_0_12_2_enexo_3;
  reg reg_act_regs_data_3_12_2_enexo_3;
  reg reg_act_config_inst_counter_enexo_60;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_61;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_61;
  reg reg_act_regs_data_1_13_2_enexo_3;
  reg reg_act_regs_data_0_13_2_enexo_3;
  reg reg_act_regs_data_3_13_2_enexo_3;
  reg reg_act_regs_data_2_13_2_enexo_3;
  reg reg_act_config_inst_counter_enexo_61;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_62;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_62;
  reg reg_act_regs_data_3_14_2_enexo_3;
  reg reg_act_regs_data_0_14_2_enexo_3;
  reg reg_act_regs_data_1_14_2_enexo_3;
  reg reg_act_regs_data_2_14_2_enexo_3;
  reg reg_act_config_inst_counter_enexo_62;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_63;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_63;
  reg reg_act_regs_data_1_15_2_enexo_3;
  reg reg_act_regs_data_2_15_2_enexo_3;
  reg reg_act_regs_data_0_15_2_enexo_3;
  reg reg_act_config_inst_counter_enexo_63;
  reg reg_act_regs_data_3_15_2_enexo_3;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_64;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_64;
  reg reg_act_config_inst_counter_enexo_64;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_65;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_65;
  reg reg_act_regs_data_2_0_2_enexo_4;
  reg reg_act_regs_data_3_0_2_enexo_4;
  reg reg_act_regs_data_1_0_2_enexo_4;
  reg reg_act_regs_data_0_0_2_enexo_4;
  reg reg_act_config_inst_counter_enexo_65;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_66;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_66;
  reg reg_act_regs_data_1_1_2_enexo_4;
  reg reg_act_regs_data_3_1_2_enexo_4;
  reg reg_act_regs_data_0_1_2_enexo_4;
  reg reg_act_regs_data_2_1_2_enexo_4;
  reg reg_act_config_inst_counter_enexo_66;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_67;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_67;
  reg reg_act_regs_data_0_2_2_enexo_4;
  reg reg_act_regs_data_2_2_2_enexo_4;
  reg reg_act_regs_data_1_2_2_enexo_4;
  reg reg_act_regs_data_3_2_2_enexo_4;
  reg reg_act_config_inst_counter_enexo_67;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_68;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_68;
  reg reg_act_regs_data_2_3_2_enexo_4;
  reg reg_act_regs_data_3_3_2_enexo_4;
  reg reg_act_regs_data_1_3_2_enexo_4;
  reg reg_act_regs_data_0_3_2_enexo_4;
  reg reg_act_config_inst_counter_enexo_68;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_69;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_69;
  reg reg_act_regs_data_2_4_2_enexo_4;
  reg reg_act_regs_data_3_4_2_enexo_4;
  reg reg_act_regs_data_1_4_2_enexo_4;
  reg reg_act_regs_data_0_4_2_enexo_4;
  reg reg_act_config_inst_counter_enexo_69;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_70;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_70;
  reg reg_act_regs_data_0_5_2_enexo_4;
  reg reg_act_regs_data_2_5_2_enexo_4;
  reg reg_act_regs_data_3_5_2_enexo_4;
  reg reg_act_regs_data_1_5_2_enexo_4;
  reg reg_act_config_inst_counter_enexo_70;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_71;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_71;
  reg reg_act_regs_data_3_6_2_enexo_4;
  reg reg_act_regs_data_1_6_2_enexo_4;
  reg reg_act_regs_data_0_6_2_enexo_4;
  reg reg_act_regs_data_2_6_2_enexo_4;
  reg reg_act_config_inst_counter_enexo_71;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_72;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_72;
  reg reg_act_regs_data_2_7_2_enexo_4;
  reg reg_act_regs_data_1_7_2_enexo_4;
  reg reg_act_regs_data_0_7_2_enexo_4;
  reg reg_act_regs_data_3_7_2_enexo_4;
  reg reg_act_config_inst_counter_enexo_72;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_73;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_73;
  reg reg_act_regs_data_3_8_2_enexo_4;
  reg reg_act_regs_data_1_8_2_enexo_4;
  reg reg_act_regs_data_0_8_2_enexo_4;
  reg reg_act_regs_data_2_8_2_enexo_4;
  reg reg_act_config_inst_counter_enexo_73;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_74;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_74;
  reg reg_act_regs_data_2_11_2_enexo_4;
  reg reg_act_regs_data_3_11_2_enexo_4;
  reg reg_act_regs_data_1_11_2_enexo_4;
  reg reg_act_regs_data_0_11_2_enexo_4;
  reg reg_act_config_inst_counter_enexo_74;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_75;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_75;
  reg reg_act_regs_data_1_12_2_enexo_4;
  reg reg_act_regs_data_2_12_2_enexo_4;
  reg reg_act_regs_data_0_12_2_enexo_4;
  reg reg_act_regs_data_3_12_2_enexo_4;
  reg reg_act_config_inst_counter_enexo_75;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_76;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_76;
  reg reg_act_regs_data_1_13_2_enexo_4;
  reg reg_act_regs_data_0_13_2_enexo_4;
  reg reg_act_regs_data_3_13_2_enexo_4;
  reg reg_act_regs_data_2_13_2_enexo_4;
  reg reg_act_config_inst_counter_enexo_76;
  reg reg_act_config_inst_regs_1_sva_dfm_5_enexo_77;
  reg reg_act_config_inst_regs_17_sva_dfm_6_enexo_77;
  reg reg_act_regs_data_3_14_2_enexo_4;
  reg reg_act_regs_data_0_14_2_enexo_4;
  reg reg_act_regs_data_1_14_2_enexo_4;
  reg reg_act_regs_data_2_14_2_enexo_4;
  reg reg_act_config_inst_counter_enexo_77;
  wire act_regs_data_and_859_enex5;
  wire act_regs_data_and_860_enex5;
  wire act_regs_data_and_861_enex5;
  wire act_regs_data_and_862_enex5;
  wire act_regs_data_and_863_enex5;
  wire act_regs_data_and_864_enex5;
  wire act_regs_data_and_865_enex5;
  wire act_regs_data_and_866_enex5;
  wire act_regs_data_and_867_enex5;
  wire act_regs_data_and_868_enex5;
  wire act_regs_data_and_869_enex5;
  wire act_regs_data_and_870_enex5;
  wire act_regs_data_and_871_enex5;
  wire act_regs_data_and_872_enex5;
  wire act_regs_data_and_873_enex5;
  wire act_regs_data_and_874_enex5;
  wire act_regs_data_and_875_enex5;
  wire act_regs_data_and_876_enex5;
  wire act_regs_data_and_877_enex5;
  wire act_regs_data_and_878_enex5;
  wire act_regs_data_and_879_enex5;
  wire act_regs_data_and_880_enex5;
  wire act_regs_data_and_881_enex5;
  wire act_regs_data_and_882_enex5;
  wire act_regs_data_and_883_enex5;
  wire act_regs_data_and_884_enex5;
  wire act_regs_data_and_885_enex5;
  wire act_regs_data_and_886_enex5;
  wire act_regs_data_and_887_enex5;
  wire act_regs_data_and_888_enex5;
  wire act_regs_data_and_889_enex5;
  wire act_regs_data_and_890_enex5;
  wire act_regs_data_and_891_enex5;
  wire act_regs_data_and_892_enex5;
  wire act_regs_data_and_893_enex5;
  wire act_regs_data_and_894_enex5;
  wire act_regs_data_and_895_enex5;
  wire act_regs_data_and_896_enex5;
  wire act_regs_data_and_897_enex5;
  wire act_regs_data_and_898_enex5;
  wire act_regs_data_and_899_enex5;
  wire act_regs_data_and_900_enex5;
  wire act_regs_data_and_901_enex5;
  wire act_regs_data_and_902_enex5;
  wire act_regs_data_and_903_enex5;
  wire act_regs_data_and_904_enex5;
  wire act_regs_data_and_905_enex5;
  wire act_regs_data_and_906_enex5;
  wire act_regs_data_and_907_enex5;
  wire act_regs_data_and_908_enex5;
  wire act_regs_data_and_909_enex5;
  wire act_regs_data_and_910_enex5;
  wire act_regs_data_and_911_enex5;
  wire act_regs_data_and_912_enex5;
  wire act_regs_data_and_913_enex5;
  wire act_regs_data_and_914_enex5;
  wire act_regs_data_and_915_enex5;
  wire act_regs_data_and_916_enex5;
  wire act_regs_data_and_917_enex5;
  wire act_regs_data_and_918_enex5;
  wire act_regs_data_and_919_enex5;
  wire act_regs_data_and_920_enex5;
  wire act_regs_data_and_921_enex5;
  wire act_regs_data_and_922_enex5;
  wire act_mem_banks_read_read_data_and_16_enex5;
  wire act_mem_banks_read_read_data_and_17_enex5;
  wire act_mem_banks_read_read_data_and_18_enex5;
  wire act_mem_banks_read_read_data_and_19_enex5;
  wire act_mem_banks_read_read_data_and_20_enex5;
  wire act_mem_banks_read_read_data_and_21_enex5;
  wire act_mem_banks_read_read_data_and_22_enex5;
  wire act_mem_banks_read_read_data_and_23_enex5;
  wire act_mem_banks_read_read_data_and_24_enex5;
  wire act_mem_banks_read_read_data_and_25_enex5;
  wire act_mem_banks_read_read_data_and_26_enex5;
  wire act_mem_banks_read_read_data_and_27_enex5;
  wire act_mem_banks_read_read_data_and_28_enex5;
  wire act_mem_banks_read_read_data_and_29_enex5;
  wire act_mem_banks_read_read_data_and_30_enex5;
  wire act_mem_banks_read_read_data_and_31_enex5;
  wire act_port_read_out_data_and_16_enex5;
  wire act_port_read_out_data_and_17_enex5;
  wire act_port_read_out_data_and_18_enex5;
  wire act_port_read_out_data_and_19_enex5;
  wire act_port_read_out_data_and_20_enex5;
  wire act_port_read_out_data_and_21_enex5;
  wire act_port_read_out_data_and_22_enex5;
  wire act_port_read_out_data_and_23_enex5;
  wire act_port_read_out_data_and_24_enex5;
  wire act_port_read_out_data_and_25_enex5;
  wire act_port_read_out_data_and_26_enex5;
  wire act_port_read_out_data_and_27_enex5;
  wire act_port_read_out_data_and_28_enex5;
  wire act_port_read_out_data_and_29_enex5;
  wire act_port_read_out_data_and_30_enex5;
  wire act_port_read_out_data_and_31_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_37_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_38_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_39_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_40_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_41_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_42_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_43_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_44_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_45_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_46_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_47_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_48_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_49_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_50_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_51_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_52_enex5;
  wire Relu_for_y_qelse_and_31_enex5;
  wire Relu_for_y_qelse_and_32_enex5;
  wire Relu_for_y_qelse_and_33_enex5;
  wire Relu_for_y_qelse_and_34_enex5;
  wire Relu_for_y_qelse_and_35_enex5;
  wire Relu_for_y_qelse_and_36_enex5;
  wire Relu_for_y_qelse_and_37_enex5;
  wire Relu_for_y_qelse_and_38_enex5;
  wire Relu_for_y_qelse_and_39_enex5;
  wire Relu_for_y_qelse_and_40_enex5;
  wire Relu_for_y_qelse_and_41_enex5;
  wire Relu_for_y_qelse_and_42_enex5;
  wire Relu_for_y_qelse_and_43_enex5;
  wire Relu_for_y_qelse_and_44_enex5;
  wire Relu_for_y_qelse_and_45_enex5;
  wire Relu_for_y_qelse_and_46_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_15_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_16_enex5;
  wire ActUnit_RunInst_switch_lp_and_815_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_17_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_18_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_19_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_20_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_21_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_22_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_23_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_24_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_25_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_26_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_27_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_28_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_29_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_15_enex5;
  wire ActUnit_RunInst_switch_lp_and_816_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_16_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_17_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_18_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_19_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_20_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_21_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_22_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_23_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_24_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_25_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_26_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_27_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_28_enex5;
  wire ActUnit_RunInst_curr_inst_and_enex5;
  wire ActUnit_RunInst_switch_lp_and_817_enex5;
  wire nv_scvector_cctor_nv_scvector_3_for_and_enex5;
  wire nv_scvector_cctor_nv_scvector_3_for_and_15_enex5;
  wire nv_scvector_cctor_nv_scvector_3_for_and_16_enex5;
  wire nv_scvector_cctor_nv_scvector_3_for_and_17_enex5;
  wire nv_scvector_cctor_nv_scvector_3_for_and_18_enex5;
  wire nv_scvector_cctor_nv_scvector_3_for_and_19_enex5;
  wire nv_scvector_cctor_nv_scvector_3_for_and_20_enex5;
  wire nv_scvector_cctor_nv_scvector_3_for_and_21_enex5;
  wire nv_scvector_cctor_nv_scvector_3_for_and_22_enex5;
  wire nv_scvector_cctor_nv_scvector_3_for_and_23_enex5;
  wire nv_scvector_cctor_nv_scvector_3_for_and_24_enex5;
  wire nv_scvector_cctor_nv_scvector_3_for_and_25_enex5;
  wire w_load_and_tmp;
  wire is_start_and_tmp;
  wire and_1417_tmp;
  wire and_1415_tmp;
  wire and_1413_tmp;
  wire and_1411_tmp;
  wire and_1409_tmp;
  wire and_1407_tmp;
  wire and_1405_tmp;
  wire and_1403_tmp;
  wire and_1401_tmp;
  wire and_1399_tmp;
  wire and_1397_tmp;
  wire and_1395_tmp;
  wire and_1393_tmp;
  wire and_1391_tmp;
  wire and_1389_tmp;
  wire and_1387_tmp;
  wire and_1385_tmp;
  wire and_1383_tmp;
  wire and_1381_tmp;
  wire and_1379_tmp;
  wire and_1377_tmp;
  wire and_1375_tmp;
  wire and_1373_tmp;
  wire and_1371_tmp;
  wire and_1369_tmp;
  wire and_1367_tmp;
  wire and_1365_tmp;
  wire and_1363_tmp;
  wire and_1361_tmp;
  wire and_1359_tmp;
  wire and_1357_tmp;
  wire and_1355_tmp;
  wire and_1353_tmp;
  wire and_1351_tmp;
  wire and_1349_tmp;
  wire and_1347_tmp;
  wire and_1345_tmp;
  wire and_1343_tmp;
  wire and_1341_tmp;
  wire and_1339_tmp;
  wire and_1337_tmp;
  wire and_1335_tmp;
  wire and_1333_tmp;
  wire and_1331_tmp;
  wire and_1329_tmp;
  wire and_1327_tmp;
  wire and_1325_tmp;
  wire and_1323_tmp;
  wire and_1246_tmp;
  wire and_1321_tmp;
  wire and_1243_tmp;
  wire and_1319_tmp;
  wire and_1237_tmp;
  wire and_1317_tmp;
  wire and_1231_tmp;
  wire and_1315_tmp;
  wire and_1275_tmp;
  wire and_1313_tmp;
  wire and_1268_tmp;
  wire and_1311_tmp;
  wire and_1309_tmp;
  wire and_1240_tmp;
  wire and_1307_tmp;
  wire and_1234_tmp;
  wire and_1305_tmp;
  wire and_1228_tmp;
  wire and_1303_tmp;
  wire and_1289_tmp;
  wire and_1301_tmp;
  wire and_1282_tmp;
  wire and_1299_tmp;
  wire and_1254_tmp;
  wire and_1297_tmp;
  wire and_1250_tmp;
  wire and_1295_tmp;
  wire and_1261_tmp;
  wire and_1293_tmp;
  wire and_1225_tmp;
  wire and_1291_tmp;
  wire ActUnit_CheckStart_start_reg_and_tmp;
  wire act_config_inst_counter_and_tmp;
  wire or_71_cse;
  wire [31:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_22_itm;
  wire ActUnit_PushOutput_if_for_and_27_itm;
  wire [28:0] Silu_for_1_else_else_acc_itm_29_1;
  wire [27:0] Gelu_for_13_else_else_acc_itm_28_1;
  wire [27:0] Gelu_for_8_else_else_acc_itm_28_1;
  wire Tanh_for_else_else_and_8_cse;
  wire Tanh_for_else_else_and_9_cse;
  wire [27:0] z_out_28_1;
  wire [27:0] z_out_1_28_1;
  wire [27:0] z_out_2_28_1;
  wire [28:0] z_out_3_29_1;
  wire [28:0] z_out_4_29_1;

  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_1;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_1;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_1;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_1;
  wire mux_114_nl;
  wire nand_6_nl;
  wire mux_113_nl;
  wire mux_112_nl;
  wire mux_111_nl;
  wire nand_5_nl;
  wire or_443_nl;
  wire mux_110_nl;
  wire or_442_nl;
  wire mux_109_nl;
  wire mux_108_nl;
  wire mux_107_nl;
  wire nand_4_nl;
  wire mux_106_nl;
  wire mux_105_nl;
  wire and_603_nl;
  wire and_602_nl;
  wire mux_104_nl;
  wire and_601_nl;
  wire and_600_nl;
  wire mux_103_nl;
  wire mux_102_nl;
  wire nand_2_nl;
  wire mux_100_nl;
  wire mux_99_nl;
  wire and_598_nl;
  wire mux_98_nl;
  wire and_596_nl;
  wire and_595_nl;
  wire nand_1_nl;
  wire mux_97_nl;
  wire nor_160_nl;
  wire mux_96_nl;
  wire and_594_nl;
  wire mux_95_nl;
  wire or_419_nl;
  wire or_417_nl;
  wire nor_161_nl;
  wire mux_134_nl;
  wire nand_12_nl;
  wire mux_133_nl;
  wire mux_132_nl;
  wire mux_131_nl;
  wire nand_11_nl;
  wire or_471_nl;
  wire mux_130_nl;
  wire or_470_nl;
  wire mux_129_nl;
  wire mux_128_nl;
  wire mux_127_nl;
  wire nand_10_nl;
  wire mux_126_nl;
  wire mux_125_nl;
  wire and_615_nl;
  wire and_614_nl;
  wire mux_124_nl;
  wire and_613_nl;
  wire and_612_nl;
  wire mux_123_nl;
  wire mux_122_nl;
  wire nand_8_nl;
  wire mux_120_nl;
  wire mux_119_nl;
  wire and_610_nl;
  wire and_609_nl;
  wire mux_118_nl;
  wire and_608_nl;
  wire and_607_nl;
  wire nand_7_nl;
  wire mux_117_nl;
  wire nor_162_nl;
  wire mux_116_nl;
  wire and_606_nl;
  wire mux_115_nl;
  wire or_447_nl;
  wire or_445_nl;
  wire nor_163_nl;
  wire mux_140_nl;
  wire mux_139_nl;
  wire mux_138_nl;
  wire or_477_nl;
  wire or_476_nl;
  wire mux_137_nl;
  wire mux_136_nl;
  wire mux_135_nl;
  wire or_475_nl;
  wire or_474_nl;
  wire or_472_nl;
  wire mux_141_nl;
  wire nor_164_nl;
  wire nor_165_nl;
  wire mux_151_nl;
  wire or_499_nl;
  wire mux_150_nl;
  wire or_497_nl;
  wire mux_149_nl;
  wire or_496_nl;
  wire mux_148_nl;
  wire mux_147_nl;
  wire mux_146_nl;
  wire nand_207_nl;
  wire mux_145_nl;
  wire and_631_nl;
  wire mux_144_nl;
  wire nor_167_nl;
  wire mux_143_nl;
  wire mux_142_nl;
  wire or_485_nl;
  wire or_484_nl;
  wire or_481_nl;
  wire mux_165_nl;
  wire nor_171_nl;
  wire mux_164_nl;
  wire nor_172_nl;
  wire mux_163_nl;
  wire or_522_nl;
  wire mux_162_nl;
  wire mux_161_nl;
  wire mux_160_nl;
  wire mux_159_nl;
  wire nor_170_nl;
  wire nand_209_nl;
  wire nand_210_nl;
  wire mux_158_nl;
  wire mux_157_nl;
  wire mux_156_nl;
  wire and_655_nl;
  wire mux_155_nl;
  wire mux_154_nl;
  wire mux_153_nl;
  wire and_651_nl;
  wire and_649_nl;
  wire and_647_nl;
  wire or_504_nl;
  wire mux_179_nl;
  wire nor_197_nl;
  wire mux_178_nl;
  wire nor_198_nl;
  wire mux_177_nl;
  wire or_542_nl;
  wire mux_176_nl;
  wire mux_175_nl;
  wire mux_174_nl;
  wire mux_173_nl;
  wire nor_195_nl;
  wire nand_211_nl;
  wire nand_212_nl;
  wire mux_172_nl;
  wire mux_171_nl;
  wire mux_170_nl;
  wire mux_168_nl;
  wire mux_167_nl;
  wire mux_166_nl;
  wire nor_196_nl;
  wire and_706_nl;
  wire or_526_nl;
  wire mux_180_nl;
  wire nor_199_nl;
  wire nor_200_nl;
  wire mux_181_nl;
  wire nor_201_nl;
  wire nor_202_nl;
  wire mux_182_nl;
  wire nor_203_nl;
  wire nor_204_nl;
  wire mux_183_nl;
  wire nor_205_nl;
  wire nor_206_nl;
  wire mux_184_nl;
  wire nor_207_nl;
  wire nor_208_nl;
  wire mux_185_nl;
  wire nor_209_nl;
  wire nor_210_nl;
  wire mux_186_nl;
  wire nor_211_nl;
  wire nor_212_nl;
  wire mux_187_nl;
  wire nor_213_nl;
  wire nor_214_nl;
  wire mux_188_nl;
  wire nor_215_nl;
  wire nor_216_nl;
  wire mux_189_nl;
  wire nor_217_nl;
  wire nor_218_nl;
  wire mux_190_nl;
  wire nor_219_nl;
  wire nor_220_nl;
  wire mux_191_nl;
  wire nor_221_nl;
  wire nor_222_nl;
  wire mux_192_nl;
  wire nor_223_nl;
  wire nor_224_nl;
  wire mux_193_nl;
  wire nor_225_nl;
  wire nor_226_nl;
  wire and_843_nl;
  wire mux_53_nl;
  wire mux_52_nl;
  wire nor_62_nl;
  wire or_172_nl;
  wire nor_18_nl;
  wire while_else_1_while_else_1_nand_1_nl;
  wire mux_80_nl;
  wire nor_74_nl;
  wire mux_79_nl;
  wire or_242_nl;
  wire mux_78_nl;
  wire mux_77_nl;
  wire or_240_nl;
  wire mux_76_nl;
  wire mux_75_nl;
  wire nor_347_nl;
  wire or_238_nl;
  wire[7:0] act_config_InstIncr_if_act_config_InstIncr_if_and_1_nl;
  wire[7:0] operator_8_false_acc_nl;
  wire[8:0] nl_operator_8_false_acc_nl;
  wire act_config_InstIncr_if_not_nl;
  wire[4:0] act_config_InstIncr_act_config_InstIncr_and_1_nl;
  wire[4:0] operator_5_false_acc_nl;
  wire[5:0] nl_operator_5_false_acc_nl;
  wire act_config_InstIncr_if_not_7_nl;
  wire and_880_nl;
  wire mux_296_nl;
  wire and_1426_nl;
  wire mux_295_nl;
  wire mux_294_nl;
  wire mux_293_nl;
  wire mux_292_nl;
  wire mux_291_nl;
  wire nor_678_nl;
  wire nor_679_nl;
  wire mux_290_nl;
  wire nor_680_nl;
  wire nor_681_nl;
  wire mux_289_nl;
  wire mux_288_nl;
  wire nor_682_nl;
  wire nor_683_nl;
  wire mux_287_nl;
  wire nor_684_nl;
  wire nor_685_nl;
  wire mux_286_nl;
  wire mux_285_nl;
  wire mux_284_nl;
  wire nor_686_nl;
  wire nor_687_nl;
  wire mux_283_nl;
  wire nor_688_nl;
  wire nor_689_nl;
  wire mux_282_nl;
  wire mux_281_nl;
  wire nor_690_nl;
  wire nor_691_nl;
  wire mux_280_nl;
  wire nor_692_nl;
  wire nor_693_nl;
  wire mux_279_nl;
  wire mux_278_nl;
  wire mux_277_nl;
  wire mux_276_nl;
  wire nor_694_nl;
  wire nor_695_nl;
  wire mux_275_nl;
  wire nor_696_nl;
  wire nor_697_nl;
  wire mux_274_nl;
  wire mux_273_nl;
  wire nor_698_nl;
  wire nor_699_nl;
  wire mux_272_nl;
  wire nor_700_nl;
  wire nor_701_nl;
  wire mux_271_nl;
  wire mux_270_nl;
  wire mux_269_nl;
  wire nor_702_nl;
  wire nor_703_nl;
  wire mux_268_nl;
  wire nor_704_nl;
  wire nor_705_nl;
  wire mux_267_nl;
  wire mux_266_nl;
  wire nor_706_nl;
  wire nor_707_nl;
  wire mux_nl;
  wire nor_708_nl;
  wire nor_709_nl;
  wire nor_nl;
  wire mux_199_nl;
  wire mux_198_nl;
  wire mux_298_nl;
  wire mux_297_nl;
  wire and_nl;
  wire nor_710_nl;
  wire nor_711_nl;
  wire[31:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_13_nl;
  wire[31:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_12_nl;
  wire[31:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_11_nl;
  wire[31:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_10_nl;
  wire[31:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_9_nl;
  wire[31:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_8_nl;
  wire[31:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_7_nl;
  wire[31:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_6_nl;
  wire[31:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_5_nl;
  wire[31:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_4_nl;
  wire[31:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_3_nl;
  wire[31:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_nl;
  wire mux_202_nl;
  wire mux_201_nl;
  wire mux_200_nl;
  wire and_1094_nl;
  wire[7:0] and_1111_nl;
  wire[7:0] mux_252_nl;
  wire not_1290_nl;
  wire[7:0] and_1113_nl;
  wire[7:0] mux_253_nl;
  wire not_1292_nl;
  wire[7:0] and_1115_nl;
  wire[7:0] mux_254_nl;
  wire not_1294_nl;
  wire[7:0] and_1117_nl;
  wire[7:0] mux_255_nl;
  wire not_1296_nl;
  wire[7:0] and_1119_nl;
  wire[7:0] mux_256_nl;
  wire not_1298_nl;
  wire[7:0] and_1121_nl;
  wire[7:0] mux_257_nl;
  wire not_1300_nl;
  wire[7:0] and_1123_nl;
  wire[7:0] mux_258_nl;
  wire not_1302_nl;
  wire[7:0] and_1125_nl;
  wire[7:0] mux_259_nl;
  wire not_1304_nl;
  wire[7:0] and_1127_nl;
  wire[7:0] mux_260_nl;
  wire not_1306_nl;
  wire[7:0] and_1129_nl;
  wire[7:0] mux_261_nl;
  wire not_1308_nl;
  wire[1:0] and_1131_nl;
  wire[1:0] mux_262_nl;
  wire not_1310_nl;
  wire[6:0] and_1133_nl;
  wire[6:0] mux_263_nl;
  wire not_1312_nl;
  wire[6:0] and_1135_nl;
  wire[6:0] mux_264_nl;
  wire not_1314_nl;
  wire[2:0] and_1137_nl;
  wire[2:0] mux_265_nl;
  wire not_1316_nl;
  wire ActUnit_RunInst_switch_lp_mux_1_nl;
  wire ActUnit_RunInst_switch_lp_mux_2_nl;
  wire ActUnit_RunInst_switch_lp_mux_4_nl;
  wire ActUnit_RunInst_switch_lp_mux_5_nl;
  wire ActUnit_RunInst_switch_lp_mux_7_nl;
  wire ActUnit_RunInst_switch_lp_mux_9_nl;
  wire ActUnit_RunInst_switch_lp_mux_11_nl;
  wire ActUnit_RunInst_switch_lp_mux_13_nl;
  wire mux_204_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_14_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_13_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_12_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_11_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_10_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_9_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_8_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_7_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_6_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_5_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_4_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_3_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_2_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_1_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_nl;
  wire ActUnit_RunInst_switch_lp_not_1_nl;
  wire mux_206_nl;
  wire mux_208_nl;
  wire mux_207_nl;
  wire mux_209_nl;
  wire and_1096_nl;
  wire mux_210_nl;
  wire mux_211_nl;
  wire ActUnit_RunInst_switch_lp_or_3_nl;
  wire ActUnit_PushOutput_if_for_i_not_nl;
  wire mux_213_nl;
  wire nor_232_nl;
  wire reg_act_regs_data_0_0_1_rgt_nl;
  wire act_regs_data_nor_1_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_68_nl;
  wire[30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_141_nl;
  wire reg_act_regs_data_0_1_1_rgt_nl;
  wire act_regs_data_or_1_nl;
  wire act_regs_data_mux1h_74_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_4_nl;
  wire[30:0] act_regs_data_mux1h_575_nl;
  wire not_3696_nl;
  wire reg_act_regs_data_0_10_1_rgt_nl;
  wire act_regs_data_or_2_nl;
  wire act_regs_data_mux1h_79_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_11_nl;
  wire[30:0] act_regs_data_mux1h_567_nl;
  wire not_3697_nl;
  wire reg_act_regs_data_0_11_1_rgt_nl;
  wire act_regs_data_or_4_nl;
  wire act_regs_data_mux1h_84_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_73_nl;
  wire[30:0] act_regs_data_mux1h_566_nl;
  wire not_3698_nl;
  wire reg_act_regs_data_0_12_1_rgt_nl;
  wire act_regs_data_or_6_nl;
  wire act_regs_data_mux1h_89_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_80_nl;
  wire[30:0] act_regs_data_mux1h_565_nl;
  wire not_3699_nl;
  wire reg_act_regs_data_0_13_1_rgt_nl;
  wire act_regs_data_or_8_nl;
  wire act_regs_data_mux1h_94_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_87_nl;
  wire[30:0] act_regs_data_mux1h_564_nl;
  wire not_3700_nl;
  wire reg_act_regs_data_0_14_1_rgt_nl;
  wire act_regs_data_or_10_nl;
  wire act_regs_data_mux1h_99_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_94_nl;
  wire[30:0] act_regs_data_mux1h_563_nl;
  wire not_3701_nl;
  wire reg_act_regs_data_0_15_1_rgt_nl;
  wire act_regs_data_or_12_nl;
  wire act_regs_data_mux1h_104_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_101_nl;
  wire[30:0] act_regs_data_mux1h_562_nl;
  wire not_3702_nl;
  wire reg_act_regs_data_0_2_1_rgt_nl;
  wire act_regs_data_or_14_nl;
  wire act_regs_data_mux1h_109_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_108_nl;
  wire[30:0] act_regs_data_mux1h_574_nl;
  wire not_3703_nl;
  wire reg_act_regs_data_0_3_1_rgt_nl;
  wire act_regs_data_or_16_nl;
  wire act_regs_data_mux1h_114_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_18_nl;
  wire[30:0] act_regs_data_mux1h_573_nl;
  wire not_3704_nl;
  wire reg_act_regs_data_0_4_1_rgt_nl;
  wire act_regs_data_or_18_nl;
  wire act_regs_data_mux1h_119_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_25_nl;
  wire[30:0] act_regs_data_mux1h_572_nl;
  wire not_3705_nl;
  wire reg_act_regs_data_0_5_1_rgt_nl;
  wire act_regs_data_or_20_nl;
  wire act_regs_data_mux1h_124_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_32_nl;
  wire[30:0] act_regs_data_mux1h_571_nl;
  wire not_3706_nl;
  wire reg_act_regs_data_0_6_1_rgt_nl;
  wire act_regs_data_or_22_nl;
  wire act_regs_data_mux1h_129_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_39_nl;
  wire[30:0] act_regs_data_mux1h_570_nl;
  wire not_3707_nl;
  wire reg_act_regs_data_0_7_1_rgt_nl;
  wire act_regs_data_or_24_nl;
  wire act_regs_data_mux1h_134_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_46_nl;
  wire[30:0] act_regs_data_mux1h_569_nl;
  wire not_3708_nl;
  wire reg_act_regs_data_0_8_1_rgt_nl;
  wire act_regs_data_or_26_nl;
  wire act_regs_data_mux1h_139_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_53_nl;
  wire[30:0] act_regs_data_mux1h_568_nl;
  wire not_3709_nl;
  wire ActUnit_RunInst_case_2_for_ActUnit_RunInst_case_2_for_and_nl;
  wire Gelu_for_Gelu_for_and_11_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_6_nl;
  wire[30:0] ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_90_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_and_34_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_and_35_nl;
  wire nor_771_nl;
  wire nor_340_nl;
  wire and_1140_nl;
  wire mux_217_nl;
  wire ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_5_nl;
  wire ActUnit_DecodeAxiRead_else_mux_1_nl;
  wire mux_218_nl;
  wire ActUnit_DecodeAxi_mux_93_nl;
  wire ActUnit_DecodeAxi_if_mux_91_nl;
  wire ActUnit_DecodeAxiRead_mux_33_nl;
  wire act_config_ActConfigRead_mux_19_nl;
  wire act_config_ActConfigRead_else_mux_19_nl;
  wire act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_24_nl;
  wire ActUnit_DecodeAxi_mux_94_nl;
  wire ActUnit_DecodeAxi_if_mux_89_nl;
  wire ActUnit_DecodeAxiRead_mux_31_nl;
  wire act_config_ActConfigRead_mux_17_nl;
  wire act_config_ActConfigRead_else_mux_17_nl;
  wire act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_18_nl;
  wire[5:0] act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_20_nl;
  wire[7:0] act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_21_nl;
  wire[4:0] act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_22_nl;
  wire[7:0] act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_23_nl;
  wire mux_219_nl;
  wire mux_220_nl;
  wire or_829_nl;
  wire or_997_nl;
  wire[1:0] ActUnit_DecodeAxiWrite_if_mux_5_nl;
  wire[1:0] ActUnit_DecodeAxiWrite_if_mux_7_nl;
  wire[1:0] ActUnit_DecodeAxiWrite_if_mux_9_nl;
  wire[1:0] ActUnit_DecodeAxiWrite_if_mux_11_nl;
  wire[1:0] ActUnit_DecodeAxiWrite_if_mux_13_nl;
  wire[1:0] ActUnit_DecodeAxiWrite_if_mux_15_nl;
  wire[1:0] ActUnit_DecodeAxiWrite_if_mux_17_nl;
  wire[1:0] ActUnit_DecodeAxiWrite_if_mux_19_nl;
  wire[1:0] ActUnit_DecodeAxiWrite_if_mux_21_nl;
  wire[1:0] ActUnit_DecodeAxiWrite_if_mux_23_nl;
  wire[1:0] ActUnit_DecodeAxiWrite_if_mux_25_nl;
  wire[1:0] ActUnit_DecodeAxiWrite_if_mux_27_nl;
  wire[1:0] ActUnit_DecodeAxiWrite_if_mux_29_nl;
  wire[1:0] ActUnit_DecodeAxiWrite_if_mux_31_nl;
  wire[1:0] ActUnit_DecodeAxiWrite_if_mux_33_nl;
  wire[1:0] ActUnit_DecodeAxiWrite_if_mux_35_nl;
  wire act_regs_data_mux_128_nl;
  wire act_regs_data_or_126_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_69_nl;
  wire[30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_174_nl;
  wire act_regs_data_mux_129_nl;
  wire act_regs_data_or_127_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_104_nl;
  wire[30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_173_nl;
  wire act_regs_data_mux_130_nl;
  wire act_regs_data_or_128_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_97_nl;
  wire[30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_171_nl;
  wire act_regs_data_mux_131_nl;
  wire act_regs_data_or_129_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_90_nl;
  wire[30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_169_nl;
  wire act_regs_data_mux_132_nl;
  wire act_regs_data_or_130_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_83_nl;
  wire[30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_167_nl;
  wire act_regs_data_mux_133_nl;
  wire act_regs_data_or_131_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_76_nl;
  wire[30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_165_nl;
  wire act_regs_data_mux_134_nl;
  wire act_regs_data_or_132_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_12_nl;
  wire[30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_163_nl;
  wire act_regs_data_mux_135_nl;
  wire act_regs_data_or_133_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_62_nl;
  wire[30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_161_nl;
  wire act_regs_data_mux_136_nl;
  wire act_regs_data_or_134_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_54_nl;
  wire[30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_159_nl;
  wire act_regs_data_mux_137_nl;
  wire act_regs_data_or_135_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_47_nl;
  wire[30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_157_nl;
  wire act_regs_data_mux_138_nl;
  wire act_regs_data_or_136_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_40_nl;
  wire[30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_155_nl;
  wire act_regs_data_mux_139_nl;
  wire act_regs_data_or_137_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_33_nl;
  wire[30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_153_nl;
  wire act_regs_data_mux_140_nl;
  wire act_regs_data_or_138_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_26_nl;
  wire[30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_151_nl;
  wire act_regs_data_mux_141_nl;
  wire act_regs_data_or_139_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_19_nl;
  wire[30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_149_nl;
  wire act_regs_data_mux_142_nl;
  wire act_regs_data_or_140_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_111_nl;
  wire[30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_147_nl;
  wire act_regs_data_mux_143_nl;
  wire act_regs_data_or_141_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_5_nl;
  wire[30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_145_nl;
  wire act_regs_data_mux_144_nl;
  wire act_regs_data_or_142_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_67_nl;
  wire[30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_143_nl;
  wire act_regs_data_mux_145_nl;
  wire act_regs_data_or_143_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_102_nl;
  wire[30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_142_nl;
  wire act_regs_data_mux_146_nl;
  wire act_regs_data_or_144_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_95_nl;
  wire[30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_144_nl;
  wire act_regs_data_mux_147_nl;
  wire act_regs_data_or_145_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_88_nl;
  wire[30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_146_nl;
  wire act_regs_data_mux_148_nl;
  wire act_regs_data_or_146_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_81_nl;
  wire[30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_148_nl;
  wire act_regs_data_mux_149_nl;
  wire act_regs_data_or_147_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_74_nl;
  wire[30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_150_nl;
  wire act_regs_data_mux_150_nl;
  wire act_regs_data_or_148_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_10_nl;
  wire[30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_152_nl;
  wire act_regs_data_mux_151_nl;
  wire act_regs_data_or_149_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_60_nl;
  wire[30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_154_nl;
  wire act_regs_data_mux_152_nl;
  wire act_regs_data_or_150_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_52_nl;
  wire[30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_156_nl;
  wire act_regs_data_mux_153_nl;
  wire act_regs_data_or_151_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_45_nl;
  wire[30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_158_nl;
  wire act_regs_data_mux_154_nl;
  wire act_regs_data_or_152_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_38_nl;
  wire[30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_160_nl;
  wire act_regs_data_mux_155_nl;
  wire act_regs_data_or_153_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_31_nl;
  wire[30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_162_nl;
  wire act_regs_data_mux_156_nl;
  wire act_regs_data_or_154_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_24_nl;
  wire[30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_164_nl;
  wire act_regs_data_mux_157_nl;
  wire act_regs_data_or_155_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_17_nl;
  wire[30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_166_nl;
  wire act_regs_data_mux_158_nl;
  wire act_regs_data_or_156_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_109_nl;
  wire[30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_168_nl;
  wire act_regs_data_mux_159_nl;
  wire act_regs_data_or_157_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_3_nl;
  wire[30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_170_nl;
  wire act_regs_data_mux_160_nl;
  wire act_regs_data_or_158_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_66_nl;
  wire[30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_172_nl;
  wire act_regs_data_mux_161_nl;
  wire act_regs_data_or_159_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_59_nl;
  wire[30:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_175_nl;
  wire ActUnit_DecodeAxiWrite_mux_4_nl;
  wire act_config_ActConfigWrite_mux_1_nl;
  wire ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_23_nl;
  wire ActUnit_DecodeAxiRead_else_mux_3_nl;
  wire while_and_64_nl;
  wire[30:0] Silu_for_else_mux_1_nl;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_not_34_nl;
  wire[29:0] Silu_for_1_else_else_acc_nl;
  wire[30:0] nl_Silu_for_1_else_else_acc_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_10_nl;
  wire Silu_for_Silu_for_and_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_48_nl;
  wire mux_223_nl;
  wire mux_222_nl;
  wire[30:0] ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_83_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_and_36_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_and_37_nl;
  wire nor_772_nl;
  wire mux_224_nl;
  wire[30:0] Silu_for_else_mux_3_nl;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_not_36_nl;
  wire[30:0] Silu_for_else_mux_2_nl;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_not_35_nl;
  wire mux_226_nl;
  wire mux_225_nl;
  wire[30:0] Silu_for_else_mux_5_nl;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_not_38_nl;
  wire[30:0] Silu_for_else_mux_4_nl;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_not_37_nl;
  wire mux_227_nl;
  wire or_993_nl;
  wire or_994_nl;
  wire[30:0] Silu_for_else_mux_7_nl;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_not_40_nl;
  wire[30:0] Silu_for_else_mux_6_nl;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_not_39_nl;
  wire[30:0] Silu_for_else_mux_8_nl;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_not_41_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_15_nl;
  wire Gelu_for_Gelu_for_and_1_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_89_nl;
  wire[30:0] ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_78_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_and_38_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_and_39_nl;
  wire nor_773_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_20_nl;
  wire Silu_for_Silu_for_and_9_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_55_nl;
  wire[30:0] ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_82_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_and_40_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_and_41_nl;
  wire nor_774_nl;
  wire Gelu_for_Gelu_for_and_nl;
  wire[30:0] Gelu_for_Gelu_for_and_19_nl;
  wire[30:0] Gelu_for_else_mux_nl;
  wire operator_32_8_true_AC_TRN_AC_WRAP_3_not_34_nl;
  wire[30:0] Silu_for_else_mux_11_nl;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_not_42_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_25_nl;
  wire Gelu_for_Gelu_for_and_2_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_96_nl;
  wire[30:0] ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_77_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_and_42_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_and_43_nl;
  wire nor_775_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_30_nl;
  wire Silu_for_Silu_for_and_10_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_61_nl;
  wire[30:0] ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_81_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_and_44_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_and_45_nl;
  wire nor_776_nl;
  wire mux_232_nl;
  wire[30:0] Silu_for_else_mux_13_nl;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_not_44_nl;
  wire[30:0] Silu_for_else_mux_12_nl;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_not_43_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_35_nl;
  wire Gelu_for_Gelu_for_and_3_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_103_nl;
  wire[30:0] ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_76_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_and_46_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_and_47_nl;
  wire nor_777_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_40_nl;
  wire Gelu_for_Gelu_for_and_4_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_110_nl;
  wire[30:0] ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_88_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_and_48_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_and_49_nl;
  wire nor_778_nl;
  wire[30:0] Silu_for_else_mux_15_nl;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_not_46_nl;
  wire[30:0] Silu_for_else_mux_14_nl;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_not_45_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_45_nl;
  wire Gelu_for_Gelu_for_and_5_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_20_nl;
  wire[30:0] ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_87_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_and_50_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_and_51_nl;
  wire nor_779_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_50_nl;
  wire Gelu_for_Gelu_for_and_6_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_27_nl;
  wire[30:0] ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_86_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_and_52_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_and_53_nl;
  wire nor_780_nl;
  wire[28:0] Gelu_for_13_else_else_acc_nl;
  wire[29:0] nl_Gelu_for_13_else_else_acc_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_55_nl;
  wire Gelu_for_Gelu_for_and_12_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_13_nl;
  wire[30:0] ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_89_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_and_54_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_and_55_nl;
  wire nor_781_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_60_nl;
  wire Gelu_for_Gelu_for_and_13_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_75_nl;
  wire[30:0] ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_80_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_and_56_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_and_57_nl;
  wire nor_782_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_65_nl;
  wire Gelu_for_Gelu_for_and_14_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_82_nl;
  wire[30:0] ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_79_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_and_58_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_and_59_nl;
  wire nor_783_nl;
  wire[28:0] Gelu_for_8_else_else_acc_nl;
  wire[29:0] nl_Gelu_for_8_else_else_acc_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_70_nl;
  wire Gelu_for_Gelu_for_and_7_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_34_nl;
  wire[30:0] ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_85_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_and_60_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_and_61_nl;
  wire nor_784_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_75_nl;
  wire Gelu_for_Gelu_for_and_8_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_41_nl;
  wire[30:0] ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_84_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_and_62_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_and_63_nl;
  wire nor_785_nl;
  wire while_and_273_nl;
  wire while_while_mux1h_84_nl;
  wire and_1460_nl;
  wire mux_354_nl;
  wire while_and_272_nl;
  wire while_while_mux1h_85_nl;
  wire while_and_271_nl;
  wire while_while_mux1h_86_nl;
  wire while_and_270_nl;
  wire while_while_mux1h_87_nl;
  wire while_and_269_nl;
  wire while_while_mux1h_88_nl;
  wire while_and_268_nl;
  wire while_while_mux1h_89_nl;
  wire while_and_267_nl;
  wire while_while_mux1h_90_nl;
  wire while_and_266_nl;
  wire while_while_mux1h_91_nl;
  wire while_and_265_nl;
  wire while_while_mux1h_92_nl;
  wire while_and_264_nl;
  wire while_while_mux1h_93_nl;
  wire while_and_263_nl;
  wire while_while_mux1h_94_nl;
  wire while_and_262_nl;
  wire while_while_mux1h_95_nl;
  wire while_and_261_nl;
  wire while_while_mux1h_96_nl;
  wire while_and_260_nl;
  wire while_while_mux1h_97_nl;
  wire while_and_259_nl;
  wire while_while_mux1h_98_nl;
  wire while_and_258_nl;
  wire while_while_mux1h_99_nl;
  wire while_and_257_nl;
  wire while_while_mux1h_100_nl;
  wire and_1496_nl;
  wire mux_410_nl;
  wire while_and_256_nl;
  wire while_while_mux1h_101_nl;
  wire while_and_255_nl;
  wire while_while_mux1h_102_nl;
  wire while_and_254_nl;
  wire while_while_mux1h_103_nl;
  wire while_and_253_nl;
  wire while_while_mux1h_104_nl;
  wire while_and_252_nl;
  wire while_while_mux1h_105_nl;
  wire while_and_251_nl;
  wire while_while_mux1h_106_nl;
  wire while_and_250_nl;
  wire while_while_mux1h_107_nl;
  wire while_and_249_nl;
  wire while_while_mux1h_108_nl;
  wire while_and_248_nl;
  wire while_while_mux1h_109_nl;
  wire while_and_247_nl;
  wire while_while_mux1h_110_nl;
  wire while_and_246_nl;
  wire while_while_mux1h_111_nl;
  wire while_and_245_nl;
  wire while_while_mux1h_112_nl;
  wire while_and_244_nl;
  wire while_while_mux1h_113_nl;
  wire while_and_243_nl;
  wire while_while_mux1h_114_nl;
  wire while_and_242_nl;
  wire while_while_mux1h_115_nl;
  wire while_and_241_nl;
  wire while_while_mux1h_116_nl;
  wire and_1532_nl;
  wire mux_466_nl;
  wire while_and_240_nl;
  wire while_while_mux1h_117_nl;
  wire while_and_239_nl;
  wire while_while_mux1h_118_nl;
  wire while_and_238_nl;
  wire while_while_mux1h_119_nl;
  wire while_and_237_nl;
  wire while_while_mux1h_120_nl;
  wire while_and_236_nl;
  wire while_while_mux1h_121_nl;
  wire while_and_235_nl;
  wire while_while_mux1h_122_nl;
  wire while_and_234_nl;
  wire while_while_mux1h_123_nl;
  wire while_and_233_nl;
  wire while_while_mux1h_124_nl;
  wire while_and_232_nl;
  wire while_while_mux1h_125_nl;
  wire while_and_231_nl;
  wire while_while_mux1h_126_nl;
  wire while_and_230_nl;
  wire while_while_mux1h_127_nl;
  wire while_and_229_nl;
  wire while_while_mux1h_128_nl;
  wire while_and_228_nl;
  wire while_while_mux1h_129_nl;
  wire while_and_227_nl;
  wire while_while_mux1h_130_nl;
  wire while_and_226_nl;
  wire while_while_mux1h_131_nl;
  wire while_and_225_nl;
  wire while_while_mux1h_132_nl;
  wire and_1568_nl;
  wire mux_522_nl;
  wire while_and_224_nl;
  wire while_while_mux1h_133_nl;
  wire while_and_223_nl;
  wire while_while_mux1h_134_nl;
  wire while_and_222_nl;
  wire while_while_mux1h_135_nl;
  wire while_and_221_nl;
  wire while_while_mux1h_136_nl;
  wire while_and_220_nl;
  wire while_while_mux1h_137_nl;
  wire while_and_219_nl;
  wire while_while_mux1h_138_nl;
  wire while_and_218_nl;
  wire while_while_mux1h_139_nl;
  wire while_and_217_nl;
  wire while_while_mux1h_140_nl;
  wire while_and_216_nl;
  wire while_while_mux1h_141_nl;
  wire while_and_215_nl;
  wire while_while_mux1h_142_nl;
  wire while_and_214_nl;
  wire while_while_mux1h_143_nl;
  wire while_and_213_nl;
  wire while_while_mux1h_144_nl;
  wire while_and_212_nl;
  wire while_while_mux1h_145_nl;
  wire while_and_211_nl;
  wire while_while_mux1h_146_nl;
  wire while_and_nl;
  wire while_while_mux1h_147_nl;
  wire mux_82_nl;
  wire or_399_nl;
  wire act_config_InstIncr_mux_2_nl;
  wire act_config_InstIncr_if_act_config_InstIncr_if_and_nl;
  wire ActUnit_RunInst_switch_lp_nor_nl;
  wire[4:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_6_nl;
  wire[4:0] ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_and_18_nl;
  wire ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_nl;
  wire ActUnit_DecodeAxiWrite_else_not_17_nl;
  wire[31:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_7_nl;
  wire[31:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_8_nl;
  wire[31:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_9_nl;
  wire[31:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_10_nl;
  wire[31:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_11_nl;
  wire[31:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_12_nl;
  wire[31:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_13_nl;
  wire[31:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_14_nl;
  wire[31:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_15_nl;
  wire[31:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_16_nl;
  wire[31:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_17_nl;
  wire[31:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_18_nl;
  wire[31:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_19_nl;
  wire[31:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_20_nl;
  wire[31:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_21_nl;
  wire while_mux_32_nl;
  wire[30:0] while_mux_395_nl;
  wire while_while_nand_nl;
  wire[30:0] Gelu_for_else_mux_15_nl;
  wire operator_32_8_true_AC_TRN_AC_WRAP_3_not_31_nl;
  wire[30:0] Gelu_for_else_mux_10_nl;
  wire operator_32_8_true_AC_TRN_AC_WRAP_3_not_32_nl;
  wire[30:0] Gelu_for_else_mux_9_nl;
  wire operator_32_8_true_AC_TRN_AC_WRAP_3_not_33_nl;
  wire[30:0] Tanh_for_16_else_else_acc_nl;
  wire[31:0] nl_Tanh_for_16_else_else_acc_nl;
  wire Tanh_for_Tanh_for_nor_15_nl;
  wire Tanh_for_and_79_nl;
  wire[30:0] Tanh_for_15_else_else_acc_nl;
  wire[31:0] nl_Tanh_for_15_else_else_acc_nl;
  wire Tanh_for_Tanh_for_nor_14_nl;
  wire Tanh_for_and_77_nl;
  wire[30:0] Tanh_for_14_else_else_acc_nl;
  wire[31:0] nl_Tanh_for_14_else_else_acc_nl;
  wire Tanh_for_Tanh_for_nor_13_nl;
  wire Tanh_for_and_75_nl;
  wire[30:0] Tanh_for_13_else_else_acc_nl;
  wire[31:0] nl_Tanh_for_13_else_else_acc_nl;
  wire Tanh_for_Tanh_for_nor_12_nl;
  wire Tanh_for_and_73_nl;
  wire[30:0] Tanh_for_12_else_else_acc_nl;
  wire[31:0] nl_Tanh_for_12_else_else_acc_nl;
  wire Tanh_for_Tanh_for_nor_11_nl;
  wire Tanh_for_and_71_nl;
  wire[30:0] Tanh_for_11_else_else_acc_nl;
  wire[31:0] nl_Tanh_for_11_else_else_acc_nl;
  wire Tanh_for_Tanh_for_nor_10_nl;
  wire Tanh_for_and_69_nl;
  wire[30:0] Tanh_for_10_else_else_acc_nl;
  wire[31:0] nl_Tanh_for_10_else_else_acc_nl;
  wire Tanh_for_Tanh_for_nor_9_nl;
  wire Tanh_for_and_67_nl;
  wire[30:0] Tanh_for_9_else_else_acc_nl;
  wire[31:0] nl_Tanh_for_9_else_else_acc_nl;
  wire Tanh_for_Tanh_for_nor_8_nl;
  wire Tanh_for_and_65_nl;
  wire[30:0] Tanh_for_8_else_else_acc_nl;
  wire[31:0] nl_Tanh_for_8_else_else_acc_nl;
  wire Tanh_for_Tanh_for_nor_7_nl;
  wire Tanh_for_and_63_nl;
  wire[30:0] Tanh_for_7_else_else_acc_nl;
  wire[31:0] nl_Tanh_for_7_else_else_acc_nl;
  wire Tanh_for_Tanh_for_nor_6_nl;
  wire Tanh_for_and_61_nl;
  wire[30:0] Tanh_for_6_else_else_acc_nl;
  wire[31:0] nl_Tanh_for_6_else_else_acc_nl;
  wire Tanh_for_Tanh_for_nor_5_nl;
  wire Tanh_for_and_59_nl;
  wire[30:0] Tanh_for_5_else_else_acc_nl;
  wire[31:0] nl_Tanh_for_5_else_else_acc_nl;
  wire Tanh_for_Tanh_for_nor_4_nl;
  wire Tanh_for_and_57_nl;
  wire[30:0] Tanh_for_4_else_else_acc_nl;
  wire[31:0] nl_Tanh_for_4_else_else_acc_nl;
  wire Tanh_for_Tanh_for_nor_3_nl;
  wire Tanh_for_and_55_nl;
  wire[30:0] Tanh_for_3_else_else_acc_nl;
  wire[31:0] nl_Tanh_for_3_else_else_acc_nl;
  wire Tanh_for_Tanh_for_nor_2_nl;
  wire Tanh_for_and_53_nl;
  wire[30:0] Tanh_for_2_else_else_acc_nl;
  wire[31:0] nl_Tanh_for_2_else_else_acc_nl;
  wire Tanh_for_Tanh_for_nor_1_nl;
  wire Tanh_for_and_51_nl;
  wire[30:0] Tanh_for_1_else_else_acc_nl;
  wire[31:0] nl_Tanh_for_1_else_else_acc_nl;
  wire Tanh_for_Tanh_for_nor_nl;
  wire Tanh_for_and_49_nl;
  wire[4:0] ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_and_1_nl;
  wire nor_60_nl;
  wire or_170_nl;
  wire mux_54_nl;
  wire nor_63_nl;
  wire mux_48_nl;
  wire nand_nl;
  wire or_86_nl;
  wire nor_128_nl;
  wire nor_129_nl;
  wire nor_130_nl;
  wire nor_131_nl;
  wire mux_152_nl;
  wire and_710_nl;
  wire and_709_nl;
  wire mux_216_nl;
  wire mux_228_nl;
  wire mux_230_nl;
  wire mux_233_nl;
  wire mux_212_nl;
  wire nand_214_nl;
  wire or_605_nl;
  wire mux_578_nl;
  wire nor_768_nl;
  wire or_1509_nl;
  wire mux_94_nl;
  wire mux_93_nl;
  wire mux_92_nl;
  wire and_568_nl;
  wire mux_91_nl;
  wire mux_577_nl;
  wire mux_576_nl;
  wire and_1602_nl;
  wire mux_573_nl;
  wire mux_564_nl;
  wire or_1495_nl;
  wire mux_569_nl;
  wire mux_568_nl;
  wire and_1596_nl;
  wire mux_565_nl;
  wire mux_622_nl;
  wire or_1481_nl;
  wire mux_561_nl;
  wire nand_448_nl;
  wire mux_558_nl;
  wire or_1467_nl;
  wire mux_555_nl;
  wire or_1460_nl;
  wire mux_552_nl;
  wire or_1453_nl;
  wire mux_549_nl;
  wire mux_540_nl;
  wire or_1446_nl;
  wire mux_545_nl;
  wire mux_621_nl;
  wire or_1439_nl;
  wire mux_541_nl;
  wire mux_620_nl;
  wire or_1432_nl;
  wire mux_537_nl;
  wire mux_536_nl;
  wire or_1425_nl;
  wire mux_533_nl;
  wire or_1418_nl;
  wire mux_530_nl;
  wire or_1411_nl;
  wire mux_527_nl;
  wire or_1404_nl;
  wire mux_524_nl;
  wire or_1397_nl;
  wire mux_521_nl;
  wire mux_512_nl;
  wire or_1391_nl;
  wire mux_517_nl;
  wire mux_508_nl;
  wire or_1385_nl;
  wire mux_513_nl;
  wire mux_619_nl;
  wire or_1379_nl;
  wire mux_509_nl;
  wire mux_618_nl;
  wire or_1373_nl;
  wire mux_505_nl;
  wire or_1367_nl;
  wire mux_502_nl;
  wire or_1361_nl;
  wire mux_499_nl;
  wire or_1355_nl;
  wire mux_496_nl;
  wire or_1349_nl;
  wire mux_493_nl;
  wire mux_484_nl;
  wire or_1343_nl;
  wire mux_489_nl;
  wire mux_617_nl;
  wire or_1337_nl;
  wire mux_485_nl;
  wire mux_616_nl;
  wire or_1331_nl;
  wire mux_481_nl;
  wire mux_480_nl;
  wire or_1325_nl;
  wire mux_477_nl;
  wire or_1319_nl;
  wire mux_474_nl;
  wire or_1313_nl;
  wire mux_471_nl;
  wire or_1307_nl;
  wire mux_468_nl;
  wire or_1301_nl;
  wire mux_465_nl;
  wire mux_456_nl;
  wire or_1294_nl;
  wire mux_461_nl;
  wire mux_452_nl;
  wire or_1287_nl;
  wire mux_457_nl;
  wire mux_615_nl;
  wire or_1280_nl;
  wire mux_453_nl;
  wire mux_614_nl;
  wire or_1273_nl;
  wire mux_449_nl;
  wire or_1266_nl;
  wire mux_446_nl;
  wire or_1259_nl;
  wire mux_443_nl;
  wire or_1252_nl;
  wire mux_440_nl;
  wire or_1245_nl;
  wire mux_437_nl;
  wire mux_428_nl;
  wire or_1238_nl;
  wire mux_433_nl;
  wire mux_613_nl;
  wire or_1231_nl;
  wire mux_429_nl;
  wire mux_612_nl;
  wire or_1224_nl;
  wire mux_425_nl;
  wire mux_424_nl;
  wire or_1217_nl;
  wire mux_421_nl;
  wire or_1210_nl;
  wire mux_418_nl;
  wire or_1203_nl;
  wire mux_415_nl;
  wire or_1196_nl;
  wire mux_412_nl;
  wire or_1189_nl;
  wire mux_349_nl;
  wire or_1078_nl;
  wire mux_409_nl;
  wire mux_400_nl;
  wire or_1183_nl;
  wire mux_345_nl;
  wire and_1456_nl;
  wire mux_405_nl;
  wire mux_396_nl;
  wire or_1177_nl;
  wire mux_338_nl;
  wire and_1454_nl;
  wire mux_401_nl;
  wire mux_611_nl;
  wire or_1171_nl;
  wire mux_331_nl;
  wire nor_362_nl;
  wire mux_397_nl;
  wire mux_610_nl;
  wire or_1165_nl;
  wire mux_393_nl;
  wire or_1159_nl;
  wire mux_390_nl;
  wire or_1153_nl;
  wire mux_387_nl;
  wire or_1147_nl;
  wire mux_341_nl;
  wire or_1076_nl;
  wire mux_384_nl;
  wire or_1141_nl;
  wire mux_335_nl;
  wire or_1074_nl;
  wire mux_381_nl;
  wire mux_372_nl;
  wire or_1135_nl;
  wire mux_327_nl;
  wire mux_326_nl;
  wire mux_325_nl;
  wire and_1449_nl;
  wire mux_324_nl;
  wire and_1450_nl;
  wire mux_377_nl;
  wire mux_609_nl;
  wire or_1129_nl;
  wire mux_373_nl;
  wire mux_608_nl;
  wire or_1123_nl;
  wire mux_369_nl;
  wire mux_368_nl;
  wire or_1117_nl;
  wire mux_353_nl;
  wire nor_372_nl;
  wire mux_365_nl;
  wire or_1111_nl;
  wire mux_351_nl;
  wire or_1080_nl;
  wire mux_362_nl;
  wire or_1105_nl;
  wire mux_359_nl;
  wire or_1099_nl;
  wire mux_323_nl;
  wire mux_322_nl;
  wire mux_321_nl;
  wire or_1069_nl;
  wire mux_356_nl;
  wire or_1093_nl;
  wire mux_221_nl;
  wire or_991_nl;
  wire[28:0] Gelu_for_12_else_else_acc_rg_1_nl;
  wire[29:0] nl_Gelu_for_12_else_else_acc_rg_1_nl;
  wire[25:0] Gelu_for_else_else_mux1h_10_nl;
  wire and_1143_nl;
  wire and_1146_nl;
  wire and_1148_nl;
  wire[28:0] Gelu_for_10_else_else_acc_rg_1_nl;
  wire[29:0] nl_Gelu_for_10_else_else_acc_rg_1_nl;
  wire[25:0] Gelu_for_else_else_mux1h_12_nl;
  wire and_1162_nl;
  wire[28:0] Gelu_for_11_else_else_acc_rg_1_nl;
  wire[29:0] nl_Gelu_for_11_else_else_acc_rg_1_nl;
  wire[25:0] Gelu_for_else_else_mux1h_14_nl;
  wire and_1175_nl;
  wire[29:0] Silu_for_10_else_else_acc_rg_1_nl;
  wire[30:0] nl_Silu_for_10_else_else_acc_rg_1_nl;
  wire[26:0] Silu_for_else_else_mux1h_1_nl;
  wire and_1179_nl;
  wire[29:0] Silu_for_11_else_else_acc_rg_1_nl;
  wire[30:0] nl_Silu_for_11_else_else_acc_rg_1_nl;
  wire[26:0] Silu_for_else_else_mux1h_3_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [25:0] nl_Tanh_for_3_else_else_mul_1_cmp_b;
  assign nl_Tanh_for_3_else_else_mul_1_cmp_b = nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[25:0];
  wire [25:0] nl_Tanh_for_3_else_else_mul_1_cmp_1_b;
  assign nl_Tanh_for_3_else_else_mul_1_cmp_1_b = nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[25:0];
  wire [25:0] nl_Tanh_for_3_else_else_mul_1_cmp_2_b;
  assign nl_Tanh_for_3_else_else_mul_1_cmp_2_b = nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[25:0];
  wire [25:0] nl_Tanh_for_3_else_else_mul_1_cmp_3_b;
  assign nl_Tanh_for_3_else_else_mul_1_cmp_3_b = nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[25:0];
  wire [25:0] nl_Tanh_for_3_else_else_mul_1_cmp_4_b;
  assign nl_Tanh_for_3_else_else_mul_1_cmp_4_b = nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[25:0];
  wire [25:0] nl_Tanh_for_3_else_else_mul_1_cmp_5_b;
  assign nl_Tanh_for_3_else_else_mul_1_cmp_5_b = nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[25:0];
  wire [25:0] nl_Tanh_for_3_else_else_mul_1_cmp_6_b;
  assign nl_Tanh_for_3_else_else_mul_1_cmp_6_b = nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[25:0];
  wire [25:0] nl_Tanh_for_3_else_else_mul_1_cmp_7_b;
  assign nl_Tanh_for_3_else_else_mul_1_cmp_7_b = nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[25:0];
  wire [25:0] nl_Tanh_for_3_else_else_mul_1_cmp_8_b;
  assign nl_Tanh_for_3_else_else_mul_1_cmp_8_b = nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[25:0];
  wire [25:0] nl_Tanh_for_3_else_else_mul_1_cmp_9_b;
  assign nl_Tanh_for_3_else_else_mul_1_cmp_9_b = nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[25:0];
  wire [25:0] nl_Tanh_for_3_else_else_mul_1_cmp_10_b;
  assign nl_Tanh_for_3_else_else_mul_1_cmp_10_b = nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[25:0];
  wire [25:0] nl_Tanh_for_3_else_else_mul_1_cmp_11_b;
  assign nl_Tanh_for_3_else_else_mul_1_cmp_11_b = nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[25:0];
  wire [25:0] nl_Tanh_for_3_else_else_mul_1_cmp_12_b;
  assign nl_Tanh_for_3_else_else_mul_1_cmp_12_b = nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[25:0];
  wire [25:0] nl_Tanh_for_3_else_else_mul_1_cmp_13_b;
  assign nl_Tanh_for_3_else_else_mul_1_cmp_13_b = nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[25:0];
  wire [25:0] nl_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_1_a;
  assign nl_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_1_a = nv_scvector_cctor_nv_scvector_6_for_16_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0];
  wire [25:0] nl_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_6_a;
  assign nl_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_6_a = nv_scvector_cctor_nv_scvector_6_for_11_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0];
  wire [25:0] nl_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_7_a;
  assign nl_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_7_a = nv_scvector_cctor_nv_scvector_6_for_10_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0];
  wire [25:0] nl_Tanh_for_1_else_else_mul_cmp_a;
  assign nl_Tanh_for_1_else_else_mul_cmp_a = MUX1HOT_v_26_7_2((nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[25:0]),
      reg_ActUnit_RunInst_case_11_nv_scvector_cctor_data_0_ftd_6, (ActUnit_RunInst_case_15_nv_scvector_cctor_data_0_sva_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_6_for_5_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_6_for_7_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_6_for_14_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_6_for_11_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      {and_dcpl_554 , and_dcpl_604 , and_dcpl_612 , and_dcpl_614 , and_dcpl_600 ,
      and_dcpl_576 , and_dcpl_578});
  wire[1:0] Tanh_for_else_else_and_nl;
  wire[1:0] Tanh_for_else_else_mux1h_31_nl;
  wire not_1260_nl;
  wire Tanh_for_else_else_and_1_nl;
  wire Tanh_for_else_else_mux1h_59_nl;
  wire[45:0] Tanh_for_else_else_mux1h_60_nl;
  wire [48:0] nl_Tanh_for_1_else_else_mul_cmp_b;
  assign Tanh_for_else_else_mux1h_31_nl = MUX1HOT_v_2_4_2((Tanh_for_1_else_else_mul_1_cmp_z[48:47]),
      (signext_2_1(Tanh_for_1_else_else_mul_1_cmp_z[46])), (signext_2_1(Tanh_for_1_else_else_mul_1_cmp_1_z[46])),
      (signext_2_1(Gelu_for_else_else_slc_Tanh_for_1_else_else_mul_cmp_z_46_0_itm[46])),
      {and_dcpl_604 , and_dcpl_612 , and_dcpl_609 , and_dcpl_576});
  assign not_1260_nl = ~ and_dcpl_554;
  assign Tanh_for_else_else_and_nl = MUX_v_2_2_2(2'b00, Tanh_for_else_else_mux1h_31_nl,
      not_1260_nl);
  assign Tanh_for_else_else_mux1h_59_nl = MUX1HOT_s_1_3_2((Tanh_for_1_else_else_mul_1_cmp_z[46]),
      (Tanh_for_1_else_else_mul_1_cmp_1_z[46]), (Gelu_for_else_else_slc_Tanh_for_1_else_else_mul_cmp_z_46_0_itm[46]),
      {Tanh_for_else_else_or_1_cse , and_dcpl_609 , and_dcpl_576});
  assign Tanh_for_else_else_and_1_nl = Tanh_for_else_else_mux1h_59_nl & (~ and_dcpl_554);
  assign Tanh_for_else_else_mux1h_60_nl = MUX1HOT_v_46_4_2(46'b0000000000000000000000000110011000100001000101,
      (Tanh_for_1_else_else_mul_1_cmp_z[45:0]), (Tanh_for_1_else_else_mul_1_cmp_1_z[45:0]),
      (Gelu_for_else_else_slc_Tanh_for_1_else_else_mul_cmp_z_46_0_itm[45:0]), {and_dcpl_554
      , Tanh_for_else_else_or_1_cse , and_dcpl_609 , and_dcpl_576});
  assign nl_Tanh_for_1_else_else_mul_cmp_b = {Tanh_for_else_else_and_nl , Tanh_for_else_else_and_1_nl
      , Tanh_for_else_else_mux1h_60_nl};
  wire [25:0] nl_Tanh_for_1_else_else_mul_cmp_1_a;
  assign nl_Tanh_for_1_else_else_mul_cmp_1_a = nv_scvector_cctor_nv_scvector_6_for_16_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0];
  wire [25:0] nl_Tanh_for_1_else_else_mul_cmp_6_a;
  assign nl_Tanh_for_1_else_else_mul_cmp_6_a = nv_scvector_cctor_nv_scvector_6_for_11_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0];
  wire [25:0] nl_Tanh_for_1_else_else_mul_cmp_7_a;
  assign nl_Tanh_for_1_else_else_mul_cmp_7_a = nv_scvector_cctor_nv_scvector_6_for_10_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0];
  wire [25:0] nl_Tanh_for_1_else_else_mul_cmp_12_a;
  assign nl_Tanh_for_1_else_else_mul_cmp_12_a = MUX1HOT_v_26_8_2((nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[25:0]),
      reg_nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6,
      (nv_scvector_cctor_nv_scvector_6_for_2_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_6_for_3_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_6_for_4_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_6_for_6_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_6_for_15_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_6_for_10_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      {and_dcpl_554 , and_dcpl_604 , and_dcpl_612 , and_dcpl_613 , and_dcpl_614 ,
      and_dcpl_600 , and_dcpl_576 , and_dcpl_578});
  wire and_640_nl;
  wire [48:0] nl_Tanh_for_1_else_else_mul_cmp_12_b;
  assign and_640_nl = (~((~((act_config_in_InstFetch_return_sva_7_2[4]) | (fsm_output[0])))
      | (fsm_output[3]))) & (fsm_output[2]) & (~ (fsm_output[1])) & (~ (fsm_output[4]));
  assign nl_Tanh_for_1_else_else_mul_cmp_12_b = MUX1HOT_v_49_5_2(49'b0000000000000000000000000000110011000100001000101,
      Tanh_for_3_else_else_mul_1_cmp_12_z, (signext_49_47(Tanh_for_1_else_else_mul_1_cmp_1_z[46:0])),
      (signext_49_47(Tanh_for_1_else_else_mul_1_cmp_z[46:0])), ({{2{Gelu_for_else_else_slc_Tanh_for_1_else_else_mul_cmp_12_z_46_0_itm[46]}},
      Gelu_for_else_else_slc_Tanh_for_1_else_else_mul_cmp_12_z_46_0_itm}), {and_dcpl_554
      , and_dcpl_604 , and_640_nl , and_dcpl_609 , and_dcpl_576});
  wire [25:0] nl_Tanh_for_1_else_else_mul_cmp_13_a;
  assign nl_Tanh_for_1_else_else_mul_cmp_13_a = MUX1HOT_v_26_5_2((nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[25:0]),
      reg_nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6,
      (nv_scvector_cctor_nv_scvector_6_for_12_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_6_for_9_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_6_for_16_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      {and_dcpl_554 , and_dcpl_592 , and_dcpl_600 , and_dcpl_576 , and_dcpl_578});
  wire [48:0] nl_Tanh_for_1_else_else_mul_cmp_13_b;
  assign nl_Tanh_for_1_else_else_mul_cmp_13_b = MUX1HOT_v_49_5_2(49'b0000000000000000000000000000110011000100001000101,
      Tanh_for_3_else_else_mul_1_cmp_13_z, ({{2{Gelu_for_else_else_slc_Tanh_for_1_else_else_mul_1_cmp_z_46_0_itm[46]}},
      Gelu_for_else_else_slc_Tanh_for_1_else_else_mul_1_cmp_z_46_0_itm}), (signext_49_47(Tanh_for_1_else_else_mul_1_cmp_1_z[46:0])),
      ({{2{Gelu_for_else_else_slc_Tanh_for_1_else_else_mul_cmp_13_z_46_0_itm[46]}},
      Gelu_for_else_else_slc_Tanh_for_1_else_else_mul_cmp_13_z_46_0_itm}), {and_dcpl_554
      , and_dcpl_592 , and_dcpl_600 , and_dcpl_576 , and_dcpl_578});
  wire [25:0] nl_Tanh_for_1_else_else_mul_cmp_14_a;
  assign nl_Tanh_for_1_else_else_mul_cmp_14_a = MUX_v_26_2_2(reg_nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6,
      (nv_scvector_cctor_nv_scvector_6_for_8_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      and_dcpl_576);
  wire [48:0] nl_Tanh_for_1_else_else_mul_cmp_14_b;
  assign nl_Tanh_for_1_else_else_mul_cmp_14_b = MUX_v_49_2_2(Tanh_for_3_else_else_mul_1_cmp_z,
      (signext_49_47(Tanh_for_1_else_else_mul_1_cmp_z[46:0])), and_dcpl_576);
  wire [25:0] nl_Tanh_for_1_else_else_mul_cmp_15_a;
  assign nl_Tanh_for_1_else_else_mul_cmp_15_a = MUX1HOT_v_26_3_2((nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[25:0]),
      reg_nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6,
      (nv_scvector_cctor_nv_scvector_6_for_13_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      {and_dcpl_554 , and_dcpl_592 , and_dcpl_576});
  wire [48:0] nl_Tanh_for_1_else_else_mul_cmp_15_b;
  assign nl_Tanh_for_1_else_else_mul_cmp_15_b = MUX1HOT_v_49_3_2(49'b0000000000000000000000000000110011000100001000101,
      (Tanh_for_1_else_else_mul_1_cmp_1_z[48:0]), ({{2{Gelu_for_else_else_slc_Tanh_for_1_else_else_mul_cmp_15_z_46_0_itm[46]}},
      Gelu_for_else_else_slc_Tanh_for_1_else_else_mul_cmp_15_z_46_0_itm}), {and_dcpl_554
      , and_dcpl_592 , and_dcpl_576});
  wire Tanh_for_else_else_mux1h_13_nl;
  wire[25:0] Tanh_for_else_else_mux1h_61_nl;
  wire [26:0] nl_Tanh_for_1_else_else_mul_1_cmp_a;
  assign Tanh_for_else_else_mux1h_13_nl = MUX1HOT_s_1_14_2((ActUnit_RunInst_case_11_nv_scvector_cctor_data_0_sva_1_30_0[26]),
      (ActUnit_RunInst_case_11_nv_scvector_cctor_data_0_sva_1_30_0[25]), (nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[26]),
      (nv_scvector_cctor_nv_scvector_6_for_12_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25]),
      (nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[26]),
      (nv_scvector_cctor_nv_scvector_6_for_4_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25]),
      (nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[26]),
      (nv_scvector_cctor_nv_scvector_6_for_6_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25]),
      (nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[26]),
      (nv_scvector_cctor_nv_scvector_6_for_8_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25]),
      (nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[26]),
      (nv_scvector_cctor_nv_scvector_6_for_10_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25]),
      (nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[26]),
      (nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[26]),
      {Tanh_for_else_else_and_8_cse , Tanh_for_else_else_and_9_cse , and_dcpl_562
      , and_dcpl_581 , and_dcpl_566 , and_dcpl_583 , and_dcpl_569 , and_dcpl_584
      , and_dcpl_572 , and_dcpl_585 , and_dcpl_573 , and_dcpl_586 , and_dcpl_576
      , and_dcpl_578});
  assign Tanh_for_else_else_mux1h_61_nl = MUX1HOT_v_26_13_2((ActUnit_RunInst_case_11_nv_scvector_cctor_data_0_sva_1_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_6_for_12_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_6_for_4_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_6_for_6_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_6_for_8_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_6_for_10_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      {and_dcpl_554 , and_dcpl_562 , and_dcpl_581 , and_dcpl_566 , and_dcpl_583 ,
      and_dcpl_569 , and_dcpl_584 , and_dcpl_572 , and_dcpl_585 , and_dcpl_573 ,
      and_dcpl_586 , and_dcpl_576 , and_dcpl_578});
  assign nl_Tanh_for_1_else_else_mul_1_cmp_a = {Tanh_for_else_else_mux1h_13_nl ,
      Tanh_for_else_else_mux1h_61_nl};
  wire [26:0] nl_Tanh_for_1_else_else_mul_1_cmp_b;
  assign nl_Tanh_for_1_else_else_mul_1_cmp_b = MUX1HOT_v_27_10_2(27'b111110101010101010101010101,
      (ActUnit_RunInst_case_11_nv_scvector_cctor_data_0_sva_1_30_0[26:0]), 27'b000000110011000100001000101,
      (nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[26:0]),
      (nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[26:0]),
      (nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[26:0]),
      (nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[26:0]),
      (nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[26:0]),
      (nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[26:0]),
      (nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[26:0]),
      {Tanh_for_else_else_and_2_cse , Tanh_for_else_else_and_3_cse , Tanh_for_else_else_or_cse
      , and_dcpl_562 , and_dcpl_566 , and_dcpl_569 , and_dcpl_572 , and_dcpl_573
      , and_dcpl_576 , and_dcpl_578});
  wire Tanh_for_else_else_mux1h_6_nl;
  wire[25:0] Tanh_for_else_else_mux1h_62_nl;
  wire [26:0] nl_Tanh_for_1_else_else_mul_1_cmp_1_a;
  assign Tanh_for_else_else_mux1h_6_nl = MUX1HOT_s_1_14_2((nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[26]),
      (nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[25]),
      (nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[26]),
      (nv_scvector_cctor_nv_scvector_6_for_3_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25]),
      (nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[26]),
      (nv_scvector_cctor_nv_scvector_6_for_5_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25]),
      (nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[26]),
      (nv_scvector_cctor_nv_scvector_6_for_7_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25]),
      (nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[26]),
      (nv_scvector_cctor_nv_scvector_6_for_9_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25]),
      (nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[26]),
      (nv_scvector_cctor_nv_scvector_6_for_11_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25]),
      (nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[26]),
      (nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[26]),
      {Tanh_for_else_else_and_8_cse , Tanh_for_else_else_and_9_cse , and_dcpl_562
      , and_dcpl_581 , and_dcpl_566 , and_dcpl_583 , and_dcpl_569 , and_dcpl_584
      , and_dcpl_572 , and_dcpl_585 , and_dcpl_573 , and_dcpl_586 , and_dcpl_576
      , and_dcpl_578});
  assign Tanh_for_else_else_mux1h_62_nl = MUX1HOT_v_26_13_2((nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_6_for_3_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_6_for_5_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_6_for_7_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_6_for_9_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_6_for_11_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      {and_dcpl_554 , and_dcpl_562 , and_dcpl_581 , and_dcpl_566 , and_dcpl_583 ,
      and_dcpl_569 , and_dcpl_584 , and_dcpl_572 , and_dcpl_585 , and_dcpl_573 ,
      and_dcpl_586 , and_dcpl_576 , and_dcpl_578});
  assign nl_Tanh_for_1_else_else_mul_1_cmp_1_a = {Tanh_for_else_else_mux1h_6_nl ,
      Tanh_for_else_else_mux1h_62_nl};
  wire [26:0] nl_Tanh_for_1_else_else_mul_1_cmp_1_b;
  assign nl_Tanh_for_1_else_else_mul_1_cmp_1_b = MUX1HOT_v_27_10_2(27'b111110101010101010101010101,
      (nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[26:0]),
      27'b000000110011000100001000101, (nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[26:0]),
      (nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[26:0]),
      (nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[26:0]),
      (nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[26:0]),
      (nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[26:0]),
      (nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[26:0]),
      (nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[26:0]),
      {Tanh_for_else_else_and_2_cse , Tanh_for_else_else_and_3_cse , Tanh_for_else_else_or_cse
      , and_dcpl_562 , and_dcpl_566 , and_dcpl_569 , and_dcpl_572 , and_dcpl_573
      , and_dcpl_576 , and_dcpl_578});
  wire  nl_ActUnit_ActUnitRun_rva_out_Push_mioi_inst_ActUnitRun_wten;
  assign nl_ActUnit_ActUnitRun_rva_out_Push_mioi_inst_ActUnitRun_wten = ~ ActUnitRun_wen;
  wire[31:0] ActUnit_PushAxiRsp_if_mux_11_nl;
  wire[31:0] ActUnit_PushAxiRsp_if_mux_10_nl;
  wire[31:0] ActUnit_PushAxiRsp_if_mux_9_nl;
  wire[31:0] ActUnit_PushAxiRsp_if_mux_8_nl;
  wire[31:0] ActUnit_PushAxiRsp_if_mux_7_nl;
  wire[31:0] ActUnit_PushAxiRsp_if_mux_6_nl;
  wire[31:0] ActUnit_PushAxiRsp_if_mux_5_nl;
  wire[31:0] ActUnit_PushAxiRsp_if_mux_4_nl;
  wire[31:0] ActUnit_PushAxiRsp_if_mux_3_nl;
  wire[31:0] ActUnit_PushAxiRsp_if_mux_2_nl;
  wire[31:0] ActUnit_PushAxiRsp_if_mux_1_nl;
  wire[31:0] ActUnit_PushAxiRsp_if_mux_nl;
  wire[7:0] act_mem_banks_read_read_data_mux_19_nl;
  wire[7:0] act_mem_banks_read_read_data_mux_18_nl;
  wire[7:0] act_mem_banks_read_read_data_mux_17_nl;
  wire[7:0] act_mem_banks_read_read_data_mux_16_nl;
  wire[7:0] act_mem_banks_read_read_data_mux_15_nl;
  wire[7:0] act_mem_banks_read_read_data_mux_14_nl;
  wire[7:0] act_mem_banks_read_read_data_mux_13_nl;
  wire[7:0] act_mem_banks_read_read_data_mux_12_nl;
  wire[7:0] act_mem_banks_read_read_data_mux_11_nl;
  wire[2:0] act_mem_banks_read_read_data_mux_10_nl;
  wire[4:0] act_mem_banks_read_read_data_mux_9_nl;
  wire[7:0] act_mem_banks_read_read_data_mux_8_nl;
  wire[7:0] act_mem_banks_read_read_data_mux_7_nl;
  wire[1:0] act_mem_banks_read_read_data_mux_6_nl;
  wire[5:0] act_mem_banks_read_read_data_mux_5_nl;
  wire[7:0] act_mem_banks_read_read_data_mux_4_nl;
  wire[6:0] act_mem_banks_read_read_data_mux_3_nl;
  wire act_mem_banks_read_read_data_mux_2_nl;
  wire[6:0] act_mem_banks_read_read_data_mux_1_nl;
  wire act_mem_banks_read_read_data_mux_nl;
  wire [511:0] nl_ActUnit_ActUnitRun_rva_out_Push_mioi_inst_rva_out_Push_mioi_m_data_rsc_dat_ActUnitRun;
  assign ActUnit_PushAxiRsp_if_mux_11_nl = MUX_v_32_2_2(rva_out_reg_data_511_480_sva_dfm_3,
      act_mem_banks_read_read_data_lpi_1_dfm_1_511_480_mx1, act_read_req_valid_lpi_1_dfm_6);
  assign ActUnit_PushAxiRsp_if_mux_10_nl = MUX_v_32_2_2(rva_out_reg_data_479_448_sva_dfm_3,
      act_mem_banks_read_read_data_lpi_1_dfm_1_479_448_mx1, act_read_req_valid_lpi_1_dfm_6);
  assign ActUnit_PushAxiRsp_if_mux_9_nl = MUX_v_32_2_2(rva_out_reg_data_447_416_sva_dfm_3,
      act_mem_banks_read_read_data_lpi_1_dfm_1_447_416_mx1, act_read_req_valid_lpi_1_dfm_6);
  assign ActUnit_PushAxiRsp_if_mux_8_nl = MUX_v_32_2_2(rva_out_reg_data_415_384_sva_dfm_3,
      act_mem_banks_read_read_data_lpi_1_dfm_1_415_384_mx1, act_read_req_valid_lpi_1_dfm_6);
  assign ActUnit_PushAxiRsp_if_mux_7_nl = MUX_v_32_2_2(rva_out_reg_data_383_352_sva_dfm_3,
      act_mem_banks_read_read_data_lpi_1_dfm_1_383_352_mx1, act_read_req_valid_lpi_1_dfm_6);
  assign ActUnit_PushAxiRsp_if_mux_6_nl = MUX_v_32_2_2(rva_out_reg_data_351_320_sva_dfm_3,
      act_mem_banks_read_read_data_lpi_1_dfm_1_351_320_mx1, act_read_req_valid_lpi_1_dfm_6);
  assign ActUnit_PushAxiRsp_if_mux_5_nl = MUX_v_32_2_2(rva_out_reg_data_319_288_sva_dfm_3,
      act_mem_banks_read_read_data_lpi_1_dfm_1_319_288_mx1, act_read_req_valid_lpi_1_dfm_6);
  assign ActUnit_PushAxiRsp_if_mux_4_nl = MUX_v_32_2_2(rva_out_reg_data_287_256_sva_dfm_3,
      act_mem_banks_read_read_data_lpi_1_dfm_1_287_256_mx1, act_read_req_valid_lpi_1_dfm_6);
  assign ActUnit_PushAxiRsp_if_mux_3_nl = MUX_v_32_2_2(rva_out_reg_data_255_224_sva_dfm_3,
      act_mem_banks_read_read_data_lpi_1_dfm_1_255_224_mx1, act_read_req_valid_lpi_1_dfm_6);
  assign ActUnit_PushAxiRsp_if_mux_2_nl = MUX_v_32_2_2(rva_out_reg_data_223_192_sva_dfm_3,
      act_mem_banks_read_read_data_lpi_1_dfm_1_223_192_mx1, act_read_req_valid_lpi_1_dfm_6);
  assign ActUnit_PushAxiRsp_if_mux_1_nl = MUX_v_32_2_2(rva_out_reg_data_191_160_sva_dfm_3,
      act_mem_banks_read_read_data_lpi_1_dfm_1_191_160_mx1, act_read_req_valid_lpi_1_dfm_6);
  assign ActUnit_PushAxiRsp_if_mux_nl = MUX_v_32_2_2(rva_out_reg_data_159_128_sva_dfm_3,
      act_mem_banks_read_read_data_lpi_1_dfm_1_159_128_mx1, act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_19_nl = MUX_v_8_2_2(rva_out_reg_data_127_120_sva_dfm_3,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_127_96_mx1[31:24]), act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_18_nl = MUX_v_8_2_2(rva_out_reg_data_119_112_sva_dfm_3,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_127_96_mx1[23:16]), act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_17_nl = MUX_v_8_2_2(rva_out_reg_data_111_104_sva_dfm_3,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_127_96_mx1[15:8]), act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_16_nl = MUX_v_8_2_2(rva_out_reg_data_103_96_sva_dfm_3,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_127_96_mx1[7:0]), act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_15_nl = MUX_v_8_2_2(rva_out_reg_data_95_88_sva_dfm_3,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_95_64_mx1[31:24]), act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_14_nl = MUX_v_8_2_2(rva_out_reg_data_87_80_sva_dfm_3,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_95_64_mx1[23:16]), act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_13_nl = MUX_v_8_2_2(rva_out_reg_data_79_72_sva_dfm_3,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_95_64_mx1[15:8]), act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_12_nl = MUX_v_8_2_2(rva_out_reg_data_71_64_sva_dfm_3,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_95_64_mx1[7:0]), act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_11_nl = MUX_v_8_2_2(rva_out_reg_data_63_56_sva_dfm_3,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_63_32_mx1[31:24]), act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_10_nl = MUX_v_3_2_2(rva_out_reg_data_55_53_sva_dfm_3,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_63_32_mx1[23:21]), act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_9_nl = MUX_v_5_2_2(rva_out_reg_data_52_48_sva_dfm_3,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_63_32_mx1[20:16]), act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_8_nl = MUX_v_8_2_2(rva_out_reg_data_47_40_sva_dfm_3,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_63_32_mx1[15:8]), act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_7_nl = MUX_v_8_2_2(rva_out_reg_data_39_32_sva_dfm_3,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_63_32_mx1[7:0]), act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_6_nl = MUX_v_2_2_2(rva_out_reg_data_31_30_sva_dfm_3,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_31_0_mx1[31:30]), act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_5_nl = MUX_v_6_2_2(rva_out_reg_data_29_24_sva_dfm_3,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_31_0_mx1[29:24]), act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_4_nl = MUX_v_8_2_2(rva_out_reg_data_23_16_sva_dfm_3,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_31_0_mx1[23:16]), act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_3_nl = MUX_v_7_2_2(rva_out_reg_data_15_9_sva_dfm_3,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_31_0_mx1[15:9]), act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_2_nl = MUX_s_1_2_2(rva_out_reg_data_8_sva_dfm_3,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_31_0_mx1[8]), act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_1_nl = MUX_v_7_2_2(rva_out_reg_data_7_1_sva_dfm_3,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_31_0_mx1[7:1]), act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_nl = MUX_s_1_2_2(rva_out_reg_data_0_sva_dfm_3,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_31_0_mx1[0]), act_read_req_valid_lpi_1_dfm_6);
  assign nl_ActUnit_ActUnitRun_rva_out_Push_mioi_inst_rva_out_Push_mioi_m_data_rsc_dat_ActUnitRun
      = {ActUnit_PushAxiRsp_if_mux_11_nl , ActUnit_PushAxiRsp_if_mux_10_nl , ActUnit_PushAxiRsp_if_mux_9_nl
      , ActUnit_PushAxiRsp_if_mux_8_nl , ActUnit_PushAxiRsp_if_mux_7_nl , ActUnit_PushAxiRsp_if_mux_6_nl
      , ActUnit_PushAxiRsp_if_mux_5_nl , ActUnit_PushAxiRsp_if_mux_4_nl , ActUnit_PushAxiRsp_if_mux_3_nl
      , ActUnit_PushAxiRsp_if_mux_2_nl , ActUnit_PushAxiRsp_if_mux_1_nl , ActUnit_PushAxiRsp_if_mux_nl
      , act_mem_banks_read_read_data_mux_19_nl , act_mem_banks_read_read_data_mux_18_nl
      , act_mem_banks_read_read_data_mux_17_nl , act_mem_banks_read_read_data_mux_16_nl
      , act_mem_banks_read_read_data_mux_15_nl , act_mem_banks_read_read_data_mux_14_nl
      , act_mem_banks_read_read_data_mux_13_nl , act_mem_banks_read_read_data_mux_12_nl
      , act_mem_banks_read_read_data_mux_11_nl , act_mem_banks_read_read_data_mux_10_nl
      , act_mem_banks_read_read_data_mux_9_nl , act_mem_banks_read_read_data_mux_8_nl
      , act_mem_banks_read_read_data_mux_7_nl , act_mem_banks_read_read_data_mux_6_nl
      , act_mem_banks_read_read_data_mux_5_nl , act_mem_banks_read_read_data_mux_4_nl
      , act_mem_banks_read_read_data_mux_3_nl , act_mem_banks_read_read_data_mux_2_nl
      , act_mem_banks_read_read_data_mux_1_nl , act_mem_banks_read_read_data_mux_nl};
  wire  nl_ActUnit_ActUnitRun_output_port_Push_mioi_inst_ActUnitRun_wten;
  assign nl_ActUnit_ActUnitRun_output_port_Push_mioi_inst_ActUnitRun_wten = ~ ActUnitRun_wen;
  wire ActUnit_PushOutput_if_for_ActUnit_PushOutput_if_for_and_nl;
  wire[30:0] ActUnit_PushOutput_if_for_ActUnit_PushOutput_if_for_and_1_nl;
  wire [511:0] nl_ActUnit_ActUnitRun_output_port_Push_mioi_inst_output_port_Push_mioi_m_data_data_rsc_dat_ActUnitRun;
  assign ActUnit_PushOutput_if_for_ActUnit_PushOutput_if_for_and_nl = ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_31
      & ActUnit_PushOutput_if_for_and_27_itm;
  assign ActUnit_PushOutput_if_for_ActUnit_PushOutput_if_for_and_1_nl = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_30_0, ActUnit_PushOutput_if_for_and_27_itm);
  assign nl_ActUnit_ActUnitRun_output_port_Push_mioi_inst_output_port_Push_mioi_m_data_data_rsc_dat_ActUnitRun
      = {ActUnit_PushOutput_if_for_ActUnit_PushOutput_if_for_and_nl , ActUnit_PushOutput_if_for_ActUnit_PushOutput_if_for_and_1_nl
      , ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_31 , ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_30_0
      , ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_31 , ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_30_0
      , ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_31 , ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_30_0
      , ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_31 , ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_30_0
      , ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_31 , ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_30_0
      , ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_31 , ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_30_0
      , ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_31 , ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_30_0
      , ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_31 , ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_30_0
      , ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_31 , ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_30_0
      , ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_31 , ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_30_0
      , ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_31 , ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_30_0
      , ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_31 , ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_30_0
      , ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_31 , ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_30_0
      , ActUnit_PushOutput_if_output_port_reg_data_data_1_sva_31 , ActUnit_PushOutput_if_output_port_reg_data_data_1_sva_30_0
      , ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_31 , ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_30_0};
  wire [8:0] nl_ActUnit_ActUnitRun_output_port_Push_mioi_inst_output_port_Push_mioi_m_logical_addr_rsc_dat_ActUnitRun;
  assign nl_ActUnit_ActUnitRun_output_port_Push_mioi_inst_output_port_Push_mioi_m_logical_addr_rsc_dat_ActUnitRun
      = act_config_output_counter_sva_dfm_3 + act_config_output_addr_base_sva;
  wire  nl_ActUnit_ActUnitRun_done_Push_mioi_inst_ActUnitRun_wten;
  assign nl_ActUnit_ActUnitRun_done_Push_mioi_inst_ActUnitRun_wten = ~ ActUnitRun_wen;
  wire  nl_ActUnit_ActUnitRun_ActUnitRun_fsm_inst_while_C_0_tr0;
  assign nl_ActUnit_ActUnitRun_ActUnitRun_fsm_inst_while_C_0_tr0 = (~(is_start_sva
      & (act_config_in_InstFetch_mux_tmp[5]))) | (act_config_in_InstFetch_mux_tmp[7])
      | (act_config_in_InstFetch_mux_tmp[6]) | (act_config_in_InstFetch_mux_tmp[4]);
  wire  nl_ActUnit_ActUnitRun_ActUnitRun_fsm_inst_ActUnit_RunInst_case_2_for_C_0_tr0;
  assign nl_ActUnit_ActUnitRun_ActUnitRun_fsm_inst_ActUnit_RunInst_case_2_for_C_0_tr0
      = ActUnit_RunInst_case_2_for_i_4_0_sva_2[4];
  wire  nl_ActUnit_ActUnitRun_ActUnitRun_fsm_inst_while_C_11_tr0;
  assign nl_ActUnit_ActUnitRun_ActUnitRun_fsm_inst_while_C_11_tr0 = ~(is_start_sva
      & ActUnit_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva);
  wire  nl_ActUnit_ActUnitRun_ActUnitRun_fsm_inst_ActUnit_PushOutput_if_for_C_0_tr0;
  assign nl_ActUnit_ActUnitRun_ActUnitRun_fsm_inst_ActUnit_PushOutput_if_for_C_0_tr0
      = ActUnit_RunInst_case_2_for_i_4_0_sva_2[4];
  wire  nl_ActUnit_ActUnitRun_ActUnitRun_fsm_inst_while_C_13_tr0;
  assign nl_ActUnit_ActUnitRun_ActUnitRun_fsm_inst_while_C_13_tr0 = (~ w_load_lpi_1_dfm_1)
      | act_config_is_zero_first_sva | (~ is_start_sva);
  wire  nl_ActUnit_ActUnitRun_ActUnitRun_fsm_inst_ActUnit_RunLoad_if_else_for_C_0_tr0;
  assign nl_ActUnit_ActUnitRun_ActUnitRun_fsm_inst_ActUnit_RunLoad_if_else_for_C_0_tr0
      = ActUnit_RunInst_case_2_for_i_4_0_sva_2[4];
  ActUnit_mgc_mul_pipe #(.width_a(32'sd23),
  .signd_a(32'sd1),
  .width_b(32'sd26),
  .signd_b(32'sd1),
  .width_z(32'sd49),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Tanh_for_3_else_else_mul_1_cmp (
      .a(23'b10101010101010101010101),
      .b(nl_Tanh_for_3_else_else_mul_1_cmp_b[25:0]),
      .clk(clk),
      .en(Tanh_for_3_else_else_mul_1_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_3_else_else_mul_1_cmp_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd23),
  .signd_a(32'sd1),
  .width_b(32'sd26),
  .signd_b(32'sd1),
  .width_z(32'sd49),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Tanh_for_3_else_else_mul_1_cmp_1 (
      .a(23'b10101010101010101010101),
      .b(nl_Tanh_for_3_else_else_mul_1_cmp_1_b[25:0]),
      .clk(clk),
      .en(Tanh_for_3_else_else_mul_1_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_3_else_else_mul_1_cmp_1_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd23),
  .signd_a(32'sd1),
  .width_b(32'sd26),
  .signd_b(32'sd1),
  .width_z(32'sd49),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Tanh_for_3_else_else_mul_1_cmp_2 (
      .a(23'b10101010101010101010101),
      .b(nl_Tanh_for_3_else_else_mul_1_cmp_2_b[25:0]),
      .clk(clk),
      .en(Tanh_for_3_else_else_mul_1_cmp_2_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_3_else_else_mul_1_cmp_2_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd23),
  .signd_a(32'sd1),
  .width_b(32'sd26),
  .signd_b(32'sd1),
  .width_z(32'sd49),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Tanh_for_3_else_else_mul_1_cmp_3 (
      .a(23'b10101010101010101010101),
      .b(nl_Tanh_for_3_else_else_mul_1_cmp_3_b[25:0]),
      .clk(clk),
      .en(Tanh_for_3_else_else_mul_1_cmp_3_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_3_else_else_mul_1_cmp_3_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd23),
  .signd_a(32'sd1),
  .width_b(32'sd26),
  .signd_b(32'sd1),
  .width_z(32'sd49),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Tanh_for_3_else_else_mul_1_cmp_4 (
      .a(23'b10101010101010101010101),
      .b(nl_Tanh_for_3_else_else_mul_1_cmp_4_b[25:0]),
      .clk(clk),
      .en(Tanh_for_3_else_else_mul_1_cmp_4_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_3_else_else_mul_1_cmp_4_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd23),
  .signd_a(32'sd1),
  .width_b(32'sd26),
  .signd_b(32'sd1),
  .width_z(32'sd49),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Tanh_for_3_else_else_mul_1_cmp_5 (
      .a(23'b10101010101010101010101),
      .b(nl_Tanh_for_3_else_else_mul_1_cmp_5_b[25:0]),
      .clk(clk),
      .en(Tanh_for_3_else_else_mul_1_cmp_5_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_3_else_else_mul_1_cmp_5_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd23),
  .signd_a(32'sd1),
  .width_b(32'sd26),
  .signd_b(32'sd1),
  .width_z(32'sd49),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Tanh_for_3_else_else_mul_1_cmp_6 (
      .a(23'b10101010101010101010101),
      .b(nl_Tanh_for_3_else_else_mul_1_cmp_6_b[25:0]),
      .clk(clk),
      .en(Tanh_for_3_else_else_mul_1_cmp_6_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_3_else_else_mul_1_cmp_6_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd23),
  .signd_a(32'sd1),
  .width_b(32'sd26),
  .signd_b(32'sd1),
  .width_z(32'sd49),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Tanh_for_3_else_else_mul_1_cmp_7 (
      .a(23'b10101010101010101010101),
      .b(nl_Tanh_for_3_else_else_mul_1_cmp_7_b[25:0]),
      .clk(clk),
      .en(Tanh_for_3_else_else_mul_1_cmp_7_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_3_else_else_mul_1_cmp_7_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd23),
  .signd_a(32'sd1),
  .width_b(32'sd26),
  .signd_b(32'sd1),
  .width_z(32'sd49),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Tanh_for_3_else_else_mul_1_cmp_8 (
      .a(23'b10101010101010101010101),
      .b(nl_Tanh_for_3_else_else_mul_1_cmp_8_b[25:0]),
      .clk(clk),
      .en(Tanh_for_3_else_else_mul_1_cmp_8_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_3_else_else_mul_1_cmp_8_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd23),
  .signd_a(32'sd1),
  .width_b(32'sd26),
  .signd_b(32'sd1),
  .width_z(32'sd49),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Tanh_for_3_else_else_mul_1_cmp_9 (
      .a(23'b10101010101010101010101),
      .b(nl_Tanh_for_3_else_else_mul_1_cmp_9_b[25:0]),
      .clk(clk),
      .en(Tanh_for_3_else_else_mul_1_cmp_9_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_3_else_else_mul_1_cmp_9_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd23),
  .signd_a(32'sd1),
  .width_b(32'sd26),
  .signd_b(32'sd1),
  .width_z(32'sd49),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Tanh_for_3_else_else_mul_1_cmp_10 (
      .a(23'b10101010101010101010101),
      .b(nl_Tanh_for_3_else_else_mul_1_cmp_10_b[25:0]),
      .clk(clk),
      .en(Tanh_for_3_else_else_mul_1_cmp_10_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_3_else_else_mul_1_cmp_10_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd23),
  .signd_a(32'sd1),
  .width_b(32'sd26),
  .signd_b(32'sd1),
  .width_z(32'sd49),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Tanh_for_3_else_else_mul_1_cmp_11 (
      .a(23'b10101010101010101010101),
      .b(nl_Tanh_for_3_else_else_mul_1_cmp_11_b[25:0]),
      .clk(clk),
      .en(Tanh_for_3_else_else_mul_1_cmp_11_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_3_else_else_mul_1_cmp_11_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd23),
  .signd_a(32'sd1),
  .width_b(32'sd26),
  .signd_b(32'sd1),
  .width_z(32'sd49),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Tanh_for_3_else_else_mul_1_cmp_12 (
      .a(23'b10101010101010101010101),
      .b(nl_Tanh_for_3_else_else_mul_1_cmp_12_b[25:0]),
      .clk(clk),
      .en(Tanh_for_3_else_else_mul_1_cmp_12_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_3_else_else_mul_1_cmp_12_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd23),
  .signd_a(32'sd1),
  .width_b(32'sd26),
  .signd_b(32'sd1),
  .width_z(32'sd49),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Tanh_for_3_else_else_mul_1_cmp_13 (
      .a(23'b10101010101010101010101),
      .b(nl_Tanh_for_3_else_else_mul_1_cmp_13_b[25:0]),
      .clk(clk),
      .en(Tanh_for_3_else_else_mul_1_cmp_13_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_3_else_else_mul_1_cmp_13_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd26),
  .signd_a(32'sd1),
  .width_b(32'sd75),
  .signd_b(32'sd1),
  .width_z(32'sd101),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd5),
  .n_inreg(32'sd1)) Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp (
      .a(reg_ActUnit_RunInst_case_11_nv_scvector_cctor_data_0_ftd_6),
      .b(Tanh_for_1_else_else_mul_cmp_z),
      .clk(clk),
      .en(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd26),
  .signd_a(32'sd1),
  .width_b(32'sd75),
  .signd_b(32'sd1),
  .width_z(32'sd101),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd5),
  .n_inreg(32'sd1)) Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_1 (
      .a(nl_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_1_a[25:0]),
      .b(Tanh_for_1_else_else_mul_cmp_1_z),
      .clk(clk),
      .en(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_1_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd26),
  .signd_a(32'sd1),
  .width_b(32'sd75),
  .signd_b(32'sd1),
  .width_z(32'sd101),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd5),
  .n_inreg(32'sd1)) Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_2 (
      .a(reg_nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6),
      .b(Tanh_for_1_else_else_mul_cmp_2_z),
      .clk(clk),
      .en(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_2_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_2_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd26),
  .signd_a(32'sd1),
  .width_b(32'sd75),
  .signd_b(32'sd1),
  .width_z(32'sd101),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd5),
  .n_inreg(32'sd1)) Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_3 (
      .a(reg_nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6),
      .b(Tanh_for_1_else_else_mul_cmp_3_z),
      .clk(clk),
      .en(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_3_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_3_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd26),
  .signd_a(32'sd1),
  .width_b(32'sd75),
  .signd_b(32'sd1),
  .width_z(32'sd101),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd5),
  .n_inreg(32'sd1)) Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_4 (
      .a(reg_nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6),
      .b(Tanh_for_1_else_else_mul_cmp_4_z),
      .clk(clk),
      .en(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_4_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_4_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd26),
  .signd_a(32'sd1),
  .width_b(32'sd75),
  .signd_b(32'sd1),
  .width_z(32'sd101),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd5),
  .n_inreg(32'sd1)) Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_5 (
      .a(reg_nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6),
      .b(Tanh_for_1_else_else_mul_cmp_5_z),
      .clk(clk),
      .en(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_5_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_5_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd26),
  .signd_a(32'sd1),
  .width_b(32'sd75),
  .signd_b(32'sd1),
  .width_z(32'sd101),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd5),
  .n_inreg(32'sd1)) Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_6 (
      .a(nl_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_6_a[25:0]),
      .b(Tanh_for_1_else_else_mul_cmp_6_z),
      .clk(clk),
      .en(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_6_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_6_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd26),
  .signd_a(32'sd1),
  .width_b(32'sd75),
  .signd_b(32'sd1),
  .width_z(32'sd101),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd5),
  .n_inreg(32'sd1)) Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_7 (
      .a(nl_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_7_a[25:0]),
      .b(Tanh_for_1_else_else_mul_cmp_7_z),
      .clk(clk),
      .en(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_7_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_7_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd26),
  .signd_a(32'sd1),
  .width_b(32'sd75),
  .signd_b(32'sd1),
  .width_z(32'sd101),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd5),
  .n_inreg(32'sd1)) Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_8 (
      .a(reg_nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6),
      .b(Tanh_for_1_else_else_mul_cmp_8_z),
      .clk(clk),
      .en(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_8_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_8_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd26),
  .signd_a(32'sd1),
  .width_b(32'sd75),
  .signd_b(32'sd1),
  .width_z(32'sd101),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd5),
  .n_inreg(32'sd1)) Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_9 (
      .a(reg_nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6),
      .b(Tanh_for_1_else_else_mul_cmp_9_z),
      .clk(clk),
      .en(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_9_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_9_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd26),
  .signd_a(32'sd1),
  .width_b(32'sd75),
  .signd_b(32'sd1),
  .width_z(32'sd101),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd5),
  .n_inreg(32'sd1)) Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_10 (
      .a(reg_nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6),
      .b(Tanh_for_1_else_else_mul_cmp_10_z),
      .clk(clk),
      .en(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_10_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_10_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd26),
  .signd_a(32'sd1),
  .width_b(32'sd75),
  .signd_b(32'sd1),
  .width_z(32'sd101),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd5),
  .n_inreg(32'sd1)) Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_11 (
      .a(reg_nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6),
      .b(Tanh_for_1_else_else_mul_cmp_11_z),
      .clk(clk),
      .en(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_11_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_11_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd26),
  .signd_a(32'sd1),
  .width_b(32'sd75),
  .signd_b(32'sd1),
  .width_z(32'sd101),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd5),
  .n_inreg(32'sd1)) Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_12 (
      .a(reg_nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6),
      .b(Tanh_for_1_else_else_mul_cmp_12_z),
      .clk(clk),
      .en(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_12_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_12_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd26),
  .signd_a(32'sd1),
  .width_b(32'sd75),
  .signd_b(32'sd1),
  .width_z(32'sd101),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd5),
  .n_inreg(32'sd1)) Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_13 (
      .a(reg_nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6),
      .b(Tanh_for_1_else_else_mul_cmp_13_z),
      .clk(clk),
      .en(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_13_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_13_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd26),
  .signd_a(32'sd1),
  .width_b(32'sd75),
  .signd_b(32'sd1),
  .width_z(32'sd101),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd5),
  .n_inreg(32'sd1)) Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_14 (
      .a(reg_nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6),
      .b(Tanh_for_1_else_else_mul_cmp_14_z),
      .clk(clk),
      .en(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_14_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_14_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd26),
  .signd_a(32'sd1),
  .width_b(32'sd75),
  .signd_b(32'sd1),
  .width_z(32'sd101),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd5),
  .n_inreg(32'sd1)) Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_15 (
      .a(reg_nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6),
      .b(Tanh_for_1_else_else_mul_cmp_15_z),
      .clk(clk),
      .en(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_15_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_15_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd26),
  .signd_a(32'sd1),
  .width_b(32'sd49),
  .signd_b(32'sd1),
  .width_z(32'sd75),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd4),
  .n_inreg(32'sd1)) Tanh_for_1_else_else_mul_cmp (
      .a(nl_Tanh_for_1_else_else_mul_cmp_a[25:0]),
      .b(nl_Tanh_for_1_else_else_mul_cmp_b[48:0]),
      .clk(clk),
      .en(Tanh_for_1_else_else_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_1_else_else_mul_cmp_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd26),
  .signd_a(32'sd1),
  .width_b(32'sd49),
  .signd_b(32'sd1),
  .width_z(32'sd75),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd4),
  .n_inreg(32'sd1)) Tanh_for_1_else_else_mul_cmp_1 (
      .a(nl_Tanh_for_1_else_else_mul_cmp_1_a[25:0]),
      .b(Tanh_for_3_else_else_mul_1_cmp_1_z),
      .clk(clk),
      .en(Tanh_for_1_else_else_mul_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_1_else_else_mul_cmp_1_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd26),
  .signd_a(32'sd1),
  .width_b(32'sd49),
  .signd_b(32'sd1),
  .width_z(32'sd75),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd4),
  .n_inreg(32'sd1)) Tanh_for_1_else_else_mul_cmp_2 (
      .a(reg_nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6),
      .b(Tanh_for_3_else_else_mul_1_cmp_2_z),
      .clk(clk),
      .en(Tanh_for_1_else_else_mul_cmp_2_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_1_else_else_mul_cmp_2_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd26),
  .signd_a(32'sd1),
  .width_b(32'sd49),
  .signd_b(32'sd1),
  .width_z(32'sd75),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd4),
  .n_inreg(32'sd1)) Tanh_for_1_else_else_mul_cmp_3 (
      .a(reg_nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6),
      .b(Tanh_for_3_else_else_mul_1_cmp_3_z),
      .clk(clk),
      .en(Tanh_for_1_else_else_mul_cmp_3_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_1_else_else_mul_cmp_3_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd26),
  .signd_a(32'sd1),
  .width_b(32'sd49),
  .signd_b(32'sd1),
  .width_z(32'sd75),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd4),
  .n_inreg(32'sd1)) Tanh_for_1_else_else_mul_cmp_4 (
      .a(reg_nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6),
      .b(Tanh_for_3_else_else_mul_1_cmp_4_z),
      .clk(clk),
      .en(Tanh_for_1_else_else_mul_cmp_4_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_1_else_else_mul_cmp_4_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd26),
  .signd_a(32'sd1),
  .width_b(32'sd49),
  .signd_b(32'sd1),
  .width_z(32'sd75),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd4),
  .n_inreg(32'sd1)) Tanh_for_1_else_else_mul_cmp_5 (
      .a(reg_nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6),
      .b(Tanh_for_3_else_else_mul_1_cmp_5_z),
      .clk(clk),
      .en(Tanh_for_1_else_else_mul_cmp_5_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_1_else_else_mul_cmp_5_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd26),
  .signd_a(32'sd1),
  .width_b(32'sd49),
  .signd_b(32'sd1),
  .width_z(32'sd75),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd4),
  .n_inreg(32'sd1)) Tanh_for_1_else_else_mul_cmp_6 (
      .a(nl_Tanh_for_1_else_else_mul_cmp_6_a[25:0]),
      .b(Tanh_for_3_else_else_mul_1_cmp_6_z),
      .clk(clk),
      .en(Tanh_for_1_else_else_mul_cmp_6_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_1_else_else_mul_cmp_6_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd26),
  .signd_a(32'sd1),
  .width_b(32'sd49),
  .signd_b(32'sd1),
  .width_z(32'sd75),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd4),
  .n_inreg(32'sd1)) Tanh_for_1_else_else_mul_cmp_7 (
      .a(nl_Tanh_for_1_else_else_mul_cmp_7_a[25:0]),
      .b(Tanh_for_3_else_else_mul_1_cmp_7_z),
      .clk(clk),
      .en(Tanh_for_1_else_else_mul_cmp_7_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_1_else_else_mul_cmp_7_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd26),
  .signd_a(32'sd1),
  .width_b(32'sd49),
  .signd_b(32'sd1),
  .width_z(32'sd75),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd4),
  .n_inreg(32'sd1)) Tanh_for_1_else_else_mul_cmp_8 (
      .a(reg_nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6),
      .b(Tanh_for_3_else_else_mul_1_cmp_8_z),
      .clk(clk),
      .en(Tanh_for_1_else_else_mul_cmp_8_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_1_else_else_mul_cmp_8_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd26),
  .signd_a(32'sd1),
  .width_b(32'sd49),
  .signd_b(32'sd1),
  .width_z(32'sd75),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd4),
  .n_inreg(32'sd1)) Tanh_for_1_else_else_mul_cmp_9 (
      .a(reg_nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6),
      .b(Tanh_for_3_else_else_mul_1_cmp_9_z),
      .clk(clk),
      .en(Tanh_for_1_else_else_mul_cmp_9_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_1_else_else_mul_cmp_9_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd26),
  .signd_a(32'sd1),
  .width_b(32'sd49),
  .signd_b(32'sd1),
  .width_z(32'sd75),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd4),
  .n_inreg(32'sd1)) Tanh_for_1_else_else_mul_cmp_10 (
      .a(reg_nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6),
      .b(Tanh_for_3_else_else_mul_1_cmp_10_z),
      .clk(clk),
      .en(Tanh_for_1_else_else_mul_cmp_10_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_1_else_else_mul_cmp_10_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd26),
  .signd_a(32'sd1),
  .width_b(32'sd49),
  .signd_b(32'sd1),
  .width_z(32'sd75),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd4),
  .n_inreg(32'sd1)) Tanh_for_1_else_else_mul_cmp_11 (
      .a(reg_nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6),
      .b(Tanh_for_3_else_else_mul_1_cmp_11_z),
      .clk(clk),
      .en(Tanh_for_1_else_else_mul_cmp_11_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_1_else_else_mul_cmp_11_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd26),
  .signd_a(32'sd1),
  .width_b(32'sd49),
  .signd_b(32'sd1),
  .width_z(32'sd75),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd4),
  .n_inreg(32'sd1)) Tanh_for_1_else_else_mul_cmp_12 (
      .a(nl_Tanh_for_1_else_else_mul_cmp_12_a[25:0]),
      .b(nl_Tanh_for_1_else_else_mul_cmp_12_b[48:0]),
      .clk(clk),
      .en(Tanh_for_1_else_else_mul_cmp_12_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_1_else_else_mul_cmp_12_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd26),
  .signd_a(32'sd1),
  .width_b(32'sd49),
  .signd_b(32'sd1),
  .width_z(32'sd75),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd4),
  .n_inreg(32'sd1)) Tanh_for_1_else_else_mul_cmp_13 (
      .a(nl_Tanh_for_1_else_else_mul_cmp_13_a[25:0]),
      .b(nl_Tanh_for_1_else_else_mul_cmp_13_b[48:0]),
      .clk(clk),
      .en(Tanh_for_1_else_else_mul_cmp_13_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_1_else_else_mul_cmp_13_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd26),
  .signd_a(32'sd1),
  .width_b(32'sd49),
  .signd_b(32'sd1),
  .width_z(32'sd75),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd4),
  .n_inreg(32'sd1)) Tanh_for_1_else_else_mul_cmp_14 (
      .a(nl_Tanh_for_1_else_else_mul_cmp_14_a[25:0]),
      .b(nl_Tanh_for_1_else_else_mul_cmp_14_b[48:0]),
      .clk(clk),
      .en(Tanh_for_1_else_else_mul_cmp_14_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_1_else_else_mul_cmp_14_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd26),
  .signd_a(32'sd1),
  .width_b(32'sd49),
  .signd_b(32'sd1),
  .width_z(32'sd75),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd4),
  .n_inreg(32'sd1)) Tanh_for_1_else_else_mul_cmp_15 (
      .a(nl_Tanh_for_1_else_else_mul_cmp_15_a[25:0]),
      .b(nl_Tanh_for_1_else_else_mul_cmp_15_b[48:0]),
      .clk(clk),
      .en(Tanh_for_1_else_else_mul_cmp_15_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_1_else_else_mul_cmp_15_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd27),
  .signd_a(32'sd1),
  .width_b(32'sd27),
  .signd_b(32'sd1),
  .width_z(32'sd54),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Tanh_for_1_else_else_mul_1_cmp (
      .a(nl_Tanh_for_1_else_else_mul_1_cmp_a[26:0]),
      .b(nl_Tanh_for_1_else_else_mul_1_cmp_b[26:0]),
      .clk(clk),
      .en(Tanh_for_1_else_else_mul_1_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_1_else_else_mul_1_cmp_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd27),
  .signd_a(32'sd1),
  .width_b(32'sd27),
  .signd_b(32'sd1),
  .width_z(32'sd54),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Tanh_for_1_else_else_mul_1_cmp_1 (
      .a(nl_Tanh_for_1_else_else_mul_1_cmp_1_a[26:0]),
      .b(nl_Tanh_for_1_else_else_mul_1_cmp_1_b[26:0]),
      .clk(clk),
      .en(Tanh_for_1_else_else_mul_1_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Tanh_for_1_else_else_mul_1_cmp_1_z)
    );
  ActUnit_ActUnit_ActUnitRun_rva_in_PopNB_mioi ActUnit_ActUnitRun_rva_in_PopNB_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_in_vld(rva_in_vld),
      .rva_in_rdy(rva_in_rdy),
      .rva_in_dat(rva_in_dat),
      .ActUnitRun_wen(ActUnitRun_wen),
      .ActUnitRun_wten(ActUnitRun_wten),
      .rva_in_PopNB_mioi_oswt(reg_rva_in_PopNB_mioi_iswt0_cse),
      .rva_in_PopNB_mioi_data_data_rsc_z_mxwt(rva_in_PopNB_mioi_data_data_rsc_z_mxwt),
      .rva_in_PopNB_mioi_data_addr_rsc_z_mxwt(rva_in_PopNB_mioi_data_addr_rsc_z_mxwt),
      .rva_in_PopNB_mioi_data_rw_rsc_z_mxwt(rva_in_PopNB_mioi_data_rw_rsc_z_mxwt),
      .rva_in_PopNB_mioi_return_rsc_z_mxwt(rva_in_PopNB_mioi_return_rsc_z_mxwt),
      .rva_in_PopNB_mioi_oswt_pff(and_837_rmff)
    );
  ActUnit_ActUnit_ActUnitRun_act_port_PopNB_mioi ActUnit_ActUnitRun_act_port_PopNB_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .act_port_vld(act_port_vld),
      .act_port_rdy(act_port_rdy),
      .act_port_dat(act_port_dat),
      .ActUnitRun_wen(ActUnitRun_wen),
      .ActUnitRun_wten(ActUnitRun_wten),
      .act_port_PopNB_mioi_oswt(reg_act_port_PopNB_mioi_iswt0_cse),
      .act_port_PopNB_mioi_data_data_rsc_z_mxwt(act_port_PopNB_mioi_data_data_rsc_z_mxwt),
      .act_port_PopNB_mioi_return_rsc_z_mxwt(act_port_PopNB_mioi_return_rsc_z_mxwt),
      .act_port_PopNB_mioi_oswt_pff(and_835_rmff)
    );
  ActUnit_ActUnit_ActUnitRun_rva_out_Push_mioi ActUnit_ActUnitRun_rva_out_Push_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_out_vld(rva_out_vld),
      .rva_out_rdy(rva_out_rdy),
      .rva_out_dat(rva_out_dat),
      .ActUnitRun_wten(nl_ActUnit_ActUnitRun_rva_out_Push_mioi_inst_ActUnitRun_wten),
      .rva_out_Push_mioi_oswt(reg_rva_out_Push_mioi_iswt0_cse),
      .rva_out_Push_mioi_wen_comp(rva_out_Push_mioi_wen_comp),
      .rva_out_Push_mioi_m_data_rsc_dat_ActUnitRun(nl_ActUnit_ActUnitRun_rva_out_Push_mioi_inst_rva_out_Push_mioi_m_data_rsc_dat_ActUnitRun[511:0]),
      .rva_out_Push_mioi_oswt_pff(and_830_rmff)
    );
  ActUnit_ActUnit_ActUnitRun_start_PopNB_mioi ActUnit_ActUnitRun_start_PopNB_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .start_vld(start_vld),
      .start_rdy(start_rdy),
      .start_dat(start_dat),
      .ActUnitRun_wen(ActUnitRun_wen),
      .ActUnitRun_wten(ActUnitRun_wten),
      .start_PopNB_mioi_oswt(reg_start_PopNB_mioi_iswt0_cse),
      .start_PopNB_mioi_data_rsc_z_mxwt(start_PopNB_mioi_data_rsc_z_mxwt),
      .start_PopNB_mioi_return_rsc_z_mxwt(start_PopNB_mioi_return_rsc_z_mxwt),
      .start_PopNB_mioi_oswt_pff(and_826_rmff)
    );
  ActUnit_ActUnit_ActUnitRun_output_port_Push_mioi ActUnit_ActUnitRun_output_port_Push_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .output_port_vld(output_port_vld),
      .output_port_rdy(output_port_rdy),
      .output_port_dat(output_port_dat),
      .ActUnitRun_wten(nl_ActUnit_ActUnitRun_output_port_Push_mioi_inst_ActUnitRun_wten),
      .output_port_Push_mioi_oswt(reg_output_port_Push_mioi_iswt0_cse),
      .output_port_Push_mioi_wen_comp(output_port_Push_mioi_wen_comp),
      .output_port_Push_mioi_m_data_data_rsc_dat_ActUnitRun(nl_ActUnit_ActUnitRun_output_port_Push_mioi_inst_output_port_Push_mioi_m_data_data_rsc_dat_ActUnitRun[511:0]),
      .output_port_Push_mioi_m_logical_addr_rsc_dat_ActUnitRun(nl_ActUnit_ActUnitRun_output_port_Push_mioi_inst_output_port_Push_mioi_m_logical_addr_rsc_dat_ActUnitRun[7:0]),
      .output_port_Push_mioi_oswt_pff(and_823_rmff)
    );
  ActUnit_ActUnit_ActUnitRun_done_Push_mioi ActUnit_ActUnitRun_done_Push_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .done_vld(done_vld),
      .done_rdy(done_rdy),
      .done_dat(done_dat),
      .ActUnitRun_wten(nl_ActUnit_ActUnitRun_done_Push_mioi_inst_ActUnitRun_wten),
      .done_Push_mioi_oswt(reg_done_Push_mioi_iswt0_cse),
      .done_Push_mioi_wen_comp(done_Push_mioi_wen_comp),
      .done_Push_mioi_oswt_pff(and_819_rmff)
    );
  ActUnit_ActUnit_ActUnitRun_wait_dp ActUnit_ActUnitRun_wait_dp_inst (
      .ActUnitRun_wen(ActUnitRun_wen),
      .Tanh_for_3_else_else_mul_1_cmp_cgo(reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_cse),
      .Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg(and_812_rmff),
      .Tanh_for_3_else_else_mul_1_cmp_en(Tanh_for_3_else_else_mul_1_cmp_en),
      .Tanh_for_3_else_else_mul_1_cmp_cgo_1(reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_1_cse),
      .Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_1(and_811_rmff),
      .Tanh_for_3_else_else_mul_1_cmp_1_en(Tanh_for_3_else_else_mul_1_cmp_1_en),
      .Tanh_for_3_else_else_mul_1_cmp_cgo_2(reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_2_cse),
      .Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_2(and_810_rmff),
      .Tanh_for_3_else_else_mul_1_cmp_2_en(Tanh_for_3_else_else_mul_1_cmp_2_en),
      .Tanh_for_3_else_else_mul_1_cmp_cgo_3(reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_3_cse),
      .Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_3(and_809_rmff),
      .Tanh_for_3_else_else_mul_1_cmp_3_en(Tanh_for_3_else_else_mul_1_cmp_3_en),
      .Tanh_for_3_else_else_mul_1_cmp_cgo_4(reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_4_cse),
      .Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_4(and_808_rmff),
      .Tanh_for_3_else_else_mul_1_cmp_4_en(Tanh_for_3_else_else_mul_1_cmp_4_en),
      .Tanh_for_3_else_else_mul_1_cmp_cgo_5(reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_5_cse),
      .Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_5(and_807_rmff),
      .Tanh_for_3_else_else_mul_1_cmp_5_en(Tanh_for_3_else_else_mul_1_cmp_5_en),
      .Tanh_for_3_else_else_mul_1_cmp_cgo_6(reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_6_cse),
      .Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_6(and_806_rmff),
      .Tanh_for_3_else_else_mul_1_cmp_6_en(Tanh_for_3_else_else_mul_1_cmp_6_en),
      .Tanh_for_3_else_else_mul_1_cmp_cgo_7(reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_7_cse),
      .Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_7(and_805_rmff),
      .Tanh_for_3_else_else_mul_1_cmp_7_en(Tanh_for_3_else_else_mul_1_cmp_7_en),
      .Tanh_for_3_else_else_mul_1_cmp_cgo_8(reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_8_cse),
      .Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_8(and_804_rmff),
      .Tanh_for_3_else_else_mul_1_cmp_8_en(Tanh_for_3_else_else_mul_1_cmp_8_en),
      .Tanh_for_3_else_else_mul_1_cmp_cgo_9(reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_9_cse),
      .Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_9(and_803_rmff),
      .Tanh_for_3_else_else_mul_1_cmp_9_en(Tanh_for_3_else_else_mul_1_cmp_9_en),
      .Tanh_for_3_else_else_mul_1_cmp_cgo_10(reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_10_cse),
      .Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_10(and_802_rmff),
      .Tanh_for_3_else_else_mul_1_cmp_10_en(Tanh_for_3_else_else_mul_1_cmp_10_en),
      .Tanh_for_3_else_else_mul_1_cmp_cgo_11(reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_11_cse),
      .Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_11(and_801_rmff),
      .Tanh_for_3_else_else_mul_1_cmp_11_en(Tanh_for_3_else_else_mul_1_cmp_11_en),
      .Tanh_for_3_else_else_mul_1_cmp_cgo_12(reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_12_cse),
      .Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_12(and_800_rmff),
      .Tanh_for_3_else_else_mul_1_cmp_12_en(Tanh_for_3_else_else_mul_1_cmp_12_en),
      .Tanh_for_3_else_else_mul_1_cmp_cgo_13(reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_13_cse),
      .Tanh_for_3_else_else_mul_1_cmp_cgo_ir_unreg_13(and_799_rmff),
      .Tanh_for_3_else_else_mul_1_cmp_13_en(Tanh_for_3_else_else_mul_1_cmp_13_en),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo(reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_cse),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg(and_794_rmff),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_en(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_en),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_1(reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_1_cse),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_1(and_789_rmff),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_1_en(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_1_en),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_2(reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_2_cse),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_2(and_784_rmff),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_2_en(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_2_en),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_3(reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_3_cse),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_3(and_779_rmff),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_3_en(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_3_en),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_4(reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_4_cse),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_4(and_774_rmff),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_4_en(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_4_en),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_5(reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_5_cse),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_5(and_769_rmff),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_5_en(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_5_en),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_6(reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_6_cse),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_6(and_764_rmff),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_6_en(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_6_en),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_7(reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_7_cse),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_7(and_759_rmff),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_7_en(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_7_en),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_8(reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_8_cse),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_8(and_754_rmff),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_8_en(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_8_en),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_9(reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_9_cse),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_9(and_749_rmff),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_9_en(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_9_en),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_10(reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_10_cse),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_10(and_744_rmff),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_10_en(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_10_en),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_11(reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_11_cse),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_11(and_739_rmff),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_11_en(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_11_en),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_12(reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_12_cse),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_12(and_734_rmff),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_12_en(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_12_en),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_13(reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_13_cse),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_13(and_729_rmff),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_13_en(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_13_en),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_14(reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_14_cse),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_14(and_724_rmff),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_14_en(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_14_en),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_15(reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_15_cse),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_unreg_15(and_719_rmff),
      .Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_15_en(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_15_en),
      .Tanh_for_1_else_else_mul_cmp_cgo(reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_cse),
      .Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg(and_713_rmff),
      .Tanh_for_1_else_else_mul_cmp_en(Tanh_for_1_else_else_mul_cmp_en),
      .Tanh_for_1_else_else_mul_cmp_cgo_1(reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_1_cse),
      .Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_1(and_705_rmff),
      .Tanh_for_1_else_else_mul_cmp_1_en(Tanh_for_1_else_else_mul_cmp_1_en),
      .Tanh_for_1_else_else_mul_cmp_cgo_2(reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_2_cse),
      .Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_2(and_701_rmff),
      .Tanh_for_1_else_else_mul_cmp_2_en(Tanh_for_1_else_else_mul_cmp_2_en),
      .Tanh_for_1_else_else_mul_cmp_cgo_3(reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_3_cse),
      .Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_3(and_697_rmff),
      .Tanh_for_1_else_else_mul_cmp_3_en(Tanh_for_1_else_else_mul_cmp_3_en),
      .Tanh_for_1_else_else_mul_cmp_cgo_4(reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_4_cse),
      .Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_4(and_693_rmff),
      .Tanh_for_1_else_else_mul_cmp_4_en(Tanh_for_1_else_else_mul_cmp_4_en),
      .Tanh_for_1_else_else_mul_cmp_cgo_5(reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_5_cse),
      .Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_5(and_689_rmff),
      .Tanh_for_1_else_else_mul_cmp_5_en(Tanh_for_1_else_else_mul_cmp_5_en),
      .Tanh_for_1_else_else_mul_cmp_cgo_6(reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_6_cse),
      .Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_6(and_685_rmff),
      .Tanh_for_1_else_else_mul_cmp_6_en(Tanh_for_1_else_else_mul_cmp_6_en),
      .Tanh_for_1_else_else_mul_cmp_cgo_7(reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_7_cse),
      .Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_7(and_681_rmff),
      .Tanh_for_1_else_else_mul_cmp_7_en(Tanh_for_1_else_else_mul_cmp_7_en),
      .Tanh_for_1_else_else_mul_cmp_cgo_8(reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_8_cse),
      .Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_8(and_677_rmff),
      .Tanh_for_1_else_else_mul_cmp_8_en(Tanh_for_1_else_else_mul_cmp_8_en),
      .Tanh_for_1_else_else_mul_cmp_cgo_9(reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_9_cse),
      .Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_9(and_673_rmff),
      .Tanh_for_1_else_else_mul_cmp_9_en(Tanh_for_1_else_else_mul_cmp_9_en),
      .Tanh_for_1_else_else_mul_cmp_cgo_10(reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_10_cse),
      .Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_10(and_669_rmff),
      .Tanh_for_1_else_else_mul_cmp_10_en(Tanh_for_1_else_else_mul_cmp_10_en),
      .Tanh_for_1_else_else_mul_cmp_cgo_11(reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_11_cse),
      .Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_11(and_665_rmff),
      .Tanh_for_1_else_else_mul_cmp_11_en(Tanh_for_1_else_else_mul_cmp_11_en),
      .Tanh_for_1_else_else_mul_cmp_cgo_12(reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_12_cse),
      .Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_12(and_658_rmff),
      .Tanh_for_1_else_else_mul_cmp_12_en(Tanh_for_1_else_else_mul_cmp_12_en),
      .Tanh_for_1_else_else_mul_cmp_cgo_13(reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_13_cse),
      .Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_13(and_633_rmff),
      .Tanh_for_1_else_else_mul_cmp_13_en(Tanh_for_1_else_else_mul_cmp_13_en),
      .Tanh_for_1_else_else_mul_cmp_cgo_14(reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_14_cse),
      .Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_14(and_626_rmff),
      .Tanh_for_1_else_else_mul_cmp_14_en(Tanh_for_1_else_else_mul_cmp_14_en),
      .Tanh_for_1_else_else_mul_cmp_cgo_15(reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_15_cse),
      .Tanh_for_1_else_else_mul_cmp_cgo_ir_unreg_15(and_621_rmff),
      .Tanh_for_1_else_else_mul_cmp_15_en(Tanh_for_1_else_else_mul_cmp_15_en),
      .Tanh_for_1_else_else_mul_1_cmp_cgo(reg_Tanh_for_1_else_else_mul_1_cmp_cgo_ir_cse),
      .Tanh_for_1_else_else_mul_1_cmp_cgo_ir_unreg(and_617_rmff),
      .Tanh_for_1_else_else_mul_1_cmp_en(Tanh_for_1_else_else_mul_1_cmp_en),
      .Tanh_for_1_else_else_mul_1_cmp_cgo_1(reg_Tanh_for_1_else_else_mul_1_cmp_cgo_ir_1_cse),
      .Tanh_for_1_else_else_mul_1_cmp_cgo_ir_unreg_1(and_605_rmff),
      .Tanh_for_1_else_else_mul_1_cmp_1_en(Tanh_for_1_else_else_mul_1_cmp_1_en)
    );
  ActUnit_ActUnit_ActUnitRun_staller ActUnit_ActUnitRun_staller_inst (
      .clk(clk),
      .rst(rst),
      .ActUnitRun_wen(ActUnitRun_wen),
      .ActUnitRun_wten(ActUnitRun_wten),
      .rva_out_Push_mioi_wen_comp(rva_out_Push_mioi_wen_comp),
      .output_port_Push_mioi_wen_comp(output_port_Push_mioi_wen_comp),
      .done_Push_mioi_wen_comp(done_Push_mioi_wen_comp)
    );
  ActUnit_ActUnit_ActUnitRun_ActUnitRun_fsm ActUnit_ActUnitRun_ActUnitRun_fsm_inst
      (
      .clk(clk),
      .rst(rst),
      .ActUnitRun_wen(ActUnitRun_wen),
      .fsm_output(fsm_output),
      .while_C_0_tr0(nl_ActUnit_ActUnitRun_ActUnitRun_fsm_inst_while_C_0_tr0),
      .ActUnit_RunInst_case_2_for_C_0_tr0(nl_ActUnit_ActUnitRun_ActUnitRun_fsm_inst_ActUnit_RunInst_case_2_for_C_0_tr0),
      .while_C_11_tr0(nl_ActUnit_ActUnitRun_ActUnitRun_fsm_inst_while_C_11_tr0),
      .ActUnit_PushOutput_if_for_C_0_tr0(nl_ActUnit_ActUnitRun_ActUnitRun_fsm_inst_ActUnit_PushOutput_if_for_C_0_tr0),
      .while_C_13_tr0(nl_ActUnit_ActUnitRun_ActUnitRun_fsm_inst_while_C_13_tr0),
      .ActUnit_RunLoad_if_else_for_C_0_tr0(nl_ActUnit_ActUnitRun_ActUnitRun_fsm_inst_ActUnit_RunLoad_if_else_for_C_0_tr0)
    );
  assign act_mem_banks_write_if_for_if_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_369);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb = act_mem_banks_write_if_for_if_mux_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl default clock = (posedge clk);
  // psl ActUnit_ActUnitRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb );
  assign act_mem_banks_write_if_for_if_mux_1_cse = MUX1HOT_s_1_1_2(ActUnitRun_wen,
      and_dcpl_369);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb = act_mem_banks_write_if_for_if_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb = act_mem_banks_write_if_for_if_mux_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl ActUnit_ActUnitRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb = act_mem_banks_write_if_for_if_mux_1_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb
      = act_mem_banks_write_if_for_if_mux_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl ActUnit_ActUnitRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb
      = act_mem_banks_write_if_for_if_mux_1_cse;
  assign act_mem_banks_read_for_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_374);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_1 = act_mem_banks_read_for_mux_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl ActUnit_ActUnitRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_1  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_1 );
  assign act_mem_banks_read_for_mux_1_cse = MUX1HOT_s_1_1_2(ActUnitRun_wen, and_dcpl_374);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_1 = act_mem_banks_read_for_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_1 = act_mem_banks_read_for_mux_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl ActUnit_ActUnitRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_1  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_1 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_1 = act_mem_banks_read_for_mux_1_cse;
  assign nand_6_nl = ~(nor_333_cse & not_tmp_248);
  assign nand_5_nl = ~(nor_28_cse & not_tmp_248);
  assign or_442_nl = (~ (fsm_output[0])) | Tanh_for_2_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | Tanh_for_2_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs;
  assign mux_110_nl = MUX_s_1_2_2(nand_tmp_3, or_442_nl, fsm_output[1]);
  assign or_443_nl = (fsm_output[2]) | mux_110_nl;
  assign mux_111_nl = MUX_s_1_2_2(nand_5_nl, or_443_nl, act_config_in_InstFetch_return_sva_7_2[2]);
  assign nand_4_nl = ~((fsm_output[0]) & (~((Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
      | Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      & or_tmp_151)));
  assign mux_107_nl = MUX_s_1_2_2(nand_tmp_3, nand_4_nl, fsm_output[1]);
  assign and_603_nl = or_tmp_148 & or_tmp_151;
  assign and_602_nl = or_tmp_148 & or_tmp_147;
  assign mux_105_nl = MUX_s_1_2_2(and_603_nl, and_602_nl, fsm_output[0]);
  assign and_601_nl = or_tmp_147 & or_tmp_146;
  assign and_600_nl = or_tmp_131 & or_tmp_146;
  assign mux_104_nl = MUX_s_1_2_2(and_601_nl, and_600_nl, fsm_output[0]);
  assign mux_106_nl = MUX_s_1_2_2(mux_105_nl, mux_104_nl, fsm_output[1]);
  assign mux_108_nl = MUX_s_1_2_2(mux_107_nl, mux_106_nl, fsm_output[2]);
  assign nand_2_nl = ~((fsm_output[0]) & (~ and_tmp_11));
  assign mux_102_nl = MUX_s_1_2_2(nand_tmp_3, nand_2_nl, fsm_output[1]);
  assign and_598_nl = or_tmp_136 & or_tmp_139;
  assign mux_99_nl = MUX_s_1_2_2(and_598_nl, and_tmp_9, fsm_output[0]);
  assign and_596_nl = or_tmp_135 & or_tmp_134;
  assign and_595_nl = or_tmp_133 & or_tmp_134;
  assign mux_98_nl = MUX_s_1_2_2(and_596_nl, and_595_nl, fsm_output[0]);
  assign mux_100_nl = MUX_s_1_2_2(mux_99_nl, mux_98_nl, fsm_output[1]);
  assign mux_103_nl = MUX_s_1_2_2(mux_102_nl, mux_100_nl, fsm_output[2]);
  assign mux_109_nl = MUX_s_1_2_2(mux_108_nl, mux_103_nl, act_config_in_InstFetch_return_sva_7_2[2]);
  assign mux_112_nl = MUX_s_1_2_2(mux_111_nl, mux_109_nl, act_config_in_InstFetch_return_sva_7_2[4]);
  assign or_419_nl = Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
      | Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign mux_95_nl = MUX_s_1_2_2(or_tmp_131, or_419_nl, fsm_output[0]);
  assign and_594_nl = (Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
      | Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      & mux_95_nl;
  assign or_417_nl = (fsm_output[0]) | Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
      | Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign mux_96_nl = MUX_s_1_2_2(and_594_nl, or_417_nl, fsm_output[1]);
  assign nor_160_nl = ~((fsm_output[2]) | mux_96_nl);
  assign nor_161_nl = ~((fsm_output[2:0]!=3'b000) | Tanh_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
      | Tanh_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
  assign mux_97_nl = MUX_s_1_2_2(nor_160_nl, nor_161_nl, act_config_in_InstFetch_return_sva_7_2[2]);
  assign nand_1_nl = ~((act_config_in_InstFetch_return_sva_7_2[4]) & mux_97_nl);
  assign mux_113_nl = MUX_s_1_2_2(mux_112_nl, nand_1_nl, fsm_output[3]);
  assign mux_114_nl = MUX_s_1_2_2(nand_6_nl, mux_113_nl, and_1101_cse);
  assign and_605_rmff = (~ mux_114_nl) & and_dcpl_587;
  assign nand_12_nl = ~(nor_333_cse & not_tmp_255);
  assign nand_11_nl = ~(nor_28_cse & not_tmp_255);
  assign or_470_nl = (~ (fsm_output[0])) | Tanh_for_1_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | Tanh_for_1_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs;
  assign mux_130_nl = MUX_s_1_2_2(nand_tmp_9, or_470_nl, fsm_output[1]);
  assign or_471_nl = (fsm_output[2]) | mux_130_nl;
  assign mux_131_nl = MUX_s_1_2_2(nand_11_nl, or_471_nl, act_config_in_InstFetch_return_sva_7_2[2]);
  assign nand_10_nl = ~((fsm_output[0]) & (~((Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
      | Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      & or_tmp_179)));
  assign mux_127_nl = MUX_s_1_2_2(nand_tmp_9, nand_10_nl, fsm_output[1]);
  assign and_615_nl = or_tmp_176 & or_tmp_179;
  assign and_614_nl = or_tmp_176 & or_tmp_175;
  assign mux_125_nl = MUX_s_1_2_2(and_615_nl, and_614_nl, fsm_output[0]);
  assign and_613_nl = or_tmp_175 & or_tmp_174;
  assign and_612_nl = or_tmp_159 & or_tmp_174;
  assign mux_124_nl = MUX_s_1_2_2(and_613_nl, and_612_nl, fsm_output[0]);
  assign mux_126_nl = MUX_s_1_2_2(mux_125_nl, mux_124_nl, fsm_output[1]);
  assign mux_128_nl = MUX_s_1_2_2(mux_127_nl, mux_126_nl, fsm_output[2]);
  assign nand_8_nl = ~((fsm_output[0]) & (~(or_tmp_168 & or_tmp_167)));
  assign mux_122_nl = MUX_s_1_2_2(nand_tmp_9, nand_8_nl, fsm_output[1]);
  assign and_610_nl = or_tmp_164 & or_tmp_167;
  assign and_609_nl = or_tmp_164 & or_tmp_163;
  assign mux_119_nl = MUX_s_1_2_2(and_610_nl, and_609_nl, fsm_output[0]);
  assign and_608_nl = or_tmp_163 & or_tmp_162;
  assign and_607_nl = or_tmp_161 & or_tmp_162;
  assign mux_118_nl = MUX_s_1_2_2(and_608_nl, and_607_nl, fsm_output[0]);
  assign mux_120_nl = MUX_s_1_2_2(mux_119_nl, mux_118_nl, fsm_output[1]);
  assign mux_123_nl = MUX_s_1_2_2(mux_122_nl, mux_120_nl, fsm_output[2]);
  assign mux_129_nl = MUX_s_1_2_2(mux_128_nl, mux_123_nl, act_config_in_InstFetch_return_sva_7_2[2]);
  assign mux_132_nl = MUX_s_1_2_2(mux_131_nl, mux_129_nl, act_config_in_InstFetch_return_sva_7_2[4]);
  assign or_447_nl = Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
      | Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign mux_115_nl = MUX_s_1_2_2(or_tmp_159, or_447_nl, fsm_output[0]);
  assign and_606_nl = (Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
      | Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      & mux_115_nl;
  assign or_445_nl = (fsm_output[0]) | Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
      | Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign mux_116_nl = MUX_s_1_2_2(and_606_nl, or_445_nl, fsm_output[1]);
  assign nor_162_nl = ~((fsm_output[2]) | mux_116_nl);
  assign nor_163_nl = ~((fsm_output[2:0]!=3'b000) | Tanh_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
      | Tanh_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
  assign mux_117_nl = MUX_s_1_2_2(nor_162_nl, nor_163_nl, act_config_in_InstFetch_return_sva_7_2[2]);
  assign nand_7_nl = ~((act_config_in_InstFetch_return_sva_7_2[4]) & mux_117_nl);
  assign mux_133_nl = MUX_s_1_2_2(mux_132_nl, nand_7_nl, fsm_output[3]);
  assign mux_134_nl = MUX_s_1_2_2(nand_12_nl, mux_133_nl, and_1101_cse);
  assign and_617_rmff = (~ mux_134_nl) & and_dcpl_587;
  assign or_477_nl = (~ (fsm_output[0])) | operator_32_8_true_AC_TRN_AC_WRAP_2_less_3_tmp_1
      | operator_32_8_true_AC_TRN_AC_WRAP_3_less_3_tmp | (act_config_in_InstFetch_mux_tmp[7:4]!=4'b1111)
      | (fsm_output[1]) | (fsm_output[3]);
  assign or_476_nl = Tanh_for_2_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | Tanh_for_2_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
      | (fsm_output[3]);
  assign mux_138_nl = MUX_s_1_2_2(or_477_nl, or_476_nl, fsm_output[2]);
  assign or_475_nl = (~(operator_32_8_true_AC_TRN_AC_WRAP_2_less_3_tmp_1 | operator_32_8_true_AC_TRN_AC_WRAP_3_less_3_tmp
      | (act_config_in_InstFetch_mux_tmp[7:4]!=4'b1111))) | (fsm_output[1]) | (fsm_output[3]);
  assign mux_135_nl = MUX_s_1_2_2((fsm_output[3]), or_475_nl, fsm_output[0]);
  assign or_474_nl = (fsm_output[1]) | (fsm_output[3]);
  assign mux_136_nl = MUX_s_1_2_2((~ mux_135_nl), or_474_nl, fsm_output[2]);
  assign or_472_nl = Gelu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
      | Gelu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs;
  assign mux_137_nl = MUX_s_1_2_2(mux_136_nl, or_tmp_184, or_472_nl);
  assign mux_139_nl = MUX_s_1_2_2(mux_138_nl, mux_137_nl, act_config_in_InstFetch_return_sva_7_2[4]);
  assign mux_140_nl = MUX_s_1_2_2(or_tmp_184, mux_139_nl, and_1103_cse);
  assign and_621_rmff = (~ mux_140_nl) & and_dcpl_587;
  assign nor_164_nl = ~((~ (fsm_output[3])) | Gelu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      | Gelu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
      | (~ (act_config_in_InstFetch_return_sva_7_2[4])));
  assign nor_165_nl = ~((fsm_output[3]) | Tanh_for_3_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | Tanh_for_3_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
      | (act_config_in_InstFetch_return_sva_7_2[4]));
  assign mux_141_nl = MUX_s_1_2_2(nor_164_nl, nor_165_nl, fsm_output[2]);
  assign and_626_rmff = mux_141_nl & and_dcpl_596 & (act_config_in_InstFetch_return_sva_7_2[2])
      & (~ (fsm_output[4]));
  assign or_499_nl = (fsm_output[3:0]!=4'b0001) | operator_32_8_true_AC_TRN_AC_WRAP_2_less_tmp_1
      | operator_32_8_true_AC_TRN_AC_WRAP_3_less_tmp | not_tmp_262;
  assign or_496_nl = Tanh_for_4_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | Tanh_for_4_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs;
  assign mux_149_nl = MUX_s_1_2_2(or_tmp_198, or_496_nl, fsm_output[2]);
  assign or_497_nl = (fsm_output[3]) | mux_149_nl;
  assign nand_207_nl = ~((fsm_output[0]) & ((fsm_output[1]) | (~(operator_32_8_true_AC_TRN_AC_WRAP_2_less_tmp_1
      | operator_32_8_true_AC_TRN_AC_WRAP_3_less_tmp | not_tmp_262))));
  assign and_631_nl = (fsm_output[1]) & or_tmp_167;
  assign mux_145_nl = MUX_s_1_2_2((fsm_output[1]), and_631_nl, fsm_output[0]);
  assign mux_146_nl = MUX_s_1_2_2(nand_207_nl, mux_145_nl, fsm_output[2]);
  assign nor_167_nl = ~((fsm_output[1:0]!=2'b00) | (~(or_tmp_167 & or_tmp_134)));
  assign mux_144_nl = MUX_s_1_2_2(nor_167_nl, or_992_cse, fsm_output[2]);
  assign mux_147_nl = MUX_s_1_2_2(mux_146_nl, mux_144_nl, fsm_output[3]);
  assign or_485_nl = (fsm_output[1:0]!=2'b11) | Gelu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
      | Gelu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs;
  assign mux_142_nl = MUX_s_1_2_2(or_tmp_198, or_485_nl, fsm_output[2]);
  assign or_484_nl = (fsm_output[2]) | ((and_1104_cse | Gelu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
      | Gelu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & or_tmp_134);
  assign mux_143_nl = MUX_s_1_2_2(mux_142_nl, or_484_nl, fsm_output[3]);
  assign or_481_nl = Tanh_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
      | Tanh_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  assign mux_148_nl = MUX_s_1_2_2(mux_147_nl, mux_143_nl, or_481_nl);
  assign mux_150_nl = MUX_s_1_2_2(or_497_nl, mux_148_nl, act_config_in_InstFetch_return_sva_7_2[4]);
  assign mux_151_nl = MUX_s_1_2_2(or_499_nl, mux_150_nl, and_1103_cse);
  assign and_633_rmff = (~ mux_151_nl) & and_dcpl_587;
  assign nor_171_nl = ~((fsm_output[3:0]!=4'b0001) | operator_32_8_true_AC_TRN_AC_WRAP_2_less_1_tmp_1
      | operator_32_8_true_AC_TRN_AC_WRAP_3_less_1_tmp | not_tmp_262);
  assign or_522_nl = Tanh_for_5_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | Tanh_for_5_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs;
  assign mux_163_nl = MUX_s_1_2_2(or_tmp_229, or_522_nl, fsm_output[2]);
  assign nor_172_nl = ~((fsm_output[3]) | mux_163_nl);
  assign nor_170_nl = ~((~ (fsm_output[0])) | operator_32_8_true_AC_TRN_AC_WRAP_2_less_1_tmp_1
      | operator_32_8_true_AC_TRN_AC_WRAP_3_less_1_tmp | not_tmp_262);
  assign mux_159_nl = MUX_s_1_2_2(nor_170_nl, (fsm_output[0]), fsm_output[1]);
  assign nand_209_nl = ~((fsm_output[1]) & and_tmp_39);
  assign mux_160_nl = MUX_s_1_2_2(mux_159_nl, nand_209_nl, fsm_output[2]);
  assign nand_210_nl = ~((fsm_output[2]) & or_tmp_215);
  assign mux_161_nl = MUX_s_1_2_2(mux_160_nl, nand_210_nl, fsm_output[3]);
  assign and_655_nl = ((~ (fsm_output[0])) | Gelu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
      | Gelu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & or_tmp_140;
  assign mux_156_nl = MUX_s_1_2_2(and_655_nl, and_tmp_39, fsm_output[1]);
  assign mux_157_nl = MUX_s_1_2_2(or_tmp_229, mux_156_nl, fsm_output[2]);
  assign and_651_nl = or_tmp_163 & or_tmp_164 & or_tmp_139;
  assign and_649_nl = or_tmp_163 & or_tmp_164 & or_tmp_161;
  assign mux_153_nl = MUX_s_1_2_2(and_651_nl, and_649_nl, fsm_output[0]);
  assign and_647_nl = ((fsm_output[0]) | Gelu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
      | Gelu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & or_tmp_161;
  assign mux_154_nl = MUX_s_1_2_2(mux_153_nl, and_647_nl, fsm_output[1]);
  assign mux_155_nl = MUX_s_1_2_2(mux_154_nl, or_tmp_215, fsm_output[2]);
  assign mux_158_nl = MUX_s_1_2_2(mux_157_nl, mux_155_nl, fsm_output[3]);
  assign or_504_nl = Gelu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
      | Gelu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs;
  assign mux_162_nl = MUX_s_1_2_2(mux_161_nl, (~ mux_158_nl), or_504_nl);
  assign mux_164_nl = MUX_s_1_2_2(nor_172_nl, mux_162_nl, act_config_in_InstFetch_return_sva_7_2[4]);
  assign mux_165_nl = MUX_s_1_2_2(nor_171_nl, mux_164_nl, and_1103_cse);
  assign and_658_rmff = mux_165_nl & and_dcpl_587;
  assign and_665_rmff = and_dcpl_621 & (~(Tanh_for_6_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
      | Tanh_for_6_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | (fsm_output[3]))) & and_dcpl_616;
  assign and_669_rmff = and_dcpl_621 & (~(Tanh_for_7_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
      | Tanh_for_7_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | (fsm_output[3]))) & and_dcpl_616;
  assign and_673_rmff = and_dcpl_621 & (~(Tanh_for_8_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
      | Tanh_for_8_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | (fsm_output[3]))) & and_dcpl_616;
  assign and_677_rmff = and_dcpl_621 & (~(Tanh_for_9_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
      | Tanh_for_9_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | (fsm_output[3]))) & and_dcpl_616;
  assign and_681_rmff = and_dcpl_621 & (~(Tanh_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
      | Tanh_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | (fsm_output[3]))) & and_dcpl_616;
  assign and_685_rmff = and_dcpl_621 & (~(Tanh_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
      | Tanh_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | (fsm_output[3]))) & and_dcpl_616;
  assign and_689_rmff = and_dcpl_621 & (~(Tanh_for_12_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
      | Tanh_for_12_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | (fsm_output[3]))) & and_dcpl_616;
  assign and_693_rmff = and_dcpl_621 & (~(Tanh_for_13_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
      | Tanh_for_13_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | (fsm_output[3]))) & and_dcpl_616;
  assign and_697_rmff = and_dcpl_621 & (~(Tanh_for_14_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
      | Tanh_for_14_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | (fsm_output[3]))) & and_dcpl_616;
  assign and_701_rmff = and_dcpl_621 & (~(Tanh_for_15_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
      | Tanh_for_15_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | (fsm_output[3]))) & and_dcpl_616;
  assign and_705_rmff = and_dcpl_621 & (~(Tanh_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
      | Tanh_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | (fsm_output[3]))) & and_dcpl_616;
  assign Tanh_for_else_else_or_1_cse = and_dcpl_604 | and_dcpl_612;
  assign nor_197_nl = ~((fsm_output[3:0]!=4'b0001) | operator_32_8_true_AC_TRN_AC_WRAP_2_less_2_tmp_1
      | operator_32_8_true_AC_TRN_AC_WRAP_3_less_2_tmp | not_tmp_262);
  assign or_542_nl = Tanh_for_1_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | Tanh_for_1_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs;
  assign mux_177_nl = MUX_s_1_2_2(or_tmp_249, or_542_nl, fsm_output[2]);
  assign nor_198_nl = ~((fsm_output[3]) | mux_177_nl);
  assign nor_195_nl = ~((~ (fsm_output[0])) | operator_32_8_true_AC_TRN_AC_WRAP_2_less_2_tmp_1
      | operator_32_8_true_AC_TRN_AC_WRAP_3_less_2_tmp | not_tmp_262);
  assign mux_173_nl = MUX_s_1_2_2(nor_195_nl, (fsm_output[0]), fsm_output[1]);
  assign nand_211_nl = ~((fsm_output[1]) & mux_tmp_169);
  assign mux_174_nl = MUX_s_1_2_2(mux_173_nl, nand_211_nl, fsm_output[2]);
  assign nand_212_nl = ~((fsm_output[2]) & or_tmp_237);
  assign mux_175_nl = MUX_s_1_2_2(mux_174_nl, nand_212_nl, fsm_output[3]);
  assign mux_170_nl = MUX_s_1_2_2(or_tmp_168, mux_tmp_169, fsm_output[1]);
  assign mux_171_nl = MUX_s_1_2_2(or_tmp_249, mux_170_nl, fsm_output[2]);
  assign nor_196_nl = ~((fsm_output[0]) | (~ and_tmp_9));
  assign mux_166_nl = MUX_s_1_2_2(nor_196_nl, and_tmp_9, or_tmp_133);
  assign and_706_nl = or_tmp_133 & ((fsm_output[0]) | Gelu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
      | Gelu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs);
  assign mux_167_nl = MUX_s_1_2_2(mux_166_nl, and_706_nl, fsm_output[1]);
  assign mux_168_nl = MUX_s_1_2_2(mux_167_nl, or_tmp_237, fsm_output[2]);
  assign mux_172_nl = MUX_s_1_2_2(mux_171_nl, mux_168_nl, fsm_output[3]);
  assign or_526_nl = Gelu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
      | Gelu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs;
  assign mux_176_nl = MUX_s_1_2_2(mux_175_nl, (~ mux_172_nl), or_526_nl);
  assign mux_178_nl = MUX_s_1_2_2(nor_198_nl, mux_176_nl, act_config_in_InstFetch_return_sva_7_2[4]);
  assign mux_179_nl = MUX_s_1_2_2(nor_197_nl, mux_178_nl, and_1103_cse);
  assign and_713_rmff = mux_179_nl & and_dcpl_587;
  assign and_719_rmff = and_dcpl_668 & and_dcpl_620 & (~ Tanh_for_2_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)
      & (~ Tanh_for_2_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs)
      & (fsm_output[4:3]==2'b01);
  assign and_724_rmff = and_dcpl_668 & and_dcpl_620 & (~ Tanh_for_3_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs)
      & (~ Tanh_for_3_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)
      & (fsm_output[4:3]==2'b01);
  assign and_729_rmff = and_dcpl_668 & and_dcpl_620 & (~ Tanh_for_4_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs)
      & (~ Tanh_for_4_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)
      & (fsm_output[4:3]==2'b01);
  assign and_734_rmff = and_dcpl_668 & and_dcpl_620 & (~ Tanh_for_5_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs)
      & (~ Tanh_for_5_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)
      & (fsm_output[4:3]==2'b01);
  assign and_739_rmff = and_dcpl_668 & and_dcpl_620 & (~ Tanh_for_6_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs)
      & (~ Tanh_for_6_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)
      & (fsm_output[4:3]==2'b01);
  assign and_744_rmff = and_dcpl_668 & and_dcpl_620 & (~ Tanh_for_7_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs)
      & (~ Tanh_for_7_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)
      & (fsm_output[4:3]==2'b01);
  assign and_749_rmff = and_dcpl_668 & and_dcpl_620 & (~ Tanh_for_8_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs)
      & (~ Tanh_for_8_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)
      & (fsm_output[4:3]==2'b01);
  assign and_754_rmff = and_dcpl_668 & and_dcpl_620 & (~ Tanh_for_9_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs)
      & (~ Tanh_for_9_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)
      & (fsm_output[4:3]==2'b01);
  assign and_759_rmff = and_dcpl_668 & and_dcpl_620 & (~ Tanh_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs)
      & (~ Tanh_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)
      & (fsm_output[4:3]==2'b01);
  assign and_764_rmff = and_dcpl_668 & and_dcpl_620 & (~ Tanh_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs)
      & (~ Tanh_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)
      & (fsm_output[4:3]==2'b01);
  assign and_769_rmff = and_dcpl_668 & and_dcpl_620 & (~ Tanh_for_12_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs)
      & (~ Tanh_for_12_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)
      & (fsm_output[4:3]==2'b01);
  assign and_774_rmff = and_dcpl_668 & and_dcpl_620 & (~ Tanh_for_13_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs)
      & (~ Tanh_for_13_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)
      & (fsm_output[4:3]==2'b01);
  assign and_779_rmff = and_dcpl_668 & and_dcpl_620 & (~ Tanh_for_14_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs)
      & (~ Tanh_for_14_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)
      & (fsm_output[4:3]==2'b01);
  assign and_784_rmff = and_dcpl_668 & and_dcpl_620 & (~ Tanh_for_15_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs)
      & (~ Tanh_for_15_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)
      & (fsm_output[4:3]==2'b01);
  assign and_789_rmff = and_dcpl_668 & and_dcpl_620 & (~ Tanh_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs)
      & (~ Tanh_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)
      & (fsm_output[4:3]==2'b01);
  assign and_794_rmff = and_dcpl_668 & and_dcpl_620 & (~ Tanh_for_1_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs)
      & (~ Tanh_for_1_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)
      & (fsm_output[4:3]==2'b01);
  assign nor_199_nl = ~(operator_32_8_true_AC_TRN_AC_WRAP_2_less_12_tmp_1 | operator_32_8_true_AC_TRN_AC_WRAP_3_less_12_tmp
      | (~ (act_config_in_InstFetch_mux_tmp[4])) | (act_config_in_InstFetch_mux_tmp[6])
      | nand_181_cse);
  assign nor_200_nl = ~(Tanh_for_4_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | Tanh_for_4_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
      | (~ (act_config_in_InstFetch_return_sva_7_2[2])) | (act_config_in_InstFetch_return_sva_7_2[4])
      | not_tmp_311);
  assign mux_180_nl = MUX_s_1_2_2(nor_199_nl, nor_200_nl, fsm_output[1]);
  assign and_799_rmff = mux_180_nl & and_dcpl_748;
  assign nor_201_nl = ~(operator_32_8_true_AC_TRN_AC_WRAP_2_less_11_tmp_1 | operator_32_8_true_AC_TRN_AC_WRAP_3_less_11_tmp
      | (~ (act_config_in_InstFetch_mux_tmp[4])) | (act_config_in_InstFetch_mux_tmp[6])
      | nand_181_cse);
  assign nor_202_nl = ~(Tanh_for_5_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | Tanh_for_5_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
      | (~ (act_config_in_InstFetch_return_sva_7_2[2])) | (act_config_in_InstFetch_return_sva_7_2[4])
      | not_tmp_311);
  assign mux_181_nl = MUX_s_1_2_2(nor_201_nl, nor_202_nl, fsm_output[1]);
  assign and_800_rmff = mux_181_nl & and_dcpl_748;
  assign nor_203_nl = ~(operator_32_8_true_AC_TRN_AC_WRAP_2_less_10_tmp_1 | operator_32_8_true_AC_TRN_AC_WRAP_3_less_10_tmp
      | (~ (act_config_in_InstFetch_mux_tmp[4])) | (act_config_in_InstFetch_mux_tmp[6])
      | nand_181_cse);
  assign nor_204_nl = ~(Tanh_for_6_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | Tanh_for_6_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
      | (~ (act_config_in_InstFetch_return_sva_7_2[2])) | (act_config_in_InstFetch_return_sva_7_2[4])
      | not_tmp_311);
  assign mux_182_nl = MUX_s_1_2_2(nor_203_nl, nor_204_nl, fsm_output[1]);
  assign and_801_rmff = mux_182_nl & and_dcpl_748;
  assign nor_205_nl = ~(operator_32_8_true_AC_TRN_AC_WRAP_2_less_9_tmp_1 | operator_32_8_true_AC_TRN_AC_WRAP_3_less_9_tmp
      | (~ (act_config_in_InstFetch_mux_tmp[4])) | (act_config_in_InstFetch_mux_tmp[6])
      | nand_181_cse);
  assign nor_206_nl = ~(Tanh_for_7_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | Tanh_for_7_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
      | (~ (act_config_in_InstFetch_return_sva_7_2[2])) | (act_config_in_InstFetch_return_sva_7_2[4])
      | not_tmp_311);
  assign mux_183_nl = MUX_s_1_2_2(nor_205_nl, nor_206_nl, fsm_output[1]);
  assign and_802_rmff = mux_183_nl & and_dcpl_748;
  assign nor_207_nl = ~((~ (act_config_in_InstFetch_mux_tmp[4])) | (act_config_in_InstFetch_mux_tmp[6])
      | operator_32_8_true_AC_TRN_AC_WRAP_2_less_8_tmp_1 | operator_32_8_true_AC_TRN_AC_WRAP_3_less_8_tmp
      | nand_181_cse);
  assign nor_208_nl = ~(Tanh_for_8_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | Tanh_for_8_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
      | (~ (act_config_in_InstFetch_return_sva_7_2[2])) | (act_config_in_InstFetch_return_sva_7_2[4])
      | not_tmp_311);
  assign mux_184_nl = MUX_s_1_2_2(nor_207_nl, nor_208_nl, fsm_output[1]);
  assign and_803_rmff = mux_184_nl & and_dcpl_748;
  assign nor_209_nl = ~(operator_32_8_true_AC_TRN_AC_WRAP_2_less_7_tmp_1 | operator_32_8_true_AC_TRN_AC_WRAP_3_less_7_tmp
      | (~ (act_config_in_InstFetch_mux_tmp[4])) | (act_config_in_InstFetch_mux_tmp[6])
      | nand_181_cse);
  assign nor_210_nl = ~(Tanh_for_9_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | Tanh_for_9_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
      | (~ (act_config_in_InstFetch_return_sva_7_2[2])) | (act_config_in_InstFetch_return_sva_7_2[4])
      | not_tmp_311);
  assign mux_185_nl = MUX_s_1_2_2(nor_209_nl, nor_210_nl, fsm_output[1]);
  assign and_804_rmff = mux_185_nl & and_dcpl_748;
  assign nor_211_nl = ~(operator_32_8_true_AC_TRN_AC_WRAP_2_less_6_tmp_1 | operator_32_8_true_AC_TRN_AC_WRAP_3_less_6_tmp
      | (~ (act_config_in_InstFetch_mux_tmp[4])) | (act_config_in_InstFetch_mux_tmp[6])
      | nand_181_cse);
  assign nor_212_nl = ~(Tanh_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | Tanh_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
      | (~ (act_config_in_InstFetch_return_sva_7_2[2])) | (act_config_in_InstFetch_return_sva_7_2[4])
      | not_tmp_311);
  assign mux_186_nl = MUX_s_1_2_2(nor_211_nl, nor_212_nl, fsm_output[1]);
  assign and_805_rmff = mux_186_nl & and_dcpl_748;
  assign nor_213_nl = ~(operator_32_8_true_AC_TRN_AC_WRAP_2_less_5_tmp_1 | operator_32_8_true_AC_TRN_AC_WRAP_3_less_5_tmp
      | (~ (act_config_in_InstFetch_mux_tmp[4])) | (act_config_in_InstFetch_mux_tmp[6])
      | nand_181_cse);
  assign nor_214_nl = ~(Tanh_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | Tanh_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
      | (~ (act_config_in_InstFetch_return_sva_7_2[2])) | (act_config_in_InstFetch_return_sva_7_2[4])
      | not_tmp_311);
  assign mux_187_nl = MUX_s_1_2_2(nor_213_nl, nor_214_nl, fsm_output[1]);
  assign and_806_rmff = mux_187_nl & and_dcpl_748;
  assign nor_215_nl = ~(operator_32_8_true_AC_TRN_AC_WRAP_2_less_4_tmp_1 | operator_32_8_true_AC_TRN_AC_WRAP_3_less_4_tmp
      | (~ (act_config_in_InstFetch_mux_tmp[4])) | (act_config_in_InstFetch_mux_tmp[6])
      | nand_181_cse);
  assign nor_216_nl = ~(Tanh_for_12_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | Tanh_for_12_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
      | (~ (act_config_in_InstFetch_return_sva_7_2[2])) | (act_config_in_InstFetch_return_sva_7_2[4])
      | not_tmp_311);
  assign mux_188_nl = MUX_s_1_2_2(nor_215_nl, nor_216_nl, fsm_output[1]);
  assign and_807_rmff = mux_188_nl & and_dcpl_748;
  assign nor_217_nl = ~(operator_32_8_true_AC_TRN_AC_WRAP_2_less_3_tmp_1 | operator_32_8_true_AC_TRN_AC_WRAP_3_less_3_tmp
      | (~ (act_config_in_InstFetch_mux_tmp[4])) | (act_config_in_InstFetch_mux_tmp[6])
      | nand_181_cse);
  assign nor_218_nl = ~(Tanh_for_13_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | Tanh_for_13_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
      | (~ (act_config_in_InstFetch_return_sva_7_2[2])) | (act_config_in_InstFetch_return_sva_7_2[4])
      | not_tmp_311);
  assign mux_189_nl = MUX_s_1_2_2(nor_217_nl, nor_218_nl, fsm_output[1]);
  assign and_808_rmff = mux_189_nl & and_dcpl_748;
  assign nor_219_nl = ~(operator_32_8_true_AC_TRN_AC_WRAP_2_less_2_tmp_1 | operator_32_8_true_AC_TRN_AC_WRAP_3_less_2_tmp
      | (~ (act_config_in_InstFetch_mux_tmp[4])) | (act_config_in_InstFetch_mux_tmp[6])
      | nand_181_cse);
  assign nor_220_nl = ~(Tanh_for_14_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | Tanh_for_14_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
      | (~ (act_config_in_InstFetch_return_sva_7_2[2])) | (act_config_in_InstFetch_return_sva_7_2[4])
      | not_tmp_311);
  assign mux_190_nl = MUX_s_1_2_2(nor_219_nl, nor_220_nl, fsm_output[1]);
  assign and_809_rmff = mux_190_nl & and_dcpl_748;
  assign nor_221_nl = ~(operator_32_8_true_AC_TRN_AC_WRAP_2_less_1_tmp_1 | operator_32_8_true_AC_TRN_AC_WRAP_3_less_1_tmp
      | (~ (act_config_in_InstFetch_mux_tmp[4])) | (act_config_in_InstFetch_mux_tmp[6])
      | nand_181_cse);
  assign nor_222_nl = ~(Tanh_for_15_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | Tanh_for_15_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
      | (~ (act_config_in_InstFetch_return_sva_7_2[2])) | (act_config_in_InstFetch_return_sva_7_2[4])
      | not_tmp_311);
  assign mux_191_nl = MUX_s_1_2_2(nor_221_nl, nor_222_nl, fsm_output[1]);
  assign and_810_rmff = mux_191_nl & and_dcpl_748;
  assign nor_223_nl = ~(operator_32_8_true_AC_TRN_AC_WRAP_2_less_tmp_1 | operator_32_8_true_AC_TRN_AC_WRAP_3_less_tmp
      | (~ (act_config_in_InstFetch_mux_tmp[4])) | (act_config_in_InstFetch_mux_tmp[6])
      | nand_181_cse);
  assign nor_224_nl = ~(Tanh_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | Tanh_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
      | (~ (act_config_in_InstFetch_return_sva_7_2[2])) | (act_config_in_InstFetch_return_sva_7_2[4])
      | not_tmp_311);
  assign mux_192_nl = MUX_s_1_2_2(nor_223_nl, nor_224_nl, fsm_output[1]);
  assign and_811_rmff = mux_192_nl & and_dcpl_748;
  assign nor_225_nl = ~(operator_32_8_true_AC_TRN_AC_WRAP_2_less_13_tmp_1 | operator_32_8_true_AC_TRN_AC_WRAP_3_less_13_tmp
      | (~ (act_config_in_InstFetch_mux_tmp[4])) | (act_config_in_InstFetch_mux_tmp[6])
      | nand_181_cse);
  assign nor_226_nl = ~(Tanh_for_3_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | Tanh_for_3_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
      | (~ (act_config_in_InstFetch_return_sva_7_2[2])) | (act_config_in_InstFetch_return_sva_7_2[4])
      | not_tmp_311);
  assign mux_193_nl = MUX_s_1_2_2(nor_225_nl, nor_226_nl, fsm_output[1]);
  assign and_812_rmff = mux_193_nl & and_dcpl_748;
  assign and_819_rmff = and_dcpl_768 & is_incr_lpi_1_dfm_1 & (operator_6_false_acc_tmp[6:5]==2'b00)
      & act_config_InstIncr_if_equal_1_tmp & act_config_InstIncr_if_act_config_InstIncr_if_if_nor_tmp;
  assign and_823_rmff = and_dcpl_377 & and_dcpl_770 & and_dcpl_559;
  assign and_826_rmff = and_dcpl_775 & and_dcpl_564;
  assign and_830_rmff = and_dcpl_774 & (fsm_output[2]) & (~ (fsm_output[0])) & nor_57_cse
      & w_axi_rsp_lpi_1_dfm_1;
  assign and_835_rmff = is_start_sva & (act_config_in_InstFetch_mux_tmp[7:4]==4'b0011)
      & and_dcpl_554;
  assign and_837_rmff = and_dcpl_786 & and_dcpl_568;
  assign nor_62_nl = ~((~ (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[0])) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[8]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[9]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[10]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3]));
  assign or_172_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[0]) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[8]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[9]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[10]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3]);
  assign mux_52_nl = MUX_s_1_2_2(nor_62_nl, or_172_nl, act_config_is_valid_sva);
  assign nor_18_nl = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1:0]!=2'b01));
  assign mux_53_nl = MUX_s_1_2_2(act_config_is_valid_sva, mux_52_nl, nor_18_nl);
  assign ActUnit_DecodeAxi_if_and_37_cse = ActUnitRun_wen & and_dcpl_788 & (mux_53_nl
      | is_start_sva);
  assign nor_74_nl = ~(ActUnit_CheckStart_if_ActUnit_CheckStart_if_and_itm_1 | is_start_sva);
  assign or_242_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | act_config_is_zero_first_sva
      | (~ and_dcpl_370);
  assign or_240_nl = act_config_is_zero_first_sva | (~ and_dcpl_370);
  assign nor_347_nl = ~(is_start_sva | act_config_is_valid_sva);
  assign mux_75_nl = MUX_s_1_2_2(or_tmp_111, nor_347_nl, w_load_lpi_1_dfm_1);
  assign mux_76_nl = MUX_s_1_2_2(mux_75_nl, or_tmp_111, act_config_is_zero_first_sva);
  assign mux_77_nl = MUX_s_1_2_2(or_240_nl, mux_76_nl, ActUnit_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva);
  assign or_238_nl = (~ ActUnit_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva)
      | (~ act_config_is_valid_sva) | is_start_sva;
  assign mux_78_nl = MUX_s_1_2_2(mux_77_nl, or_238_nl, ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]);
  assign mux_79_nl = MUX_s_1_2_2(or_242_nl, mux_78_nl, ActUnit_CheckStart_start_reg_sva);
  assign mux_80_nl = MUX_s_1_2_2(nor_74_nl, mux_79_nl, is_incr_lpi_1_dfm_1);
  assign act_config_inst_regs_and_36_cse = ActUnitRun_wen & and_dcpl_799 & mux_80_nl;
  assign act_config_num_inst_and_cse = ActUnitRun_wen & (~(or_dcpl_320 | or_dcpl_310
      | or_dcpl_296 | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1:0]!=2'b01)));
  assign rva_out_reg_data_and_cse = ActUnitRun_wen & (and_dcpl_803 | and_dcpl_805);
  assign act_mem_banks_bank_a_and_cse = ActUnitRun_wen & (~(or_dcpl_335 | or_dcpl_333
      | or_dcpl_330));
  assign act_mem_banks_bank_a_and_1_cse = ActUnitRun_wen & (~(or_dcpl_335 | or_dcpl_338
      | or_dcpl_330));
  assign act_mem_banks_bank_a_and_2_cse = ActUnitRun_wen & (~(or_dcpl_335 | or_dcpl_333
      | or_dcpl_342));
  assign act_mem_banks_bank_a_and_3_cse = ActUnitRun_wen & (~(or_dcpl_335 | or_dcpl_338
      | or_dcpl_342));
  assign act_mem_banks_bank_a_and_4_cse = ActUnitRun_wen & (~(or_dcpl_335 | or_dcpl_333
      | or_dcpl_348));
  assign act_mem_banks_bank_a_and_5_cse = ActUnitRun_wen & (~(or_dcpl_335 | or_dcpl_338
      | or_dcpl_348));
  assign act_mem_banks_bank_a_and_6_cse = ActUnitRun_wen & (~(or_dcpl_335 | or_dcpl_333
      | or_dcpl_353));
  assign act_mem_banks_bank_a_and_7_cse = ActUnitRun_wen & (~(or_dcpl_335 | or_dcpl_338
      | or_dcpl_353));
  assign act_mem_banks_bank_a_and_8_cse = ActUnitRun_wen & (~(or_dcpl_335 | or_dcpl_333
      | or_dcpl_359));
  assign act_mem_banks_bank_a_and_9_cse = ActUnitRun_wen & (~(or_dcpl_335 | or_dcpl_338
      | or_dcpl_359));
  assign act_mem_banks_bank_a_and_10_cse = ActUnitRun_wen & (~(or_dcpl_335 | or_dcpl_333
      | or_dcpl_364));
  assign act_mem_banks_bank_a_and_11_cse = ActUnitRun_wen & (~(or_dcpl_335 | or_dcpl_338
      | or_dcpl_364));
  assign act_mem_banks_bank_a_and_12_cse = ActUnitRun_wen & (~(or_dcpl_335 | or_dcpl_333
      | or_dcpl_370));
  assign act_mem_banks_bank_a_and_13_cse = ActUnitRun_wen & (~(or_dcpl_335 | or_dcpl_338
      | or_dcpl_370));
  assign act_mem_banks_bank_a_and_14_cse = ActUnitRun_wen & (~(or_dcpl_335 | or_dcpl_333
      | or_dcpl_375));
  assign act_mem_banks_bank_a_and_15_cse = ActUnitRun_wen & (~(or_dcpl_335 | or_dcpl_338
      | or_dcpl_375));
  assign act_mem_banks_bank_a_and_16_cse = ActUnitRun_wen & (~(or_dcpl_335 | or_dcpl_333
      | or_dcpl_381));
  assign act_mem_banks_bank_a_and_17_cse = ActUnitRun_wen & (~(or_dcpl_335 | or_dcpl_338
      | or_dcpl_381));
  assign act_mem_banks_bank_a_and_18_cse = ActUnitRun_wen & (~(or_dcpl_335 | or_dcpl_333
      | or_dcpl_387));
  assign act_mem_banks_bank_a_and_19_cse = ActUnitRun_wen & (~(or_dcpl_335 | or_dcpl_338
      | or_dcpl_387));
  assign act_mem_banks_bank_a_and_20_cse = ActUnitRun_wen & (~(or_dcpl_335 | or_dcpl_333
      | or_dcpl_392));
  assign act_mem_banks_bank_a_and_21_cse = ActUnitRun_wen & (~(or_dcpl_335 | or_dcpl_338
      | or_dcpl_392));
  assign act_mem_banks_bank_a_and_22_cse = ActUnitRun_wen & (~(or_dcpl_335 | or_dcpl_333
      | or_dcpl_397));
  assign act_mem_banks_bank_a_and_23_cse = ActUnitRun_wen & (~(or_dcpl_335 | or_dcpl_338
      | or_dcpl_397));
  assign act_mem_banks_bank_a_and_24_cse = ActUnitRun_wen & (~(or_dcpl_335 | or_dcpl_333
      | or_dcpl_402));
  assign act_mem_banks_bank_a_and_25_cse = ActUnitRun_wen & (~(or_dcpl_335 | or_dcpl_338
      | or_dcpl_402));
  assign act_mem_banks_bank_a_and_26_cse = ActUnitRun_wen & (~(or_dcpl_335 | or_dcpl_333
      | or_dcpl_407));
  assign act_mem_banks_bank_a_and_27_cse = ActUnitRun_wen & (~(or_dcpl_335 | or_dcpl_338
      | or_dcpl_407));
  assign act_mem_banks_bank_a_and_28_cse = ActUnitRun_wen & (~(or_dcpl_335 | or_dcpl_333
      | or_dcpl_412));
  assign act_mem_banks_bank_a_and_29_cse = ActUnitRun_wen & (~(or_dcpl_335 | or_dcpl_338
      | or_dcpl_412));
  assign act_mem_banks_bank_a_and_30_cse = ActUnitRun_wen & (~(or_dcpl_335 | or_dcpl_333
      | or_dcpl_417));
  assign act_mem_banks_bank_a_and_31_cse = ActUnitRun_wen & (~(or_dcpl_335 | or_dcpl_338
      | or_dcpl_417));
  assign act_config_inst_regs_and_4_cse = ActUnitRun_wen & (~(or_dcpl_423 | or_dcpl_322
      | not_tmp_347));
  assign act_config_inst_regs_and_20_cse = ActUnitRun_wen & (~(or_dcpl_320 | or_dcpl_310
      | or_dcpl_296 | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1:0]!=2'b10)));
  assign act_regs_data_and_cse = ActUnitRun_wen & and_dcpl_814;
  assign act_regs_data_and_859_enex5 = act_regs_data_and_cse & (reg_w_load_lpi_1_dfm_1_enexo
      | reg_is_start_enexo | reg_act_regs_data_2_2_3_enexo | reg_act_config_is_zero_first_sva_dfm_4_enexo
      | reg_act_regs_data_3_15_sva_dfm_2_1_enexo | reg_act_regs_data_3_15_3_enexo);
  assign act_regs_data_and_860_enex5 = act_regs_data_and_cse & (reg_is_start_enexo_1
      | reg_act_regs_data_3_14_sva_dfm_2_1_enexo | reg_act_regs_data_3_14_3_enexo
      | reg_w_load_lpi_1_dfm_1_enexo_1 | reg_act_config_is_zero_first_sva_dfm_4_enexo_1
      | reg_act_regs_data_2_15_3_enexo);
  assign act_regs_data_and_861_enex5 = act_regs_data_and_cse & (reg_act_regs_data_3_13_3_enexo
      | reg_is_start_enexo_2 | reg_act_regs_data_2_14_3_enexo | reg_act_regs_data_3_13_sva_dfm_2_1_enexo
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_2 | reg_w_load_lpi_1_dfm_1_enexo_2);
  assign act_regs_data_and_862_enex5 = act_regs_data_and_cse & (reg_act_regs_data_3_12_3_enexo
      | reg_act_regs_data_2_13_3_enexo | reg_act_config_is_zero_first_sva_dfm_4_enexo_3
      | reg_w_load_lpi_1_dfm_1_enexo_3 | reg_is_start_enexo_3 | reg_act_regs_data_3_12_sva_dfm_2_1_enexo);
  assign act_regs_data_and_863_enex5 = act_regs_data_and_cse & (reg_w_load_lpi_1_dfm_1_enexo_4
      | reg_is_start_enexo_4 | reg_act_config_is_zero_first_sva_dfm_4_enexo_4 | reg_act_regs_data_2_12_3_enexo
      | reg_act_regs_data_3_11_sva_dfm_2_1_enexo | reg_act_regs_data_3_11_3_enexo);
  assign act_regs_data_and_864_enex5 = act_regs_data_and_cse & (reg_act_config_is_zero_first_sva_dfm_4_enexo_5
      | reg_w_load_lpi_1_dfm_1_enexo_5 | reg_is_start_enexo_5 | reg_act_regs_data_2_11_3_enexo
      | reg_act_regs_data_3_10_sva_dfm_2_1_enexo | reg_act_regs_data_3_10_3_enexo);
  assign act_regs_data_and_865_enex5 = act_regs_data_and_cse & (reg_act_regs_data_3_9_sva_dfm_2_1_enexo
      | reg_act_regs_data_3_9_3_enexo | reg_w_load_lpi_1_dfm_1_enexo_6 | reg_act_config_is_zero_first_sva_dfm_4_enexo_6
      | reg_is_start_enexo_6 | reg_act_regs_data_3_0_3_enexo);
  assign act_regs_data_and_866_enex5 = act_regs_data_and_cse & (reg_act_regs_data_2_9_3_enexo
      | reg_w_load_lpi_1_dfm_1_enexo_7 | reg_is_start_enexo_7 | reg_act_config_is_zero_first_sva_dfm_4_enexo_7
      | reg_act_regs_data_3_8_3_enexo | reg_act_regs_data_3_8_sva_dfm_2_1_enexo);
  assign act_regs_data_and_867_enex5 = act_regs_data_and_cse & (reg_act_regs_data_3_7_3_enexo
      | reg_w_load_lpi_1_dfm_1_enexo_8 | reg_act_regs_data_2_8_3_enexo | reg_act_regs_data_3_7_sva_dfm_2_1_enexo
      | reg_is_start_enexo_8 | reg_act_config_is_zero_first_sva_dfm_4_enexo_8);
  assign act_regs_data_and_868_enex5 = act_regs_data_and_cse & (reg_act_config_is_zero_first_sva_dfm_4_enexo_9
      | reg_act_regs_data_3_6_sva_dfm_2_1_enexo | reg_w_load_lpi_1_dfm_1_enexo_9
      | reg_act_regs_data_3_6_3_enexo | reg_act_regs_data_2_7_3_enexo | reg_is_start_enexo_9);
  assign act_regs_data_and_869_enex5 = act_regs_data_and_cse & (reg_act_regs_data_3_5_sva_dfm_2_1_enexo
      | reg_w_load_lpi_1_dfm_1_enexo_10 | reg_is_start_enexo_10 | reg_act_config_is_zero_first_sva_dfm_4_enexo_10
      | reg_act_regs_data_3_5_3_enexo | reg_act_regs_data_2_6_3_enexo);
  assign act_regs_data_and_870_enex5 = act_regs_data_and_cse & (reg_is_start_enexo_11
      | reg_act_regs_data_3_4_3_enexo | reg_w_load_lpi_1_dfm_1_enexo_11 | reg_act_config_is_zero_first_sva_dfm_4_enexo_11
      | reg_act_regs_data_2_5_3_enexo | reg_act_regs_data_3_4_sva_dfm_2_1_enexo);
  assign act_regs_data_and_871_enex5 = act_regs_data_and_cse & (reg_act_regs_data_3_3_sva_dfm_2_1_enexo
      | reg_is_start_enexo_12 | reg_act_regs_data_2_4_3_enexo | reg_act_config_is_zero_first_sva_dfm_4_enexo_12
      | reg_w_load_lpi_1_dfm_1_enexo_12 | reg_act_regs_data_3_3_3_enexo);
  assign act_regs_data_and_872_enex5 = act_regs_data_and_cse & (reg_act_regs_data_3_2_sva_dfm_2_1_enexo
      | reg_act_regs_data_3_2_3_enexo | reg_w_load_lpi_1_dfm_1_enexo_13 | reg_is_start_enexo_13
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_13 | reg_act_regs_data_2_3_3_enexo);
  assign act_regs_data_and_873_enex5 = act_regs_data_and_cse & (reg_act_regs_data_2_10_3_enexo
      | reg_is_start_enexo_14 | reg_w_load_lpi_1_dfm_1_enexo_14 | reg_act_config_is_zero_first_sva_dfm_4_enexo_14
      | reg_act_regs_data_3_1_3_enexo | reg_act_regs_data_3_1_sva_dfm_2_1_enexo);
  assign act_regs_data_and_874_enex5 = act_regs_data_and_cse & (reg_act_regs_data_3_0_sva_dfm_2_1_enexo
      | reg_is_start_enexo_15 | reg_act_regs_data_2_1_3_enexo | reg_act_regs_data_3_0_3_enexo_1
      | reg_w_load_lpi_1_dfm_1_enexo_15 | reg_act_config_is_zero_first_sva_dfm_4_enexo_15);
  assign act_regs_data_and_875_enex5 = act_regs_data_and_cse & (reg_act_regs_data_2_15_sva_dfm_2_1_enexo
      | reg_w_load_lpi_1_dfm_1_enexo_16 | reg_act_regs_data_1_2_3_enexo | reg_act_regs_data_2_15_3_enexo_1
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_16 | reg_is_start_enexo_16);
  assign act_regs_data_and_876_enex5 = act_regs_data_and_cse & (reg_act_config_is_zero_first_sva_dfm_4_enexo_17
      | reg_act_regs_data_1_15_3_enexo | reg_act_regs_data_2_14_3_enexo_1 | reg_is_start_enexo_17
      | reg_w_load_lpi_1_dfm_1_enexo_17 | reg_act_regs_data_2_14_sva_dfm_2_1_enexo);
  assign act_regs_data_and_877_enex5 = act_regs_data_and_cse & (reg_act_regs_data_2_13_sva_dfm_2_1_enexo
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_18 | reg_act_regs_data_2_13_3_enexo_1
      | reg_act_regs_data_1_14_3_enexo | reg_w_load_lpi_1_dfm_1_enexo_18 | reg_is_start_enexo_18);
  assign act_regs_data_and_878_enex5 = act_regs_data_and_cse & (reg_act_regs_data_2_12_sva_dfm_2_1_enexo
      | reg_act_regs_data_1_13_3_enexo | reg_act_config_is_zero_first_sva_dfm_4_enexo_19
      | reg_act_regs_data_2_12_3_enexo_1 | reg_is_start_enexo_19 | reg_w_load_lpi_1_dfm_1_enexo_19);
  assign act_regs_data_and_879_enex5 = act_regs_data_and_cse & (reg_act_config_is_zero_first_sva_dfm_4_enexo_20
      | reg_is_start_enexo_20 | reg_act_regs_data_2_11_3_enexo_1 | reg_w_load_lpi_1_dfm_1_enexo_20
      | reg_act_regs_data_2_11_sva_dfm_2_1_enexo | reg_act_regs_data_1_12_3_enexo);
  assign act_regs_data_and_880_enex5 = act_regs_data_and_cse & (reg_act_regs_data_1_11_3_enexo
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_21 | reg_w_load_lpi_1_dfm_1_enexo_21
      | reg_is_start_enexo_21 | reg_act_regs_data_2_10_sva_dfm_2_1_enexo | reg_act_regs_data_2_10_3_enexo_1);
  assign act_regs_data_and_881_enex5 = act_regs_data_and_cse & (reg_act_config_is_zero_first_sva_dfm_4_enexo_22
      | reg_act_regs_data_2_9_3_enexo_1 | reg_act_regs_data_2_0_3_enexo | reg_is_start_enexo_22
      | reg_w_load_lpi_1_dfm_1_enexo_22 | reg_act_regs_data_2_9_sva_dfm_2_1_enexo);
  assign act_regs_data_and_882_enex5 = act_regs_data_and_cse & (reg_act_regs_data_2_8_sva_dfm_2_1_enexo
      | reg_is_start_enexo_23 | reg_act_regs_data_2_8_3_enexo_1 | reg_act_config_is_zero_first_sva_dfm_4_enexo_23
      | reg_act_regs_data_1_9_3_enexo | reg_w_load_lpi_1_dfm_1_enexo_23);
  assign act_regs_data_and_883_enex5 = act_regs_data_and_cse & (reg_act_regs_data_1_8_3_enexo
      | reg_act_regs_data_2_7_3_enexo_1 | reg_act_config_is_zero_first_sva_dfm_4_enexo_24
      | reg_w_load_lpi_1_dfm_1_enexo_24 | reg_act_regs_data_2_7_sva_dfm_2_1_enexo
      | reg_is_start_enexo_24);
  assign act_regs_data_and_884_enex5 = act_regs_data_and_cse & (reg_act_regs_data_2_6_3_enexo_1
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_25 | reg_w_load_lpi_1_dfm_1_enexo_25
      | reg_act_regs_data_1_7_3_enexo | reg_act_regs_data_2_6_sva_dfm_2_1_enexo |
      reg_is_start_enexo_25);
  assign act_regs_data_and_885_enex5 = act_regs_data_and_cse & (reg_act_regs_data_1_6_3_enexo
      | reg_w_load_lpi_1_dfm_1_enexo_26 | reg_is_start_enexo_26 | reg_act_config_is_zero_first_sva_dfm_4_enexo_26
      | reg_act_regs_data_2_5_3_enexo_1 | reg_act_regs_data_2_5_sva_dfm_2_1_enexo);
  assign act_regs_data_and_886_enex5 = act_regs_data_and_cse & (reg_act_config_is_zero_first_sva_dfm_4_enexo_27
      | reg_is_start_enexo_27 | reg_act_regs_data_1_5_3_enexo | reg_act_regs_data_2_4_3_enexo_1
      | reg_act_regs_data_2_4_sva_dfm_2_1_enexo | reg_w_load_lpi_1_dfm_1_enexo_27);
  assign act_regs_data_and_887_enex5 = act_regs_data_and_cse & (reg_act_regs_data_2_3_sva_dfm_2_1_enexo
      | reg_act_regs_data_2_3_3_enexo_1 | reg_is_start_enexo_28 | reg_w_load_lpi_1_dfm_1_enexo_28
      | reg_act_regs_data_1_4_3_enexo | reg_act_config_is_zero_first_sva_dfm_4_enexo_28);
  assign act_regs_data_and_888_enex5 = act_regs_data_and_cse & (reg_act_regs_data_2_2_sva_dfm_2_1_enexo
      | reg_is_start_enexo_29 | reg_act_config_is_zero_first_sva_dfm_4_enexo_29 |
      reg_w_load_lpi_1_dfm_1_enexo_29 | reg_act_regs_data_2_2_3_enexo_1 | reg_act_regs_data_1_3_3_enexo);
  assign act_regs_data_and_889_enex5 = act_regs_data_and_cse & (reg_act_config_is_zero_first_sva_dfm_4_enexo_30
      | reg_w_load_lpi_1_dfm_1_enexo_30 | reg_act_regs_data_1_10_3_enexo | reg_act_regs_data_2_1_sva_dfm_2_1_enexo
      | reg_act_regs_data_2_1_3_enexo_1 | reg_is_start_enexo_30);
  assign act_regs_data_and_890_enex5 = act_regs_data_and_cse & (reg_act_regs_data_2_0_sva_dfm_2_1_enexo
      | reg_is_start_enexo_31 | reg_act_regs_data_1_1_3_enexo | reg_w_load_lpi_1_dfm_1_enexo_31
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_31 | reg_act_regs_data_2_0_3_enexo_1);
  assign act_regs_data_and_891_enex5 = act_regs_data_and_cse & (reg_act_regs_data_0_2_3_enexo
      | reg_is_start_enexo_32 | reg_act_regs_data_1_15_sva_dfm_2_1_enexo | reg_w_load_lpi_1_dfm_1_enexo_32
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_32 | reg_act_regs_data_1_15_3_enexo_1);
  assign act_regs_data_and_892_enex5 = act_regs_data_and_cse & (reg_act_regs_data_0_15_3_enexo
      | reg_act_regs_data_1_14_3_enexo_1 | reg_act_config_is_zero_first_sva_dfm_4_enexo_33
      | reg_act_regs_data_1_14_sva_dfm_2_1_enexo | reg_w_load_lpi_1_dfm_1_enexo_33
      | reg_is_start_enexo_33);
  assign act_regs_data_and_893_enex5 = act_regs_data_and_cse & (reg_act_regs_data_1_13_sva_dfm_2_1_enexo
      | reg_w_load_lpi_1_dfm_1_enexo_34 | reg_act_regs_data_0_14_3_enexo | reg_act_regs_data_1_13_3_enexo_1
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_34 | reg_is_start_enexo_34);
  assign act_regs_data_and_894_enex5 = act_regs_data_and_cse & (reg_act_regs_data_1_12_sva_dfm_2_1_enexo
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_35 | reg_act_regs_data_0_13_3_enexo
      | reg_is_start_enexo_35 | reg_act_regs_data_1_12_3_enexo_1 | reg_w_load_lpi_1_dfm_1_enexo_35);
  assign act_regs_data_and_895_enex5 = act_regs_data_and_cse & (reg_act_regs_data_1_11_sva_dfm_2_1_enexo
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_36 | reg_act_regs_data_0_12_3_enexo
      | reg_w_load_lpi_1_dfm_1_enexo_36 | reg_is_start_enexo_36 | reg_act_regs_data_1_11_3_enexo_1);
  assign act_regs_data_and_896_enex5 = act_regs_data_and_cse & (reg_act_regs_data_1_10_3_enexo_1
      | reg_w_load_lpi_1_dfm_1_enexo_37 | reg_act_regs_data_0_11_3_enexo | reg_act_config_is_zero_first_sva_dfm_4_enexo_37
      | reg_is_start_enexo_37 | reg_act_regs_data_1_10_sva_dfm_2_1_enexo);
  assign act_regs_data_and_897_enex5 = act_regs_data_and_cse & (reg_is_start_enexo_38
      | reg_act_regs_data_1_0_3_enexo | reg_act_regs_data_1_9_sva_dfm_2_1_enexo |
      reg_act_regs_data_1_9_3_enexo_1 | reg_act_config_is_zero_first_sva_dfm_4_enexo_38
      | reg_w_load_lpi_1_dfm_1_enexo_38);
  assign act_regs_data_and_898_enex5 = act_regs_data_and_cse & (reg_act_config_is_zero_first_sva_dfm_4_enexo_39
      | reg_act_regs_data_1_8_3_enexo_1 | reg_act_regs_data_1_8_sva_dfm_2_1_enexo
      | reg_w_load_lpi_1_dfm_1_enexo_39 | reg_act_regs_data_0_9_3_enexo | reg_is_start_enexo_39);
  assign act_regs_data_and_899_enex5 = act_regs_data_and_cse & (reg_is_start_enexo_40
      | reg_act_regs_data_0_8_3_enexo | reg_act_regs_data_1_7_sva_dfm_2_1_enexo |
      reg_act_config_is_zero_first_sva_dfm_4_enexo_40 | reg_act_regs_data_1_7_3_enexo_1
      | reg_w_load_lpi_1_dfm_1_enexo_40);
  assign act_regs_data_and_900_enex5 = act_regs_data_and_cse & (reg_is_start_enexo_41
      | reg_act_regs_data_1_6_3_enexo_1 | reg_act_config_is_zero_first_sva_dfm_4_enexo_41
      | reg_w_load_lpi_1_dfm_1_enexo_41 | reg_act_regs_data_1_6_sva_dfm_2_1_enexo
      | reg_act_regs_data_0_7_3_enexo);
  assign act_regs_data_and_901_enex5 = act_regs_data_and_cse & (reg_act_config_is_zero_first_sva_dfm_4_enexo_42
      | reg_w_load_lpi_1_dfm_1_enexo_42 | reg_act_regs_data_1_5_sva_dfm_2_1_enexo
      | reg_act_regs_data_1_5_3_enexo_1 | reg_act_regs_data_0_6_3_enexo | reg_is_start_enexo_42);
  assign act_regs_data_and_902_enex5 = act_regs_data_and_cse & (reg_is_start_enexo_43
      | reg_act_regs_data_0_5_3_enexo | reg_act_regs_data_1_4_3_enexo_1 | reg_w_load_lpi_1_dfm_1_enexo_43
      | reg_act_regs_data_1_4_sva_dfm_2_1_enexo | reg_act_config_is_zero_first_sva_dfm_4_enexo_43);
  assign act_regs_data_and_903_enex5 = act_regs_data_and_cse & (reg_w_load_lpi_1_dfm_1_enexo_44
      | reg_act_regs_data_1_3_sva_dfm_2_1_enexo | reg_is_start_enexo_44 | reg_act_config_is_zero_first_sva_dfm_4_enexo_44
      | reg_act_regs_data_1_3_3_enexo_1 | reg_act_regs_data_0_4_3_enexo);
  assign act_regs_data_and_904_enex5 = act_regs_data_and_cse & (reg_act_regs_data_1_2_sva_dfm_2_1_enexo
      | reg_w_load_lpi_1_dfm_1_enexo_45 | reg_is_start_enexo_45 | reg_act_regs_data_1_2_3_enexo_1
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_45 | reg_act_regs_data_0_3_3_enexo);
  assign act_regs_data_and_905_enex5 = act_regs_data_and_cse & (reg_act_regs_data_1_1_3_enexo_1
      | reg_act_regs_data_0_10_3_enexo | reg_act_regs_data_1_1_sva_dfm_2_1_enexo
      | reg_is_start_enexo_46 | reg_act_config_is_zero_first_sva_dfm_4_enexo_46 |
      reg_w_load_lpi_1_dfm_1_enexo_46);
  assign act_regs_data_and_906_enex5 = act_regs_data_and_cse & (reg_is_start_enexo_47
      | reg_w_load_lpi_1_dfm_1_enexo_47 | reg_act_regs_data_0_1_3_enexo | reg_act_config_is_zero_first_sva_dfm_4_enexo_47
      | reg_act_regs_data_1_0_3_enexo_1 | reg_act_regs_data_1_0_sva_dfm_2_1_enexo);
  assign act_regs_data_and_907_enex5 = act_regs_data_and_cse & (reg_is_start_enexo_48
      | reg_w_load_lpi_1_dfm_1_enexo_48 | reg_ActUnit_PushOutput_if_output_port_reg_data_data_2_1_enexo
      | reg_act_regs_data_0_15_sva_dfm_2_1_enexo | reg_act_config_is_zero_first_sva_dfm_4_enexo_48
      | reg_act_regs_data_0_15_3_enexo_1);
  assign act_regs_data_and_908_enex5 = act_regs_data_and_cse & (reg_is_start_enexo_49
      | reg_act_regs_data_0_14_sva_dfm_2_1_enexo | reg_act_config_is_zero_first_sva_dfm_4_enexo_49
      | reg_act_regs_data_0_14_3_enexo_1 | reg_w_load_lpi_1_dfm_1_enexo_49 | reg_ActUnit_PushOutput_if_output_port_reg_data_data_14_1_enexo);
  assign act_regs_data_and_909_enex5 = act_regs_data_and_cse & (reg_act_regs_data_0_13_sva_dfm_2_1_enexo
      | reg_w_load_lpi_1_dfm_1_enexo_50 | reg_is_start_enexo_50 | reg_ActUnit_PushOutput_if_output_port_reg_data_data_13_1_enexo
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_50 | reg_act_regs_data_0_13_3_enexo_1);
  assign act_regs_data_and_910_enex5 = act_regs_data_and_cse & (reg_is_start_enexo_51
      | reg_ActUnit_PushOutput_if_output_port_reg_data_data_12_1_enexo | reg_act_config_is_zero_first_sva_dfm_4_enexo_51
      | reg_act_regs_data_0_12_3_enexo_1 | reg_act_regs_data_0_12_sva_dfm_2_1_enexo
      | reg_w_load_lpi_1_dfm_1_enexo_51);
  assign act_regs_data_and_911_enex5 = act_regs_data_and_cse & (reg_act_config_is_zero_first_sva_dfm_4_enexo_52
      | reg_act_regs_data_0_11_sva_dfm_2_1_enexo | reg_is_start_enexo_52 | reg_ActUnit_PushOutput_if_output_port_reg_data_data_11_1_enexo
      | reg_w_load_lpi_1_dfm_1_enexo_52 | reg_act_regs_data_0_11_3_enexo_1);
  assign act_regs_data_and_912_enex5 = act_regs_data_and_cse & (reg_is_start_enexo_53
      | reg_w_load_lpi_1_dfm_1_enexo_53 | reg_act_regs_data_0_10_sva_dfm_2_1_enexo
      | reg_act_regs_data_0_10_3_enexo_1 | reg_ActUnit_PushOutput_if_output_port_reg_data_data_10_1_enexo
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_53);
  assign act_regs_data_and_913_enex5 = act_regs_data_and_cse & (reg_act_regs_data_0_9_sva_dfm_2_1_enexo
      | reg_is_start_enexo_54 | reg_w_load_lpi_1_dfm_1_enexo_54 | reg_act_config_is_zero_first_sva_dfm_4_enexo_54
      | reg_act_regs_data_0_9_3_enexo_1 | reg_act_regs_data_0_0_3_enexo);
  assign act_regs_data_and_914_enex5 = act_regs_data_and_cse & (reg_w_load_lpi_1_dfm_1_enexo_55
      | reg_is_start_enexo_55 | reg_ActUnit_PushOutput_if_output_port_reg_data_data_9_1_enexo
      | reg_act_regs_data_0_8_3_enexo_1 | reg_act_config_is_zero_first_sva_dfm_4_enexo_55
      | reg_act_regs_data_0_8_sva_dfm_2_1_enexo);
  assign act_regs_data_and_915_enex5 = act_regs_data_and_cse & (reg_is_start_enexo_56
      | reg_act_regs_data_0_7_sva_dfm_2_1_enexo | reg_w_load_lpi_1_dfm_1_enexo_56
      | reg_ActUnit_PushOutput_if_output_port_reg_data_data_8_1_enexo | reg_act_config_is_zero_first_sva_dfm_4_enexo_56
      | reg_act_regs_data_0_7_3_enexo_1);
  assign act_regs_data_and_916_enex5 = act_regs_data_and_cse & (reg_is_start_enexo_57
      | reg_ActUnit_PushOutput_if_output_port_reg_data_data_7_1_enexo | reg_w_load_lpi_1_dfm_1_enexo_57
      | reg_act_regs_data_0_6_3_enexo_1 | reg_act_regs_data_0_6_sva_dfm_2_1_enexo
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_57);
  assign act_regs_data_and_917_enex5 = act_regs_data_and_cse & (reg_is_start_enexo_58
      | reg_act_regs_data_0_5_sva_dfm_2_1_enexo | reg_act_regs_data_0_5_3_enexo_1
      | reg_ActUnit_PushOutput_if_output_port_reg_data_data_6_1_enexo | reg_w_load_lpi_1_dfm_1_enexo_58
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_58);
  assign act_regs_data_and_918_enex5 = act_regs_data_and_cse & (reg_act_config_is_zero_first_sva_dfm_4_enexo_59
      | reg_w_load_lpi_1_dfm_1_enexo_59 | reg_ActUnit_PushOutput_if_output_port_reg_data_data_5_1_enexo
      | reg_act_regs_data_0_4_3_enexo_1 | reg_is_start_enexo_59 | reg_act_regs_data_0_4_sva_dfm_2_1_enexo);
  assign act_regs_data_and_919_enex5 = act_regs_data_and_cse & (reg_ActUnit_PushOutput_if_output_port_reg_data_data_4_1_enexo
      | reg_act_regs_data_0_3_3_enexo_1 | reg_is_start_enexo_60 | reg_act_config_is_zero_first_sva_dfm_4_enexo_60
      | reg_act_regs_data_0_3_sva_dfm_2_1_enexo | reg_w_load_lpi_1_dfm_1_enexo_60);
  assign act_regs_data_and_920_enex5 = act_regs_data_and_cse & (reg_act_regs_data_0_2_3_enexo_1
      | reg_w_load_lpi_1_dfm_1_enexo_61 | reg_act_regs_data_0_2_sva_dfm_2_1_enexo
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_61 | reg_ActUnit_PushOutput_if_output_port_reg_data_data_3_1_enexo
      | reg_is_start_enexo_61);
  assign act_regs_data_and_921_enex5 = act_regs_data_and_cse & (reg_act_config_is_zero_first_sva_dfm_4_enexo_62
      | reg_w_load_lpi_1_dfm_1_enexo_62 | reg_act_regs_data_0_1_3_enexo_1 | reg_ActUnit_PushOutput_if_output_port_reg_data_data_1_1_enexo
      | reg_is_start_enexo_62 | reg_act_regs_data_0_1_sva_dfm_2_1_enexo);
  assign act_regs_data_and_922_enex5 = act_regs_data_and_cse & (reg_is_start_enexo_63
      | reg_w_load_lpi_1_dfm_1_enexo_63 | reg_ActUnit_PushOutput_if_output_port_reg_data_data_0_1_enexo
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_63 | reg_act_regs_data_0_0_sva_dfm_2_1_enexo
      | reg_act_regs_data_0_0_3_enexo_1);
  assign act_mem_banks_read_read_data_and_cse = ActUnitRun_wen & and_dcpl_590 & and_dcpl_563
      & (~ (fsm_output[4])) & act_read_req_valid_lpi_1_dfm_6 & (~ ActUnit_CheckStart_start_reg_sva);
  assign act_mem_banks_read_read_data_and_16_enex5 = act_mem_banks_read_read_data_and_cse
      & reg_act_mem_banks_read_for_mux_15_enexo;
  assign act_mem_banks_read_read_data_and_17_enex5 = act_mem_banks_read_read_data_and_cse
      & reg_act_mem_banks_read_for_mux_14_enexo;
  assign act_mem_banks_read_read_data_and_18_enex5 = act_mem_banks_read_read_data_and_cse
      & reg_act_mem_banks_read_for_mux_13_enexo;
  assign act_mem_banks_read_read_data_and_19_enex5 = act_mem_banks_read_read_data_and_cse
      & reg_act_mem_banks_read_for_mux_12_enexo;
  assign act_mem_banks_read_read_data_and_20_enex5 = act_mem_banks_read_read_data_and_cse
      & reg_act_mem_banks_read_for_mux_11_enexo;
  assign act_mem_banks_read_read_data_and_21_enex5 = act_mem_banks_read_read_data_and_cse
      & reg_act_mem_banks_read_for_mux_10_enexo;
  assign act_mem_banks_read_read_data_and_22_enex5 = act_mem_banks_read_read_data_and_cse
      & reg_act_mem_banks_read_for_mux_9_enexo;
  assign act_mem_banks_read_read_data_and_23_enex5 = act_mem_banks_read_read_data_and_cse
      & reg_act_mem_banks_read_for_mux_8_enexo;
  assign act_mem_banks_read_read_data_and_24_enex5 = act_mem_banks_read_read_data_and_cse
      & reg_act_mem_banks_read_for_mux_7_enexo;
  assign act_mem_banks_read_read_data_and_25_enex5 = act_mem_banks_read_read_data_and_cse
      & reg_act_mem_banks_read_for_mux_6_enexo;
  assign act_mem_banks_read_read_data_and_26_enex5 = act_mem_banks_read_read_data_and_cse
      & reg_act_mem_banks_read_for_mux_5_enexo;
  assign act_mem_banks_read_read_data_and_27_enex5 = act_mem_banks_read_read_data_and_cse
      & reg_act_mem_banks_read_for_mux_4_enexo;
  assign act_mem_banks_read_read_data_and_28_enex5 = act_mem_banks_read_read_data_and_cse
      & reg_act_mem_banks_read_for_mux_3_enexo;
  assign act_mem_banks_read_read_data_and_29_enex5 = act_mem_banks_read_read_data_and_cse
      & reg_act_mem_banks_read_for_mux_2_enexo;
  assign act_mem_banks_read_read_data_and_30_enex5 = act_mem_banks_read_read_data_and_cse
      & reg_act_mem_banks_read_for_mux_1_enexo;
  assign act_mem_banks_read_read_data_and_31_enex5 = act_mem_banks_read_read_data_and_cse
      & reg_act_mem_banks_read_for_mux_enexo;
  assign act_port_read_out_data_and_cse = ActUnitRun_wen & and_dcpl_591 & nor_57_cse
      & act_read_req_valid_lpi_1_dfm_6;
  assign act_port_read_out_data_and_16_enex5 = act_port_read_out_data_and_cse & (reg_act_mem_banks_read_for_mux_15_enexo_1
      | reg_act_mem_banks_read_read_data_lpi_1_dfm_1_31_0_enexo | reg_ActUnit_CheckStart_start_reg_enexo);
  assign act_port_read_out_data_and_17_enex5 = act_port_read_out_data_and_cse & (reg_ActUnit_CheckStart_start_reg_enexo_1
      | reg_act_mem_banks_read_for_mux_14_enexo_1 | reg_act_mem_banks_read_read_data_lpi_1_dfm_1_63_32_enexo);
  assign act_port_read_out_data_and_18_enex5 = act_port_read_out_data_and_cse & (reg_ActUnit_CheckStart_start_reg_enexo_2
      | reg_act_mem_banks_read_read_data_lpi_1_dfm_1_95_64_enexo | reg_act_mem_banks_read_for_mux_13_enexo_1);
  assign act_port_read_out_data_and_19_enex5 = act_port_read_out_data_and_cse & (reg_ActUnit_CheckStart_start_reg_enexo_3
      | reg_act_mem_banks_read_read_data_lpi_1_dfm_1_127_96_enexo | reg_act_mem_banks_read_for_mux_12_enexo_1);
  assign act_port_read_out_data_and_20_enex5 = act_port_read_out_data_and_cse & (reg_act_mem_banks_read_for_mux_11_enexo_1
      | reg_ActUnit_CheckStart_start_reg_enexo_4 | reg_act_mem_banks_read_read_data_lpi_1_dfm_1_159_128_enexo);
  assign act_port_read_out_data_and_21_enex5 = act_port_read_out_data_and_cse & (reg_ActUnit_CheckStart_start_reg_enexo_5
      | reg_act_mem_banks_read_read_data_lpi_1_dfm_1_191_160_enexo | reg_act_mem_banks_read_for_mux_10_enexo_1);
  assign act_port_read_out_data_and_22_enex5 = act_port_read_out_data_and_cse & (reg_act_mem_banks_read_for_mux_9_enexo_1
      | reg_ActUnit_CheckStart_start_reg_enexo_6 | reg_act_mem_banks_read_read_data_lpi_1_dfm_1_223_192_enexo);
  assign act_port_read_out_data_and_23_enex5 = act_port_read_out_data_and_cse & (reg_act_mem_banks_read_for_mux_8_enexo_1
      | reg_ActUnit_CheckStart_start_reg_enexo_7 | reg_act_mem_banks_read_read_data_lpi_1_dfm_1_255_224_enexo);
  assign act_port_read_out_data_and_24_enex5 = act_port_read_out_data_and_cse & (reg_act_mem_banks_read_for_mux_7_enexo_1
      | reg_ActUnit_CheckStart_start_reg_enexo_8 | reg_act_mem_banks_read_read_data_lpi_1_dfm_1_287_256_enexo);
  assign act_port_read_out_data_and_25_enex5 = act_port_read_out_data_and_cse & (reg_ActUnit_CheckStart_start_reg_enexo_9
      | reg_act_mem_banks_read_read_data_lpi_1_dfm_1_319_288_enexo | reg_act_mem_banks_read_for_mux_6_enexo_1);
  assign act_port_read_out_data_and_26_enex5 = act_port_read_out_data_and_cse & (reg_act_mem_banks_read_for_mux_5_enexo_1
      | reg_ActUnit_CheckStart_start_reg_enexo_10 | reg_act_mem_banks_read_read_data_lpi_1_dfm_1_351_320_enexo);
  assign act_port_read_out_data_and_27_enex5 = act_port_read_out_data_and_cse & (reg_ActUnit_CheckStart_start_reg_enexo_11
      | reg_act_mem_banks_read_read_data_lpi_1_dfm_1_383_352_enexo | reg_act_mem_banks_read_for_mux_4_enexo_1);
  assign act_port_read_out_data_and_28_enex5 = act_port_read_out_data_and_cse & (reg_act_mem_banks_read_read_data_lpi_1_dfm_1_415_384_enexo
      | reg_ActUnit_CheckStart_start_reg_enexo_12 | reg_act_mem_banks_read_for_mux_3_enexo_1);
  assign act_port_read_out_data_and_29_enex5 = act_port_read_out_data_and_cse & (reg_act_mem_banks_read_read_data_lpi_1_dfm_1_447_416_enexo
      | reg_act_mem_banks_read_for_mux_2_enexo_1 | reg_ActUnit_CheckStart_start_reg_enexo_13);
  assign act_port_read_out_data_and_30_enex5 = act_port_read_out_data_and_cse & (reg_act_mem_banks_read_for_mux_1_enexo_1
      | reg_ActUnit_CheckStart_start_reg_enexo_14 | reg_act_mem_banks_read_read_data_lpi_1_dfm_1_479_448_enexo);
  assign act_port_read_out_data_and_31_enex5 = act_port_read_out_data_and_cse & (reg_ActUnit_CheckStart_start_reg_enexo_15
      | reg_act_mem_banks_read_read_data_lpi_1_dfm_1_511_480_enexo | reg_act_mem_banks_read_for_mux_enexo_1);
  assign Tanh_for_and_85_m1c = w_axi_rsp_lpi_1_dfm_1 & and_dcpl_794;
  assign Tanh_for_or_cse = and_dcpl_768 | ((~ w_axi_rsp_lpi_1_dfm_1) & and_dcpl_794)
      | ((~ act_read_req_valid_lpi_1_dfm_6) & Tanh_for_and_85_m1c);
  assign Tanh_for_and_87_cse = act_read_req_valid_lpi_1_dfm_6 & Tanh_for_and_85_m1c;
  assign mux_198_nl = MUX_s_1_2_2(nor_tmp_46, mux_tmp_197, fsm_output[1]);
  assign mux_199_nl = MUX_s_1_2_2(mux_198_nl, or_tmp_315, fsm_output[4]);
  assign ActUnit_PushOutput_if_for_and_28_cse = ActUnitRun_wen & mux_199_nl;
  assign or_1033_cse = (fsm_output[3:2]!=2'b00);
  assign and_nl = act_read_req_valid_lpi_1_dfm_6 & w_axi_rsp_lpi_1_dfm_1 & (fsm_output[1])
      & (fsm_output[4]);
  assign nor_710_nl = ~((~ (fsm_output[1])) | (fsm_output[4]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | rva_in_PopNB_mioi_data_rw_rsc_z_mxwt | is_start_sva | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11:8]!=4'b1000));
  assign mux_297_nl = MUX_s_1_2_2(and_nl, nor_710_nl, fsm_output[0]);
  assign nor_711_nl = ~((~ (fsm_output[4])) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | rva_in_PopNB_mioi_data_rw_rsc_z_mxwt | is_start_sva | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11:8]!=4'b1000));
  assign mux_298_nl = MUX_s_1_2_2(mux_297_nl, nor_711_nl, or_1033_cse);
  assign and_1211_cse = mux_298_nl & ActUnitRun_wen;
  assign mux_201_nl = MUX_s_1_2_2((~ or_tmp_315), or_1033_cse, fsm_output[4]);
  assign mux_200_nl = MUX_s_1_2_2((~ or_tmp_315), or_tmp_317, fsm_output[4]);
  assign and_1094_nl = act_read_req_valid_lpi_1_dfm_6 & w_axi_rsp_lpi_1_dfm_1;
  assign mux_202_nl = MUX_s_1_2_2(mux_201_nl, mux_200_nl, and_1094_nl);
  assign rva_out_reg_data_and_16_cse = ActUnitRun_wen & ((~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11:9]!=3'b100)
      | or_dcpl_300 | is_start_sva | (~ mux_202_nl))) | and_dcpl_803);
  assign mux_204_nl = MUX_s_1_2_2(mux_tmp_203, and_dcpl_770, fsm_output[1]);
  assign ActUnit_RunInst_switch_lp_and_802_cse = ActUnitRun_wen & (mux_204_nl | (fsm_output[4]));
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc = ActUnit_RunInst_switch_lp_and_802_cse
      & and_dcpl_9 & (~ (act_config_in_InstFetch_mux_tmp[7])) & (act_config_in_InstFetch_mux_tmp[6])
      & (act_config_in_InstFetch_mux_tmp[4]);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_37_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_17_sva_dfm_6_enexo | reg_act_config_inst_regs_1_sva_dfm_5_enexo
      | reg_act_regs_data_0_15_2_enexo | reg_act_config_inst_counter_enexo | reg_act_regs_data_2_15_2_enexo
      | reg_act_regs_data_3_15_2_enexo | reg_act_regs_data_1_15_2_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_38_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_1_sva_dfm_5_enexo_1 | reg_act_config_inst_regs_17_sva_dfm_6_enexo_1
      | reg_act_config_inst_counter_enexo_1 | reg_act_regs_data_2_14_2_enexo | reg_act_regs_data_0_14_2_enexo
      | reg_act_regs_data_3_14_2_enexo | reg_act_regs_data_1_14_2_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_39_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_1_sva_dfm_5_enexo_2 | reg_act_config_inst_regs_17_sva_dfm_6_enexo_2
      | reg_act_config_inst_counter_enexo_2 | reg_act_regs_data_3_13_2_enexo | reg_act_regs_data_1_13_2_enexo
      | reg_act_regs_data_0_13_2_enexo | reg_act_regs_data_2_13_2_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_40_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_17_sva_dfm_6_enexo_3 | reg_act_config_inst_regs_1_sva_dfm_5_enexo_3
      | reg_act_regs_data_0_12_2_enexo | reg_act_regs_data_1_12_2_enexo | reg_act_regs_data_2_12_2_enexo
      | reg_act_regs_data_3_12_2_enexo | reg_act_config_inst_counter_enexo_3);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_41_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_1_sva_dfm_5_enexo_4 | reg_act_config_inst_regs_17_sva_dfm_6_enexo_4
      | reg_act_regs_data_0_11_2_enexo | reg_act_regs_data_3_11_2_enexo | reg_act_regs_data_2_11_2_enexo
      | reg_act_regs_data_1_11_2_enexo | reg_act_config_inst_counter_enexo_4);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_42_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_1_sva_dfm_5_enexo_5 | reg_act_config_inst_regs_17_sva_dfm_6_enexo_5
      | reg_act_regs_data_3_10_2_enexo | reg_act_regs_data_0_10_2_enexo | reg_act_regs_data_2_10_2_enexo
      | reg_act_config_inst_counter_enexo_5 | reg_act_regs_data_1_10_2_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_43_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_1_sva_dfm_5_enexo_6 | reg_act_regs_data_1_9_2_enexo
      | reg_act_config_inst_regs_17_sva_dfm_6_enexo_6 | reg_act_config_inst_counter_enexo_6
      | reg_act_regs_data_2_9_2_enexo | reg_act_regs_data_0_9_2_enexo | reg_act_regs_data_3_9_2_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_44_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_regs_data_3_8_2_enexo | reg_act_config_inst_regs_17_sva_dfm_6_enexo_7
      | reg_act_config_inst_regs_1_sva_dfm_5_enexo_7 | reg_act_regs_data_1_8_2_enexo
      | reg_act_regs_data_0_8_2_enexo | reg_act_regs_data_2_8_2_enexo | reg_act_config_inst_counter_enexo_7);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_45_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_regs_data_1_7_2_enexo | reg_act_config_inst_regs_17_sva_dfm_6_enexo_8
      | reg_act_config_inst_regs_1_sva_dfm_5_enexo_8 | reg_act_regs_data_2_7_2_enexo
      | reg_act_regs_data_3_7_2_enexo | reg_act_regs_data_0_7_2_enexo | reg_act_config_inst_counter_enexo_8);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_46_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_17_sva_dfm_6_enexo_9 | reg_act_config_inst_counter_enexo_9
      | reg_act_config_inst_regs_1_sva_dfm_5_enexo_9 | reg_act_regs_data_2_6_2_enexo
      | reg_act_regs_data_0_6_2_enexo | reg_act_regs_data_3_6_2_enexo | reg_act_regs_data_1_6_2_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_47_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_regs_data_3_5_2_enexo | reg_act_config_inst_regs_1_sva_dfm_5_enexo_10
      | reg_act_regs_data_1_5_2_enexo | reg_act_config_inst_regs_17_sva_dfm_6_enexo_10
      | reg_act_regs_data_2_5_2_enexo | reg_act_regs_data_0_5_2_enexo | reg_act_config_inst_counter_enexo_10);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_48_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_17_sva_dfm_6_enexo_11 | reg_act_config_inst_regs_1_sva_dfm_5_enexo_11
      | reg_act_config_inst_counter_enexo_11 | reg_act_regs_data_0_4_2_enexo | reg_act_regs_data_3_4_2_enexo
      | reg_act_regs_data_2_4_2_enexo | reg_act_regs_data_1_4_2_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_49_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_17_sva_dfm_6_enexo_12 | reg_act_regs_data_3_3_2_enexo
      | reg_act_config_inst_regs_1_sva_dfm_5_enexo_12 | reg_act_config_inst_counter_enexo_12
      | reg_act_regs_data_1_3_2_enexo | reg_act_regs_data_0_3_2_enexo | reg_act_regs_data_2_3_2_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_50_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_1_sva_dfm_5_enexo_13 | reg_act_config_inst_regs_17_sva_dfm_6_enexo_13
      | reg_act_regs_data_2_2_2_enexo | reg_act_regs_data_0_2_2_enexo | reg_act_regs_data_3_2_2_enexo
      | reg_act_config_inst_counter_enexo_13 | reg_act_regs_data_1_2_2_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_51_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_1_sva_dfm_5_enexo_14 | reg_act_config_inst_regs_17_sva_dfm_6_enexo_14
      | reg_act_regs_data_0_1_2_enexo | reg_act_config_inst_counter_enexo_14 | reg_act_regs_data_3_1_2_enexo
      | reg_act_regs_data_2_1_2_enexo | reg_act_regs_data_1_1_2_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_52_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_1_sva_dfm_5_enexo_15 | reg_act_regs_data_2_0_2_enexo
      | reg_act_regs_data_3_0_2_enexo | reg_act_regs_data_0_0_2_enexo | reg_act_config_inst_regs_17_sva_dfm_6_enexo_15
      | reg_act_regs_data_1_0_2_enexo | reg_act_config_inst_counter_enexo_15);
  assign Relu_for_y_qelse_and_cse = ActUnit_RunInst_switch_lp_and_802_cse & is_start_sva
      & (~ (act_config_in_InstFetch_mux_tmp[5])) & (act_config_in_InstFetch_mux_tmp[7])
      & and_dcpl_47;
  assign Relu_for_y_qelse_and_31_enex5 = Relu_for_y_qelse_and_cse & (reg_act_config_inst_regs_1_sva_dfm_5_enexo_16
      | reg_act_regs_data_0_15_2_enexo_1 | reg_act_config_inst_regs_17_sva_dfm_6_enexo_16
      | reg_act_regs_data_3_15_enexo | reg_act_regs_data_2_15_2_enexo_1 | reg_act_regs_data_3_15_2_enexo_1
      | reg_act_regs_data_1_15_2_enexo_1 | reg_act_config_inst_counter_enexo_16);
  assign Relu_for_y_qelse_and_32_enex5 = Relu_for_y_qelse_and_cse & (reg_act_regs_data_0_14_2_enexo_1
      | reg_act_config_inst_regs_1_sva_dfm_5_enexo_17 | reg_act_config_inst_regs_17_sva_dfm_6_enexo_17
      | reg_act_regs_data_1_14_enexo | reg_act_regs_data_1_14_2_enexo_1 | reg_act_config_inst_counter_enexo_17
      | reg_act_regs_data_3_14_2_enexo_1 | reg_act_regs_data_2_14_2_enexo_1);
  assign Relu_for_y_qelse_and_33_enex5 = Relu_for_y_qelse_and_cse & (reg_act_config_inst_regs_1_sva_dfm_5_enexo_18
      | reg_act_config_inst_regs_17_sva_dfm_6_enexo_18 | reg_act_regs_data_1_13_enexo
      | reg_act_config_inst_counter_enexo_18 | reg_act_regs_data_3_13_2_enexo_1 |
      reg_act_regs_data_2_13_2_enexo_1 | reg_act_regs_data_0_13_2_enexo_1 | reg_act_regs_data_1_13_2_enexo_1);
  assign Relu_for_y_qelse_and_34_enex5 = Relu_for_y_qelse_and_cse & (reg_act_config_inst_regs_1_sva_dfm_5_enexo_19
      | reg_act_regs_data_0_12_2_enexo_1 | reg_act_config_inst_regs_17_sva_dfm_6_enexo_19
      | reg_act_regs_data_1_12_enexo | reg_act_regs_data_3_12_2_enexo_1 | reg_act_config_inst_counter_enexo_19
      | reg_act_regs_data_1_12_2_enexo_1 | reg_act_regs_data_2_12_2_enexo_1);
  assign Relu_for_y_qelse_and_35_enex5 = Relu_for_y_qelse_and_cse & (reg_act_config_inst_regs_17_sva_dfm_6_enexo_20
      | reg_act_config_inst_regs_1_sva_dfm_5_enexo_20 | reg_act_regs_data_0_11_2_enexo_1
      | reg_act_config_inst_counter_enexo_20 | reg_act_regs_data_3_11_2_enexo_1 |
      reg_act_regs_data_1_11_enexo | reg_act_regs_data_1_11_2_enexo_1 | reg_act_regs_data_2_11_2_enexo_1);
  assign Relu_for_y_qelse_and_36_enex5 = Relu_for_y_qelse_and_cse & (reg_act_config_inst_regs_17_sva_dfm_6_enexo_21
      | reg_act_regs_data_2_10_enexo | reg_act_regs_data_3_10_2_enexo_1 | reg_act_config_inst_regs_1_sva_dfm_5_enexo_21
      | reg_act_regs_data_0_10_2_enexo_1 | reg_act_config_inst_counter_enexo_21 |
      reg_act_regs_data_1_10_2_enexo_1 | reg_act_regs_data_2_10_2_enexo_1);
  assign Relu_for_y_qelse_and_37_enex5 = Relu_for_y_qelse_and_cse & (reg_act_regs_data_0_9_enexo
      | reg_act_regs_data_0_9_2_enexo_1 | reg_act_config_inst_regs_17_sva_dfm_6_enexo_22
      | reg_act_config_inst_regs_1_sva_dfm_5_enexo_22 | reg_act_config_inst_counter_enexo_22
      | reg_act_regs_data_3_9_2_enexo_1 | reg_act_regs_data_1_9_2_enexo_1 | reg_act_regs_data_2_9_2_enexo_1);
  assign Relu_for_y_qelse_and_38_enex5 = Relu_for_y_qelse_and_cse & (reg_act_config_inst_regs_1_sva_dfm_5_enexo_23
      | reg_act_config_inst_regs_17_sva_dfm_6_enexo_23 | reg_act_regs_data_2_8_2_enexo_1
      | reg_act_regs_data_3_8_2_enexo_1 | reg_act_regs_data_0_8_enexo | reg_act_regs_data_0_8_2_enexo_1
      | reg_act_regs_data_1_8_2_enexo_1 | reg_act_config_inst_counter_enexo_23);
  assign Relu_for_y_qelse_and_39_enex5 = Relu_for_y_qelse_and_cse & (reg_act_config_inst_regs_17_sva_dfm_6_enexo_24
      | reg_act_regs_data_1_7_enexo | reg_act_regs_data_1_7_2_enexo_1 | reg_act_config_inst_regs_1_sva_dfm_5_enexo_24
      | reg_act_regs_data_0_7_2_enexo_1 | reg_act_regs_data_3_7_2_enexo_1 | reg_act_regs_data_2_7_2_enexo_1
      | reg_act_config_inst_counter_enexo_24);
  assign Relu_for_y_qelse_and_40_enex5 = Relu_for_y_qelse_and_cse & (reg_act_config_inst_regs_17_sva_dfm_6_enexo_25
      | reg_act_config_inst_regs_1_sva_dfm_5_enexo_25 | reg_act_regs_data_2_6_2_enexo_1
      | reg_act_regs_data_2_6_enexo | reg_act_regs_data_0_6_2_enexo_1 | reg_act_config_inst_counter_enexo_25
      | reg_act_regs_data_3_6_2_enexo_1 | reg_act_regs_data_1_6_2_enexo_1);
  assign Relu_for_y_qelse_and_41_enex5 = Relu_for_y_qelse_and_cse & (reg_act_config_inst_regs_17_sva_dfm_6_enexo_26
      | reg_act_config_inst_regs_1_sva_dfm_5_enexo_26 | reg_act_regs_data_3_5_enexo
      | reg_act_regs_data_0_5_2_enexo_1 | reg_act_regs_data_1_5_2_enexo_1 | reg_act_regs_data_2_5_2_enexo_1
      | reg_act_regs_data_3_5_2_enexo_1 | reg_act_config_inst_counter_enexo_26);
  assign Relu_for_y_qelse_and_42_enex5 = Relu_for_y_qelse_and_cse & (reg_act_config_inst_regs_17_sva_dfm_6_enexo_27
      | reg_act_regs_data_1_4_2_enexo_1 | reg_act_config_inst_counter_enexo_27 |
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_27 | reg_act_regs_data_1_4_enexo
      | reg_act_regs_data_0_4_2_enexo_1 | reg_act_regs_data_3_4_2_enexo_1 | reg_act_regs_data_2_4_2_enexo_1);
  assign Relu_for_y_qelse_and_43_enex5 = Relu_for_y_qelse_and_cse & (reg_act_config_inst_regs_17_sva_dfm_6_enexo_28
      | reg_act_regs_data_0_3_enexo | reg_act_config_inst_regs_1_sva_dfm_5_enexo_28
      | reg_act_config_inst_counter_enexo_28 | reg_act_regs_data_2_3_2_enexo_1 |
      reg_act_regs_data_1_3_2_enexo_1 | reg_act_regs_data_3_3_2_enexo_1 | reg_act_regs_data_0_3_2_enexo_1);
  assign Relu_for_y_qelse_and_44_enex5 = Relu_for_y_qelse_and_cse & (reg_act_config_inst_regs_17_sva_dfm_6_enexo_29
      | reg_act_config_inst_regs_1_sva_dfm_5_enexo_29 | reg_act_regs_data_2_2_2_enexo_1
      | reg_act_regs_data_1_2_enexo | reg_act_regs_data_0_2_2_enexo_1 | reg_act_config_inst_counter_enexo_29
      | reg_act_regs_data_3_2_2_enexo_1 | reg_act_regs_data_1_2_2_enexo_1);
  assign Relu_for_y_qelse_and_45_enex5 = Relu_for_y_qelse_and_cse & (reg_act_config_inst_regs_17_sva_dfm_6_enexo_30
      | reg_act_config_inst_regs_1_sva_dfm_5_enexo_30 | reg_act_regs_data_0_1_enexo
      | reg_act_regs_data_0_1_2_enexo_1 | reg_act_regs_data_2_1_2_enexo_1 | reg_act_config_inst_counter_enexo_30
      | reg_act_regs_data_1_1_2_enexo_1 | reg_act_regs_data_3_1_2_enexo_1);
  assign Relu_for_y_qelse_and_46_enex5 = Relu_for_y_qelse_and_cse & (reg_act_config_inst_regs_1_sva_dfm_5_enexo_31
      | reg_act_config_inst_regs_17_sva_dfm_6_enexo_31 | reg_act_regs_data_1_0_2_enexo_1
      | reg_act_regs_data_2_0_enexo | reg_act_config_inst_counter_enexo_31 | reg_act_regs_data_0_0_2_enexo_1
      | reg_act_regs_data_3_0_2_enexo_1 | reg_act_regs_data_2_0_2_enexo_1);
  assign nv_scvector_cctor_nv_scvector_5_for_and_cse = ActUnitRun_wen & (~((~ mux_205_itm)
      & and_dcpl_834));
  assign nv_scvector_cctor_nv_scvector_5_for_and_15_enex5 = nv_scvector_cctor_nv_scvector_5_for_and_cse
      & (reg_act_config_inst_regs_17_sva_dfm_6_enexo_32 | reg_act_config_inst_regs_1_sva_dfm_5_enexo_32
      | reg_act_regs_data_1_2_2_enexo_2 | reg_act_regs_data_3_2_2_enexo_2 | reg_act_regs_data_0_2_2_enexo_2
      | reg_act_config_inst_counter_enexo_32 | reg_act_regs_data_2_2_2_enexo_2);
  assign nv_scvector_cctor_nv_scvector_5_for_and_16_enex5 = nv_scvector_cctor_nv_scvector_5_for_and_cse
      & (reg_act_regs_data_0_3_2_enexo_2 | reg_act_config_inst_regs_17_sva_dfm_6_enexo_33
      | reg_act_config_inst_regs_1_sva_dfm_5_enexo_33 | reg_act_config_inst_counter_enexo_33
      | reg_act_regs_data_3_3_2_enexo_2 | reg_act_regs_data_2_3_2_enexo_2 | reg_act_regs_data_1_3_2_enexo_2);
  assign ActUnit_RunInst_switch_lp_and_812_cse = ActUnitRun_wen & (~(nor_734_cse
      & and_dcpl_366));
  assign ActUnit_RunInst_switch_lp_and_815_enex5 = ActUnit_RunInst_switch_lp_and_812_cse
      & (reg_act_config_inst_regs_1_sva_dfm_5_enexo_34 | reg_act_config_inst_regs_17_sva_dfm_6_enexo_34
      | reg_act_config_inst_counter_enexo_34 | reg_act_regs_data_0_0_2_enexo_2 |
      reg_act_regs_data_3_0_2_enexo_2 | reg_act_regs_data_1_0_2_enexo_2 | reg_act_regs_data_2_0_2_enexo_2);
  assign nv_scvector_cctor_nv_scvector_5_for_and_17_enex5 = ActUnit_RunInst_switch_lp_and_812_cse
      & (reg_act_config_inst_regs_1_sva_dfm_5_enexo_35 | reg_act_config_inst_regs_17_sva_dfm_6_enexo_35
      | reg_act_regs_data_1_1_2_enexo_2 | reg_act_config_inst_counter_enexo_35 |
      reg_act_regs_data_2_1_2_enexo_2 | reg_act_regs_data_3_1_2_enexo_2 | reg_act_regs_data_0_1_2_enexo_2);
  assign nv_scvector_cctor_nv_scvector_5_for_and_3_cse = ActUnitRun_wen & (~(((fsm_output[2])
      ^ (fsm_output[1])) & and_dcpl_834));
  assign nv_scvector_cctor_nv_scvector_5_for_and_18_enex5 = nv_scvector_cctor_nv_scvector_5_for_and_3_cse
      & (reg_act_config_inst_regs_17_sva_dfm_6_enexo_36 | reg_act_config_inst_regs_1_sva_dfm_5_enexo_36
      | reg_act_regs_data_2_4_2_enexo_2 | reg_act_regs_data_0_4_2_enexo_2 | reg_act_regs_data_1_4_2_enexo_2
      | reg_act_config_inst_counter_enexo_36 | reg_act_regs_data_3_4_2_enexo_2);
  assign nv_scvector_cctor_nv_scvector_5_for_and_19_enex5 = nv_scvector_cctor_nv_scvector_5_for_and_3_cse
      & (reg_act_regs_data_1_5_2_enexo_2 | reg_act_config_inst_counter_enexo_37 |
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_37 | reg_act_config_inst_regs_1_sva_dfm_5_enexo_37
      | reg_act_regs_data_2_5_2_enexo_2 | reg_act_regs_data_0_5_2_enexo_2 | reg_act_regs_data_3_5_2_enexo_2);
  assign mux_206_nl = MUX_s_1_2_2((fsm_output[2]), nand_195_cse, fsm_output[1]);
  assign nv_scvector_cctor_nv_scvector_5_for_and_5_cse = ActUnitRun_wen & (~(mux_206_nl
      & and_dcpl_834));
  assign nv_scvector_cctor_nv_scvector_5_for_and_20_enex5 = nv_scvector_cctor_nv_scvector_5_for_and_5_cse
      & (reg_act_config_inst_regs_1_sva_dfm_5_enexo_38 | reg_act_config_inst_counter_enexo_38
      | reg_act_config_inst_regs_17_sva_dfm_6_enexo_38 | reg_act_regs_data_3_6_2_enexo_2
      | reg_act_regs_data_0_6_2_enexo_2 | reg_act_regs_data_2_6_2_enexo_2 | reg_act_regs_data_1_6_2_enexo_2);
  assign nv_scvector_cctor_nv_scvector_5_for_and_21_enex5 = nv_scvector_cctor_nv_scvector_5_for_and_5_cse
      & (reg_act_config_inst_regs_1_sva_dfm_5_enexo_39 | reg_act_config_inst_regs_17_sva_dfm_6_enexo_39
      | reg_act_regs_data_2_7_2_enexo_2 | reg_act_config_inst_counter_enexo_39 |
      reg_act_regs_data_0_7_2_enexo_2 | reg_act_regs_data_3_7_2_enexo_2 | reg_act_regs_data_1_7_2_enexo_2);
  assign nv_scvector_cctor_nv_scvector_5_for_and_7_cse = ActUnitRun_wen & (~(or_dcpl_443
      & and_dcpl_834));
  assign nv_scvector_cctor_nv_scvector_5_for_and_22_enex5 = nv_scvector_cctor_nv_scvector_5_for_and_7_cse
      & (reg_act_config_inst_regs_17_sva_dfm_6_enexo_40 | reg_act_config_inst_regs_1_sva_dfm_5_enexo_40
      | reg_act_regs_data_0_8_2_enexo_2 | reg_act_regs_data_3_8_2_enexo_2 | reg_act_regs_data_2_8_2_enexo_2
      | reg_act_config_inst_counter_enexo_40 | reg_act_regs_data_1_8_2_enexo_2);
  assign nv_scvector_cctor_nv_scvector_5_for_and_23_enex5 = nv_scvector_cctor_nv_scvector_5_for_and_7_cse
      & (reg_act_config_inst_regs_1_sva_dfm_5_enexo_41 | reg_act_config_inst_regs_17_sva_dfm_6_enexo_41
      | reg_act_config_inst_counter_enexo_41 | reg_act_regs_data_2_9_2_enexo_2 |
      reg_act_regs_data_1_9_2_enexo_2 | reg_act_regs_data_3_9_2_enexo_2 | reg_act_regs_data_0_9_2_enexo_2);
  assign mux_207_nl = MUX_s_1_2_2(mux_tmp_196, or_tmp_211, fsm_output[0]);
  assign mux_208_nl = MUX_s_1_2_2(mux_207_nl, (fsm_output[3]), fsm_output[1]);
  assign nv_scvector_cctor_nv_scvector_5_for_and_9_cse = ActUnitRun_wen & (mux_208_nl
      | (fsm_output[4]));
  assign nv_scvector_cctor_nv_scvector_5_for_and_24_enex5 = nv_scvector_cctor_nv_scvector_5_for_and_9_cse
      & (reg_act_config_inst_regs_17_sva_dfm_6_enexo_42 | reg_act_config_inst_regs_1_sva_dfm_5_enexo_42
      | reg_act_regs_data_3_10_2_enexo_2 | reg_act_regs_data_2_10_2_enexo_2 | reg_act_regs_data_1_10_2_enexo_2
      | reg_act_regs_data_0_10_2_enexo_2 | reg_act_config_inst_counter_enexo_42);
  assign nv_scvector_cctor_nv_scvector_5_for_and_25_enex5 = nv_scvector_cctor_nv_scvector_5_for_and_9_cse
      & (reg_act_config_inst_counter_enexo_43 | reg_act_config_inst_regs_17_sva_dfm_6_enexo_43
      | reg_act_config_inst_regs_1_sva_dfm_5_enexo_43 | reg_act_regs_data_2_11_2_enexo_2
      | reg_act_regs_data_1_11_2_enexo_2 | reg_act_regs_data_3_11_2_enexo_2 | reg_act_regs_data_0_11_2_enexo_2);
  assign nv_scvector_cctor_nv_scvector_5_for_and_11_cse = ActUnitRun_wen & ((~(or_dcpl_443
      ^ (fsm_output[3]))) | (fsm_output[4]));
  assign nv_scvector_cctor_nv_scvector_5_for_and_26_enex5 = nv_scvector_cctor_nv_scvector_5_for_and_11_cse
      & (reg_act_config_inst_regs_1_sva_dfm_5_enexo_44 | reg_act_config_inst_regs_17_sva_dfm_6_enexo_44
      | reg_act_regs_data_2_12_2_enexo_2 | reg_act_regs_data_3_12_2_enexo_2 | reg_act_config_inst_counter_enexo_44
      | reg_act_regs_data_1_12_2_enexo_2 | reg_act_regs_data_0_12_2_enexo_2);
  assign nv_scvector_cctor_nv_scvector_5_for_and_27_enex5 = nv_scvector_cctor_nv_scvector_5_for_and_11_cse
      & (reg_act_config_inst_regs_17_sva_dfm_6_enexo_45 | reg_act_config_inst_regs_1_sva_dfm_5_enexo_45
      | reg_act_regs_data_0_13_2_enexo_2 | reg_act_regs_data_3_13_2_enexo_2 | reg_act_regs_data_2_13_2_enexo_2
      | reg_act_config_inst_counter_enexo_45 | reg_act_regs_data_1_13_2_enexo_2);
  assign and_1096_nl = or_1071_cse & (fsm_output[3]);
  assign mux_209_nl = MUX_s_1_2_2(mux_tmp_196, and_1096_nl, fsm_output[1]);
  assign nv_scvector_cctor_nv_scvector_5_for_and_13_cse = ActUnitRun_wen & (mux_209_nl
      | (fsm_output[4]));
  assign nv_scvector_cctor_nv_scvector_5_for_and_28_enex5 = nv_scvector_cctor_nv_scvector_5_for_and_13_cse
      & (reg_act_config_inst_regs_17_sva_dfm_6_enexo_46 | reg_act_config_inst_regs_1_sva_dfm_5_enexo_46
      | reg_act_regs_data_0_14_2_enexo_2 | reg_act_regs_data_1_14_2_enexo_2 | reg_act_regs_data_3_14_2_enexo_2
      | reg_act_regs_data_2_14_2_enexo_2 | reg_act_config_inst_counter_enexo_46);
  assign nv_scvector_cctor_nv_scvector_5_for_and_29_enex5 = nv_scvector_cctor_nv_scvector_5_for_and_13_cse
      & (reg_act_config_inst_regs_17_sva_dfm_6_enexo_47 | reg_act_config_inst_regs_1_sva_dfm_5_enexo_47
      | reg_act_regs_data_3_15_2_enexo_2 | reg_act_regs_data_2_15_2_enexo_2 | reg_act_regs_data_1_15_2_enexo_2
      | reg_act_regs_data_0_15_2_enexo_2 | reg_act_config_inst_counter_enexo_47);
  assign nv_scvector_cctor_nv_scvector_6_for_and_enex5 = nv_scvector_cctor_nv_scvector_5_for_and_9_cse
      & (reg_act_config_inst_regs_17_sva_dfm_6_enexo_48 | reg_act_config_inst_regs_1_sva_dfm_5_enexo_48
      | reg_act_regs_data_2_2_2_enexo_3 | reg_act_regs_data_1_2_2_enexo_3 | reg_act_regs_data_0_2_2_enexo_3
      | reg_act_config_inst_counter_enexo_48 | reg_act_regs_data_3_2_2_enexo_3);
  assign nv_scvector_cctor_nv_scvector_6_for_and_15_enex5 = nv_scvector_cctor_nv_scvector_5_for_and_13_cse
      & (reg_act_regs_data_0_11_2_enexo_3 | reg_act_config_inst_regs_1_sva_dfm_5_enexo_49
      | reg_act_config_inst_regs_17_sva_dfm_6_enexo_49 | reg_act_regs_data_3_11_2_enexo_3
      | reg_act_regs_data_2_11_2_enexo_3 | reg_act_regs_data_1_11_2_enexo_3 | reg_act_config_inst_counter_enexo_49);
  assign ActUnit_RunInst_switch_lp_and_816_enex5 = nv_scvector_cctor_nv_scvector_5_for_and_7_cse
      & (reg_act_config_inst_regs_17_sva_dfm_6_enexo_50 | reg_act_config_inst_regs_1_sva_dfm_5_enexo_50
      | reg_act_regs_data_2_0_2_enexo_3 | reg_act_config_inst_counter_enexo_50 |
      reg_act_regs_data_0_0_2_enexo_3 | reg_act_regs_data_1_0_2_enexo_3 | reg_act_regs_data_3_0_2_enexo_3);
  assign nv_scvector_cctor_nv_scvector_6_for_and_16_enex5 = nv_scvector_cctor_nv_scvector_5_for_and_7_cse
      & (reg_act_config_inst_regs_17_sva_dfm_6_enexo_51 | reg_act_config_inst_regs_1_sva_dfm_5_enexo_51
      | reg_act_regs_data_1_1_2_enexo_3 | reg_act_config_inst_counter_enexo_51 |
      reg_act_regs_data_0_1_2_enexo_3 | reg_act_regs_data_3_1_2_enexo_3 | reg_act_regs_data_2_1_2_enexo_3);
  assign nv_scvector_cctor_nv_scvector_6_for_and_17_enex5 = nv_scvector_cctor_nv_scvector_5_for_and_11_cse
      & (reg_act_config_inst_regs_1_sva_dfm_5_enexo_52 | reg_act_config_inst_regs_17_sva_dfm_6_enexo_52
      | reg_act_regs_data_1_3_2_enexo_3 | reg_act_config_inst_counter_enexo_52 |
      reg_act_regs_data_2_3_2_enexo_3 | reg_act_regs_data_0_3_2_enexo_3 | reg_act_regs_data_3_3_2_enexo_3);
  assign nv_scvector_cctor_nv_scvector_6_for_and_18_enex5 = nv_scvector_cctor_nv_scvector_5_for_and_11_cse
      & (reg_act_config_inst_regs_1_sva_dfm_5_enexo_53 | reg_act_config_inst_regs_17_sva_dfm_6_enexo_53
      | reg_act_regs_data_0_4_2_enexo_3 | reg_act_regs_data_3_4_2_enexo_3 | reg_act_config_inst_counter_enexo_53
      | reg_act_regs_data_2_4_2_enexo_3 | reg_act_regs_data_1_4_2_enexo_3);
  assign nv_scvector_cctor_nv_scvector_6_for_and_19_enex5 = nv_scvector_cctor_nv_scvector_5_for_and_13_cse
      & (reg_act_config_inst_regs_1_sva_dfm_5_enexo_54 | reg_act_regs_data_1_5_2_enexo_3
      | reg_act_config_inst_regs_17_sva_dfm_6_enexo_54 | reg_act_config_inst_counter_enexo_54
      | reg_act_regs_data_2_5_2_enexo_3 | reg_act_regs_data_3_5_2_enexo_3 | reg_act_regs_data_0_5_2_enexo_3);
  assign nv_scvector_cctor_nv_scvector_6_for_and_20_enex5 = nv_scvector_cctor_nv_scvector_5_for_and_13_cse
      & (reg_act_config_inst_regs_1_sva_dfm_5_enexo_55 | reg_act_regs_data_1_6_2_enexo_3
      | reg_act_config_inst_counter_enexo_55 | reg_act_config_inst_regs_17_sva_dfm_6_enexo_55
      | reg_act_regs_data_3_6_2_enexo_3 | reg_act_regs_data_0_6_2_enexo_3 | reg_act_regs_data_2_6_2_enexo_3);
  assign mux_210_nl = MUX_s_1_2_2(mux_tmp_196, and_dcpl_770, fsm_output[1]);
  assign nv_scvector_cctor_nv_scvector_6_for_and_7_cse = ActUnitRun_wen & (mux_210_nl
      | (fsm_output[4]));
  assign nv_scvector_cctor_nv_scvector_6_for_and_21_enex5 = nv_scvector_cctor_nv_scvector_6_for_and_7_cse
      & (reg_act_config_inst_regs_17_sva_dfm_6_enexo_56 | reg_act_config_inst_counter_enexo_56
      | reg_act_config_inst_regs_1_sva_dfm_5_enexo_56 | reg_act_regs_data_0_7_2_enexo_3
      | reg_act_regs_data_3_7_2_enexo_3 | reg_act_regs_data_1_7_2_enexo_3 | reg_act_regs_data_2_7_2_enexo_3);
  assign nv_scvector_cctor_nv_scvector_6_for_and_22_enex5 = nv_scvector_cctor_nv_scvector_6_for_and_7_cse
      & (reg_act_config_inst_regs_17_sva_dfm_6_enexo_57 | reg_act_config_inst_counter_enexo_57
      | reg_act_config_inst_regs_1_sva_dfm_5_enexo_57 | reg_act_regs_data_1_8_2_enexo_3
      | reg_act_regs_data_3_8_2_enexo_3 | reg_act_regs_data_2_8_2_enexo_3 | reg_act_regs_data_0_8_2_enexo_3);
  assign nv_scvector_cctor_nv_scvector_6_for_and_23_enex5 = ActUnit_RunInst_switch_lp_and_802_cse
      & (reg_act_config_inst_regs_17_sva_dfm_6_enexo_58 | reg_act_regs_data_3_9_2_enexo_3
      | reg_act_config_inst_regs_1_sva_dfm_5_enexo_58 | reg_act_config_inst_counter_enexo_58
      | reg_act_regs_data_1_9_2_enexo_3 | reg_act_regs_data_0_9_2_enexo_3 | reg_act_regs_data_2_9_2_enexo_3);
  assign nv_scvector_cctor_nv_scvector_6_for_and_24_enex5 = ActUnit_RunInst_switch_lp_and_802_cse
      & (reg_act_config_inst_regs_1_sva_dfm_5_enexo_59 | reg_act_config_inst_regs_17_sva_dfm_6_enexo_59
      | reg_act_regs_data_0_10_2_enexo_3 | reg_act_regs_data_3_10_2_enexo_3 | reg_act_config_inst_counter_enexo_59
      | reg_act_regs_data_2_10_2_enexo_3 | reg_act_regs_data_1_10_2_enexo_3);
  assign nv_scvector_cctor_nv_scvector_6_for_and_25_enex5 = nv_scvector_cctor_nv_scvector_6_for_and_7_cse
      & (reg_act_config_inst_regs_17_sva_dfm_6_enexo_60 | reg_act_config_inst_regs_1_sva_dfm_5_enexo_60
      | reg_act_regs_data_3_12_2_enexo_3 | reg_act_regs_data_0_12_2_enexo_3 | reg_act_config_inst_counter_enexo_60
      | reg_act_regs_data_2_12_2_enexo_3 | reg_act_regs_data_1_12_2_enexo_3);
  assign nv_scvector_cctor_nv_scvector_6_for_and_26_enex5 = nv_scvector_cctor_nv_scvector_6_for_and_7_cse
      & (reg_act_config_inst_regs_1_sva_dfm_5_enexo_61 | reg_act_config_inst_regs_17_sva_dfm_6_enexo_61
      | reg_act_regs_data_0_13_2_enexo_3 | reg_act_regs_data_3_13_2_enexo_3 | reg_act_regs_data_1_13_2_enexo_3
      | reg_act_regs_data_2_13_2_enexo_3 | reg_act_config_inst_counter_enexo_61);
  assign nv_scvector_cctor_nv_scvector_6_for_and_27_enex5 = nv_scvector_cctor_nv_scvector_6_for_and_7_cse
      & (reg_act_regs_data_3_14_2_enexo_3 | reg_act_config_inst_regs_1_sva_dfm_5_enexo_62
      | reg_act_config_inst_regs_17_sva_dfm_6_enexo_62 | reg_act_regs_data_2_14_2_enexo_3
      | reg_act_regs_data_0_14_2_enexo_3 | reg_act_regs_data_1_14_2_enexo_3 | reg_act_config_inst_counter_enexo_62);
  assign nv_scvector_cctor_nv_scvector_6_for_and_28_enex5 = ActUnit_RunInst_switch_lp_and_802_cse
      & (reg_act_config_inst_regs_1_sva_dfm_5_enexo_63 | reg_act_config_inst_regs_17_sva_dfm_6_enexo_63
      | reg_act_regs_data_3_15_2_enexo_3 | reg_act_regs_data_2_15_2_enexo_3 | reg_act_config_inst_counter_enexo_63
      | reg_act_regs_data_0_15_2_enexo_3 | reg_act_regs_data_1_15_2_enexo_3);
  assign ActUnit_RunInst_curr_inst_and_enex5 = ActUnit_RunInst_switch_lp_and_802_cse
      & is_start_sva & (reg_act_config_inst_regs_17_sva_dfm_6_enexo_64 | reg_act_config_inst_regs_1_sva_dfm_5_enexo_64
      | reg_act_config_inst_counter_enexo_64);
  assign operator_32_8_true_AC_TRN_AC_WRAP_and_cse = ActUnit_RunInst_switch_lp_and_802_cse
      & and_dcpl_9 & (act_config_in_InstFetch_mux_tmp[7]) & (act_config_in_InstFetch_mux_tmp[4]);
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_and_cse = nv_scvector_cctor_nv_scvector_5_for_and_cse
      & and_dcpl_78;
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_and_17_cse = ActUnit_RunInst_switch_lp_and_812_cse
      & and_dcpl_78;
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_and_19_cse = nv_scvector_cctor_nv_scvector_5_for_and_3_cse
      & and_dcpl_78;
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_and_21_cse = nv_scvector_cctor_nv_scvector_5_for_and_5_cse
      & and_dcpl_78;
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_and_23_cse = nv_scvector_cctor_nv_scvector_5_for_and_7_cse
      & and_dcpl_78;
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_and_25_cse = nv_scvector_cctor_nv_scvector_5_for_and_9_cse
      & and_dcpl_78;
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_and_27_cse = nv_scvector_cctor_nv_scvector_5_for_and_11_cse
      & and_dcpl_78;
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_and_29_cse = nv_scvector_cctor_nv_scvector_5_for_and_13_cse
      & and_dcpl_78;
  assign or_71_cse = (~(is_start_sva & (act_config_in_InstFetch_mux_tmp[5]))) | (act_config_in_InstFetch_mux_tmp[7])
      | (act_config_in_InstFetch_mux_tmp[6]) | (act_config_in_InstFetch_mux_tmp[4])
      | (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]);
  assign mux_211_nl = MUX_s_1_2_2(mux_tmp_203, mux_tmp_197, fsm_output[1]);
  assign ActUnit_RunInst_switch_lp_and_808_cse = ActUnitRun_wen & (mux_211_nl | (fsm_output[4]));
  assign act_regs_data_and_404_ssc = (~ act_regs_data_0_0_sva_8_mx3c1) & and_dcpl_849;
  assign act_regs_data_and_405_ssc = act_regs_data_0_0_sva_8_mx3c1 & and_dcpl_849;
  assign act_regs_data_nor_1_nl = ~((and_dcpl_857 & and_dcpl_854) | act_regs_data_0_0_sva_8_mx3c1);
  assign reg_act_regs_data_0_0_1_rgt_nl = MUX1HOT_s_1_3_2(or_dcpl_449, (~ act_config_is_zero_first_sva_dfm_4),
      act_regs_data_nor_1_nl, {and_dcpl_557 , and_dcpl_852 , and_dcpl_849});
  assign act_regs_data_and_64_ssc = ActUnitRun_wen & (~(reg_act_regs_data_0_0_1_rgt_nl
      | (~ mux_215_itm)));
  assign act_regs_data_and_406_ssc = (~ act_regs_data_0_1_sva_8_mx3c1) & and_dcpl_849;
  assign act_regs_data_and_407_ssc = act_regs_data_0_1_sva_8_mx3c1 & and_dcpl_849;
  assign act_regs_data_or_1_nl = (and_dcpl_857 & and_dcpl_861) | act_regs_data_0_1_sva_8_mx3c1;
  assign reg_act_regs_data_0_1_1_rgt_nl = MUX1HOT_s_1_3_2((~ or_dcpl_456), act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_1_nl, {and_dcpl_557 , and_dcpl_852 , and_dcpl_849});
  assign act_regs_data_and_65_ssc = ActUnitRun_wen & ((reg_act_regs_data_0_1_1_rgt_nl
      & mux_215_itm) | and_dcpl_554);
  assign act_regs_data_and_408_ssc = (~ act_regs_data_0_10_sva_8_mx3c1) & and_dcpl_849;
  assign act_regs_data_and_409_ssc = act_regs_data_0_10_sva_8_mx3c1 & and_dcpl_849;
  assign act_regs_data_or_2_nl = (and_dcpl_867 & and_dcpl_865) | act_regs_data_0_10_sva_8_mx3c1;
  assign reg_act_regs_data_0_10_1_rgt_nl = MUX1HOT_s_1_3_2((~ or_dcpl_462), act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_2_nl, {and_dcpl_557 , and_dcpl_852 , and_dcpl_849});
  assign act_regs_data_and_66_ssc = ActUnitRun_wen & ((reg_act_regs_data_0_10_1_rgt_nl
      & mux_215_itm) | and_dcpl_554);
  assign act_regs_data_and_410_ssc = (~ act_regs_data_0_11_sva_8_mx3c1) & and_dcpl_849;
  assign act_regs_data_and_411_ssc = act_regs_data_0_11_sva_8_mx3c1 & and_dcpl_849;
  assign act_regs_data_or_4_nl = (and_dcpl_867 & and_dcpl_871) | act_regs_data_0_11_sva_8_mx3c1;
  assign reg_act_regs_data_0_11_1_rgt_nl = MUX1HOT_s_1_3_2((~ or_dcpl_469), act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_4_nl, {and_dcpl_557 , and_dcpl_852 , and_dcpl_849});
  assign act_regs_data_and_67_ssc = ActUnitRun_wen & ((reg_act_regs_data_0_11_1_rgt_nl
      & mux_215_itm) | and_dcpl_554);
  assign act_regs_data_and_412_ssc = (~ act_regs_data_0_12_sva_8_mx3c1) & and_dcpl_849;
  assign act_regs_data_and_413_ssc = act_regs_data_0_12_sva_8_mx3c1 & and_dcpl_849;
  assign act_regs_data_or_6_nl = (and_dcpl_857 & and_dcpl_874) | act_regs_data_0_12_sva_8_mx3c1;
  assign reg_act_regs_data_0_12_1_rgt_nl = MUX1HOT_s_1_3_2((~ or_dcpl_474), act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_6_nl, {and_dcpl_557 , and_dcpl_852 , and_dcpl_849});
  assign act_regs_data_and_68_ssc = ActUnitRun_wen & ((reg_act_regs_data_0_12_1_rgt_nl
      & mux_215_itm) | and_dcpl_554);
  assign act_regs_data_and_414_ssc = (~ act_regs_data_0_13_sva_8_mx3c1) & and_dcpl_849;
  assign act_regs_data_and_415_ssc = act_regs_data_0_13_sva_8_mx3c1 & and_dcpl_849;
  assign act_regs_data_or_8_nl = (and_dcpl_857 & and_dcpl_877) | act_regs_data_0_13_sva_8_mx3c1;
  assign reg_act_regs_data_0_13_1_rgt_nl = MUX1HOT_s_1_3_2((~ or_dcpl_477), act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_8_nl, {and_dcpl_557 , and_dcpl_852 , and_dcpl_849});
  assign act_regs_data_and_69_ssc = ActUnitRun_wen & ((reg_act_regs_data_0_13_1_rgt_nl
      & mux_215_itm) | and_dcpl_554);
  assign act_regs_data_and_416_ssc = (~ act_regs_data_0_14_sva_8_mx3c1) & and_dcpl_849;
  assign act_regs_data_and_417_ssc = act_regs_data_0_14_sva_8_mx3c1 & and_dcpl_849;
  assign act_regs_data_or_10_nl = (and_dcpl_867 & and_dcpl_874) | act_regs_data_0_14_sva_8_mx3c1;
  assign reg_act_regs_data_0_14_1_rgt_nl = MUX1HOT_s_1_3_2((~ or_dcpl_480), act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_10_nl, {and_dcpl_557 , and_dcpl_852 , and_dcpl_849});
  assign act_regs_data_and_70_ssc = ActUnitRun_wen & ((reg_act_regs_data_0_14_1_rgt_nl
      & mux_215_itm) | and_dcpl_554);
  assign act_regs_data_and_418_ssc = (~ act_regs_data_0_15_sva_8_mx3c1) & and_dcpl_849;
  assign act_regs_data_and_419_ssc = act_regs_data_0_15_sva_8_mx3c1 & and_dcpl_849;
  assign act_regs_data_or_12_nl = (and_dcpl_867 & and_dcpl_877) | act_regs_data_0_15_sva_8_mx3c1;
  assign reg_act_regs_data_0_15_1_rgt_nl = MUX1HOT_s_1_3_2((~ or_dcpl_482), act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_12_nl, {and_dcpl_557 , and_dcpl_852 , and_dcpl_849});
  assign act_regs_data_and_71_ssc = ActUnitRun_wen & ((reg_act_regs_data_0_15_1_rgt_nl
      & mux_215_itm) | and_dcpl_554);
  assign act_regs_data_and_420_ssc = (~ act_regs_data_0_2_sva_8_mx3c1) & and_dcpl_849;
  assign act_regs_data_and_421_ssc = act_regs_data_0_2_sva_8_mx3c1 & and_dcpl_849;
  assign act_regs_data_or_14_nl = (and_dcpl_867 & and_dcpl_854) | act_regs_data_0_2_sva_8_mx3c1;
  assign reg_act_regs_data_0_2_1_rgt_nl = MUX1HOT_s_1_3_2((~ or_dcpl_484), act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_14_nl, {and_dcpl_557 , and_dcpl_852 , and_dcpl_849});
  assign act_regs_data_and_72_ssc = ActUnitRun_wen & ((reg_act_regs_data_0_2_1_rgt_nl
      & mux_215_itm) | and_dcpl_554);
  assign act_regs_data_and_422_ssc = (~ act_regs_data_0_3_sva_8_mx3c1) & and_dcpl_849;
  assign act_regs_data_and_423_ssc = act_regs_data_0_3_sva_8_mx3c1 & and_dcpl_849;
  assign act_regs_data_or_16_nl = (and_dcpl_867 & and_dcpl_861) | act_regs_data_0_3_sva_8_mx3c1;
  assign reg_act_regs_data_0_3_1_rgt_nl = MUX1HOT_s_1_3_2((~ or_dcpl_487), act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_16_nl, {and_dcpl_557 , and_dcpl_852 , and_dcpl_849});
  assign act_regs_data_and_73_ssc = ActUnitRun_wen & ((reg_act_regs_data_0_3_1_rgt_nl
      & mux_215_itm) | and_dcpl_554);
  assign act_regs_data_and_424_ssc = (~ act_regs_data_0_4_sva_8_mx3c1) & and_dcpl_849;
  assign act_regs_data_and_425_ssc = act_regs_data_0_4_sva_8_mx3c1 & and_dcpl_849;
  assign act_regs_data_or_18_nl = (and_dcpl_857 & and_dcpl_888) | act_regs_data_0_4_sva_8_mx3c1;
  assign reg_act_regs_data_0_4_1_rgt_nl = MUX1HOT_s_1_3_2((~ or_dcpl_489), act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_18_nl, {and_dcpl_557 , and_dcpl_852 , and_dcpl_849});
  assign act_regs_data_and_74_ssc = ActUnitRun_wen & ((reg_act_regs_data_0_4_1_rgt_nl
      & mux_215_itm) | and_dcpl_554);
  assign act_regs_data_and_426_ssc = (~ act_regs_data_0_5_sva_8_mx3c1) & and_dcpl_849;
  assign act_regs_data_and_427_ssc = act_regs_data_0_5_sva_8_mx3c1 & and_dcpl_849;
  assign act_regs_data_or_20_nl = (and_dcpl_857 & and_dcpl_891) | act_regs_data_0_5_sva_8_mx3c1;
  assign reg_act_regs_data_0_5_1_rgt_nl = MUX1HOT_s_1_3_2((~ or_dcpl_492), act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_20_nl, {and_dcpl_557 , and_dcpl_852 , and_dcpl_849});
  assign act_regs_data_and_75_ssc = ActUnitRun_wen & ((reg_act_regs_data_0_5_1_rgt_nl
      & mux_215_itm) | and_dcpl_554);
  assign act_regs_data_and_428_ssc = (~ act_regs_data_0_6_sva_8_mx3c1) & and_dcpl_849;
  assign act_regs_data_and_429_ssc = act_regs_data_0_6_sva_8_mx3c1 & and_dcpl_849;
  assign act_regs_data_or_22_nl = (and_dcpl_867 & and_dcpl_888) | act_regs_data_0_6_sva_8_mx3c1;
  assign reg_act_regs_data_0_6_1_rgt_nl = MUX1HOT_s_1_3_2((~ or_dcpl_495), act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_22_nl, {and_dcpl_557 , and_dcpl_852 , and_dcpl_849});
  assign act_regs_data_and_76_ssc = ActUnitRun_wen & ((reg_act_regs_data_0_6_1_rgt_nl
      & mux_215_itm) | and_dcpl_554);
  assign act_regs_data_and_430_ssc = (~ act_regs_data_0_7_sva_8_mx3c1) & and_dcpl_849;
  assign act_regs_data_and_431_ssc = act_regs_data_0_7_sva_8_mx3c1 & and_dcpl_849;
  assign act_regs_data_or_24_nl = (and_dcpl_867 & and_dcpl_891) | act_regs_data_0_7_sva_8_mx3c1;
  assign reg_act_regs_data_0_7_1_rgt_nl = MUX1HOT_s_1_3_2((~ or_dcpl_497), act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_24_nl, {and_dcpl_557 , and_dcpl_852 , and_dcpl_849});
  assign act_regs_data_and_77_ssc = ActUnitRun_wen & ((reg_act_regs_data_0_7_1_rgt_nl
      & mux_215_itm) | and_dcpl_554);
  assign act_regs_data_and_432_ssc = (~ act_regs_data_0_8_sva_8_mx3c1) & and_dcpl_849;
  assign act_regs_data_and_433_ssc = act_regs_data_0_8_sva_8_mx3c1 & and_dcpl_849;
  assign act_regs_data_or_26_nl = (and_dcpl_857 & and_dcpl_865) | act_regs_data_0_8_sva_8_mx3c1;
  assign reg_act_regs_data_0_8_1_rgt_nl = MUX1HOT_s_1_3_2((~ or_dcpl_499), act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_26_nl, {and_dcpl_557 , and_dcpl_852 , and_dcpl_849});
  assign act_regs_data_and_78_ssc = ActUnitRun_wen & ((reg_act_regs_data_0_8_1_rgt_nl
      & mux_215_itm) | and_dcpl_554);
  assign ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_2_31 = MUX_s_1_64_2(act_regs_data_0_0_sva_dfm_2_31,
      act_regs_data_0_1_sva_dfm_2_31, act_regs_data_0_2_sva_dfm_2_31, act_regs_data_0_3_sva_dfm_2_31,
      act_regs_data_0_4_sva_dfm_2_31, act_regs_data_0_5_sva_dfm_2_31, act_regs_data_0_6_sva_dfm_2_31,
      act_regs_data_0_7_sva_dfm_2_31, act_regs_data_0_8_sva_dfm_2_31, act_regs_data_0_9_sva_dfm_2_31,
      act_regs_data_0_10_sva_dfm_2_31, act_regs_data_0_11_sva_dfm_2_31, act_regs_data_0_12_sva_dfm_2_31,
      act_regs_data_0_13_sva_dfm_2_31, act_regs_data_0_14_sva_dfm_2_31, act_regs_data_0_15_sva_dfm_2_31,
      act_regs_data_1_0_sva_dfm_2_31, act_regs_data_1_1_sva_dfm_2_31, act_regs_data_1_2_sva_dfm_2_31,
      act_regs_data_1_3_sva_dfm_2_31, act_regs_data_1_4_sva_dfm_2_31, act_regs_data_1_5_sva_dfm_2_31,
      act_regs_data_1_6_sva_dfm_2_31, act_regs_data_1_7_sva_dfm_2_31, act_regs_data_1_8_sva_dfm_2_31,
      act_regs_data_1_9_sva_dfm_2_31, act_regs_data_1_10_sva_dfm_2_31, act_regs_data_1_11_sva_dfm_2_31,
      act_regs_data_1_12_sva_dfm_2_31, act_regs_data_1_13_sva_dfm_2_31, act_regs_data_1_14_sva_dfm_2_31,
      act_regs_data_1_15_sva_dfm_2_31, act_regs_data_2_0_sva_dfm_2_31, act_regs_data_2_1_sva_dfm_2_31,
      act_regs_data_2_2_sva_dfm_2_31, act_regs_data_2_3_sva_dfm_2_31, act_regs_data_2_4_sva_dfm_2_31,
      act_regs_data_2_5_sva_dfm_2_31, act_regs_data_2_6_sva_dfm_2_31, act_regs_data_2_7_sva_dfm_2_31,
      act_regs_data_2_8_sva_dfm_2_31, act_regs_data_2_9_sva_dfm_2_31, act_regs_data_2_10_sva_dfm_2_31,
      act_regs_data_2_11_sva_dfm_2_31, act_regs_data_2_12_sva_dfm_2_31, act_regs_data_2_13_sva_dfm_2_31,
      act_regs_data_2_14_sva_dfm_2_31, act_regs_data_2_15_sva_dfm_2_31, act_regs_data_3_0_sva_dfm_2_31,
      act_regs_data_3_1_sva_dfm_2_31, act_regs_data_3_2_sva_dfm_2_31, act_regs_data_3_3_sva_dfm_2_31,
      act_regs_data_3_4_sva_dfm_2_31, act_regs_data_3_5_sva_dfm_2_31, act_regs_data_3_6_sva_dfm_2_31,
      act_regs_data_3_7_sva_dfm_2_31, act_regs_data_3_8_sva_dfm_2_31, act_regs_data_3_9_sva_dfm_2_31,
      act_regs_data_3_10_sva_dfm_2_31, act_regs_data_3_11_sva_dfm_2_31, act_regs_data_3_12_sva_dfm_2_31,
      act_regs_data_3_13_sva_dfm_2_31, act_regs_data_3_14_sva_dfm_2_31, act_regs_data_3_15_sva_dfm_2_31,
      {nvhls_get_slc_2U_NVUINT8_return_2_sva , ActUnit_PushOutput_if_for_i_4_0_sva_3_0});
  assign ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_2_30_0 = MUX_v_31_64_2(act_regs_data_0_0_sva_dfm_2_30_0,
      act_regs_data_0_1_sva_dfm_2_30_0, act_regs_data_0_2_sva_dfm_2_30_0, act_regs_data_0_3_sva_dfm_2_30_0,
      act_regs_data_0_4_sva_dfm_2_30_0, act_regs_data_0_5_sva_dfm_2_30_0, act_regs_data_0_6_sva_dfm_2_30_0,
      act_regs_data_0_7_sva_dfm_2_30_0, act_regs_data_0_8_sva_dfm_2_30_0, act_regs_data_0_9_sva_dfm_2_30_0,
      act_regs_data_0_10_sva_dfm_2_30_0, act_regs_data_0_11_sva_dfm_2_30_0, act_regs_data_0_12_sva_dfm_2_30_0,
      act_regs_data_0_13_sva_dfm_2_30_0, act_regs_data_0_14_sva_dfm_2_30_0, act_regs_data_0_15_sva_dfm_2_30_0,
      act_regs_data_1_0_sva_dfm_2_30_0, act_regs_data_1_1_sva_dfm_2_30_0, act_regs_data_1_2_sva_dfm_2_30_0,
      act_regs_data_1_3_sva_dfm_2_30_0, act_regs_data_1_4_sva_dfm_2_30_0, act_regs_data_1_5_sva_dfm_2_30_0,
      act_regs_data_1_6_sva_dfm_2_30_0, act_regs_data_1_7_sva_dfm_2_30_0, act_regs_data_1_8_sva_dfm_2_30_0,
      act_regs_data_1_9_sva_dfm_2_30_0, act_regs_data_1_10_sva_dfm_2_30_0, act_regs_data_1_11_sva_dfm_2_30_0,
      act_regs_data_1_12_sva_dfm_2_30_0, act_regs_data_1_13_sva_dfm_2_30_0, act_regs_data_1_14_sva_dfm_2_30_0,
      act_regs_data_1_15_sva_dfm_2_30_0, act_regs_data_2_0_sva_dfm_2_30_0, act_regs_data_2_1_sva_dfm_2_30_0,
      act_regs_data_2_2_sva_dfm_2_30_0, act_regs_data_2_3_sva_dfm_2_30_0, act_regs_data_2_4_sva_dfm_2_30_0,
      act_regs_data_2_5_sva_dfm_2_30_0, act_regs_data_2_6_sva_dfm_2_30_0, act_regs_data_2_7_sva_dfm_2_30_0,
      act_regs_data_2_8_sva_dfm_2_30_0, act_regs_data_2_9_sva_dfm_2_30_0, act_regs_data_2_10_sva_dfm_2_30_0,
      act_regs_data_2_11_sva_dfm_2_30_0, act_regs_data_2_12_sva_dfm_2_30_0, act_regs_data_2_13_sva_dfm_2_30_0,
      act_regs_data_2_14_sva_dfm_2_30_0, act_regs_data_2_15_sva_dfm_2_30_0, act_regs_data_3_0_sva_dfm_2_30_0,
      act_regs_data_3_1_sva_dfm_2_30_0, act_regs_data_3_2_sva_dfm_2_30_0, act_regs_data_3_3_sva_dfm_2_30_0,
      act_regs_data_3_4_sva_dfm_2_30_0, act_regs_data_3_5_sva_dfm_2_30_0, act_regs_data_3_6_sva_dfm_2_30_0,
      act_regs_data_3_7_sva_dfm_2_30_0, act_regs_data_3_8_sva_dfm_2_30_0, act_regs_data_3_9_sva_dfm_2_30_0,
      act_regs_data_3_10_sva_dfm_2_30_0, act_regs_data_3_11_sva_dfm_2_30_0, act_regs_data_3_12_sva_dfm_2_30_0,
      act_regs_data_3_13_sva_dfm_2_30_0, act_regs_data_3_14_sva_dfm_2_30_0, act_regs_data_3_15_sva_dfm_2_30_0,
      {nvhls_get_slc_2U_NVUINT8_return_2_sva , ActUnit_PushOutput_if_for_i_4_0_sva_3_0});
  assign ActUnit_RunInst_case_2_for_and_27_seb = ActUnit_PushOutput_if_for_and_stg_2_7_sva_1
      & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign nor_734_cse = ~((fsm_output[3:2]!=2'b00));
  assign or_1071_cse = (fsm_output[0]) | (fsm_output[2]);
  assign or_996_tmp = (ActUnit_DecodeAxiRead_unequal_tmp_1 & and_dcpl_906) | and_dcpl_908;
  assign act_mem_banks_read_for_and_cse = ActUnitRun_wen & (~ mux_tmp_55);
  assign mux_218_nl = MUX_s_1_2_2(nor_734_cse, or_1097_cse, fsm_output[4]);
  assign rva_out_reg_data_and_62_cse = ActUnitRun_wen & mux_218_nl & or_tmp_68;
  assign while_and_203_cse = (~ and_dcpl_916) & while_asn_1335;
  assign while_and_204_cse = and_dcpl_916 & while_asn_1335;
  assign mux_219_nl = MUX_s_1_2_2(nor_734_cse, mux_tmp_196, or_992_cse);
  assign ActUnit_RunInst_case_3_act_port_reg_data_and_cse = ActUnitRun_wen & (mux_219_nl
      | (fsm_output[4]));
  assign or_829_nl = and_1104_cse | (fsm_output[3:2]!=2'b00);
  assign mux_220_nl = MUX_s_1_2_2(nor_734_cse, or_829_nl, fsm_output[4]);
  assign act_config_output_counter_and_1_cse = ActUnitRun_wen & mux_220_nl;
  assign act_regs_data_and_284_cse = ActUnitRun_wen & and_dcpl_849 & and_dcpl_370
      & (~ act_config_is_zero_first_sva_dfm_4) & (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]);
  assign or_832_ssc = or_dcpl_504 | or_dcpl_478;
  assign or_833_ssc = or_dcpl_504 | or_dcpl_475;
  assign or_836_ssc = or_dcpl_508 | or_dcpl_478;
  assign or_837_ssc = or_dcpl_508 | or_dcpl_475;
  assign or_838_ssc = or_dcpl_504 | or_dcpl_471;
  assign or_839_ssc = or_dcpl_504 | or_dcpl_464;
  assign or_840_ssc = or_dcpl_508 | or_dcpl_471;
  assign or_841_ssc = or_dcpl_508 | or_dcpl_464;
  assign or_842_ssc = or_dcpl_504 | or_dcpl_493;
  assign or_843_ssc = or_dcpl_504 | or_dcpl_490;
  assign or_844_ssc = or_dcpl_508 | or_dcpl_493;
  assign or_845_ssc = or_dcpl_508 | or_dcpl_490;
  assign or_846_ssc = or_dcpl_504 | or_dcpl_458;
  assign or_847_ssc = or_dcpl_504 | or_dcpl_451;
  assign or_848_ssc = or_dcpl_508 | or_dcpl_458;
  assign act_regs_data_and_434_ssc = (~ act_regs_data_3_0_sva_8_mx2c1) & and_dcpl_849;
  assign act_regs_data_and_435_ssc = act_regs_data_3_0_sva_8_mx2c1 & and_dcpl_849;
  assign act_regs_data_or_126_nl = (and_dcpl_856 & (nvhls_get_slc_2U_NVUINT8_return_3_sva==2'b11)
      & and_dcpl_854) | act_regs_data_3_0_sva_8_mx2c1;
  assign act_regs_data_mux_128_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_126_nl, and_dcpl_849);
  assign act_regs_data_and_94_ssc = ActUnitRun_wen & act_regs_data_mux_128_nl & mux_215_itm;
  assign act_regs_data_and_436_ssc = (~ act_regs_data_2_15_sva_8_mx2c1) & and_dcpl_849;
  assign act_regs_data_and_437_ssc = act_regs_data_2_15_sva_8_mx2c1 & and_dcpl_849;
  assign act_regs_data_or_127_nl = (and_dcpl_924 & and_dcpl_877) | act_regs_data_2_15_sva_8_mx2c1;
  assign act_regs_data_mux_129_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_127_nl, and_dcpl_849);
  assign act_regs_data_and_95_ssc = ActUnitRun_wen & act_regs_data_mux_129_nl & mux_215_itm;
  assign act_regs_data_and_438_ssc = (~ act_regs_data_2_14_sva_8_mx2c1) & and_dcpl_849;
  assign act_regs_data_and_439_ssc = act_regs_data_2_14_sva_8_mx2c1 & and_dcpl_849;
  assign act_regs_data_or_128_nl = (and_dcpl_924 & and_dcpl_874) | act_regs_data_2_14_sva_8_mx2c1;
  assign act_regs_data_mux_130_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_128_nl, and_dcpl_849);
  assign act_regs_data_and_96_ssc = ActUnitRun_wen & act_regs_data_mux_130_nl & mux_215_itm;
  assign act_regs_data_and_440_ssc = (~ act_regs_data_2_13_sva_8_mx2c1) & and_dcpl_849;
  assign act_regs_data_and_441_ssc = act_regs_data_2_13_sva_8_mx2c1 & and_dcpl_849;
  assign act_regs_data_or_129_nl = (and_dcpl_929 & and_dcpl_877) | act_regs_data_2_13_sva_8_mx2c1;
  assign act_regs_data_mux_131_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_129_nl, and_dcpl_849);
  assign act_regs_data_and_97_ssc = ActUnitRun_wen & act_regs_data_mux_131_nl & mux_215_itm;
  assign act_regs_data_and_442_ssc = (~ act_regs_data_2_12_sva_8_mx2c1) & and_dcpl_849;
  assign act_regs_data_and_443_ssc = act_regs_data_2_12_sva_8_mx2c1 & and_dcpl_849;
  assign act_regs_data_or_130_nl = (and_dcpl_929 & and_dcpl_874) | act_regs_data_2_12_sva_8_mx2c1;
  assign act_regs_data_mux_132_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_130_nl, and_dcpl_849);
  assign act_regs_data_and_98_ssc = ActUnitRun_wen & act_regs_data_mux_132_nl & mux_215_itm;
  assign act_regs_data_and_444_ssc = (~ act_regs_data_2_11_sva_8_mx2c1) & and_dcpl_849;
  assign act_regs_data_and_445_ssc = act_regs_data_2_11_sva_8_mx2c1 & and_dcpl_849;
  assign act_regs_data_or_131_nl = (and_dcpl_924 & and_dcpl_871) | act_regs_data_2_11_sva_8_mx2c1;
  assign act_regs_data_mux_133_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_131_nl, and_dcpl_849);
  assign act_regs_data_and_99_ssc = ActUnitRun_wen & act_regs_data_mux_133_nl & mux_215_itm;
  assign act_regs_data_and_446_ssc = (~ act_regs_data_2_10_sva_8_mx2c1) & and_dcpl_849;
  assign act_regs_data_and_447_ssc = act_regs_data_2_10_sva_8_mx2c1 & and_dcpl_849;
  assign act_regs_data_or_132_nl = (and_dcpl_924 & and_dcpl_865) | act_regs_data_2_10_sva_8_mx2c1;
  assign act_regs_data_mux_134_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_132_nl, and_dcpl_849);
  assign act_regs_data_and_100_ssc = ActUnitRun_wen & act_regs_data_mux_134_nl &
      mux_215_itm;
  assign act_regs_data_and_448_ssc = (~ act_regs_data_2_9_sva_8_mx2c1) & and_dcpl_849;
  assign act_regs_data_and_449_ssc = act_regs_data_2_9_sva_8_mx2c1 & and_dcpl_849;
  assign act_regs_data_or_133_nl = (and_dcpl_929 & and_dcpl_871) | act_regs_data_2_9_sva_8_mx2c1;
  assign act_regs_data_mux_135_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_133_nl, and_dcpl_849);
  assign act_regs_data_and_101_ssc = ActUnitRun_wen & act_regs_data_mux_135_nl &
      mux_215_itm;
  assign act_regs_data_and_450_ssc = (~ act_regs_data_2_8_sva_8_mx2c1) & and_dcpl_849;
  assign act_regs_data_and_451_ssc = act_regs_data_2_8_sva_8_mx2c1 & and_dcpl_849;
  assign act_regs_data_or_134_nl = (and_dcpl_929 & and_dcpl_865) | act_regs_data_2_8_sva_8_mx2c1;
  assign act_regs_data_mux_136_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_134_nl, and_dcpl_849);
  assign act_regs_data_and_102_ssc = ActUnitRun_wen & act_regs_data_mux_136_nl &
      mux_215_itm;
  assign act_regs_data_and_452_ssc = (~ act_regs_data_2_7_sva_8_mx2c1) & and_dcpl_849;
  assign act_regs_data_and_453_ssc = act_regs_data_2_7_sva_8_mx2c1 & and_dcpl_849;
  assign act_regs_data_or_135_nl = (and_dcpl_924 & and_dcpl_891) | act_regs_data_2_7_sva_8_mx2c1;
  assign act_regs_data_mux_137_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_135_nl, and_dcpl_849);
  assign act_regs_data_and_103_ssc = ActUnitRun_wen & act_regs_data_mux_137_nl &
      mux_215_itm;
  assign act_regs_data_and_454_ssc = (~ act_regs_data_2_6_sva_8_mx2c1) & and_dcpl_849;
  assign act_regs_data_and_455_ssc = act_regs_data_2_6_sva_8_mx2c1 & and_dcpl_849;
  assign act_regs_data_or_136_nl = (and_dcpl_924 & and_dcpl_888) | act_regs_data_2_6_sva_8_mx2c1;
  assign act_regs_data_mux_138_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_136_nl, and_dcpl_849);
  assign act_regs_data_and_104_ssc = ActUnitRun_wen & act_regs_data_mux_138_nl &
      mux_215_itm;
  assign act_regs_data_and_456_ssc = (~ act_regs_data_2_5_sva_8_mx2c1) & and_dcpl_849;
  assign act_regs_data_and_457_ssc = act_regs_data_2_5_sva_8_mx2c1 & and_dcpl_849;
  assign act_regs_data_or_137_nl = (and_dcpl_929 & and_dcpl_891) | act_regs_data_2_5_sva_8_mx2c1;
  assign act_regs_data_mux_139_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_137_nl, and_dcpl_849);
  assign act_regs_data_and_105_ssc = ActUnitRun_wen & act_regs_data_mux_139_nl &
      mux_215_itm;
  assign act_regs_data_and_458_ssc = (~ act_regs_data_2_4_sva_8_mx2c1) & and_dcpl_849;
  assign act_regs_data_and_459_ssc = act_regs_data_2_4_sva_8_mx2c1 & and_dcpl_849;
  assign act_regs_data_or_138_nl = (and_dcpl_929 & and_dcpl_888) | act_regs_data_2_4_sva_8_mx2c1;
  assign act_regs_data_mux_140_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_138_nl, and_dcpl_849);
  assign act_regs_data_and_106_ssc = ActUnitRun_wen & act_regs_data_mux_140_nl &
      mux_215_itm;
  assign act_regs_data_and_460_ssc = (~ act_regs_data_2_3_sva_8_mx2c1) & and_dcpl_849;
  assign act_regs_data_and_461_ssc = act_regs_data_2_3_sva_8_mx2c1 & and_dcpl_849;
  assign act_regs_data_or_139_nl = (and_dcpl_924 & and_dcpl_861) | act_regs_data_2_3_sva_8_mx2c1;
  assign act_regs_data_mux_141_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_139_nl, and_dcpl_849);
  assign act_regs_data_and_107_ssc = ActUnitRun_wen & act_regs_data_mux_141_nl &
      mux_215_itm;
  assign act_regs_data_and_462_ssc = (~ act_regs_data_2_2_sva_8_mx2c1) & and_dcpl_849;
  assign act_regs_data_and_463_ssc = act_regs_data_2_2_sva_8_mx2c1 & and_dcpl_849;
  assign act_regs_data_or_140_nl = (and_dcpl_924 & and_dcpl_854) | act_regs_data_2_2_sva_8_mx2c1;
  assign act_regs_data_mux_142_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_140_nl, and_dcpl_849);
  assign act_regs_data_and_108_ssc = ActUnitRun_wen & act_regs_data_mux_142_nl &
      mux_215_itm;
  assign act_regs_data_and_464_ssc = (~ act_regs_data_2_1_sva_8_mx2c1) & and_dcpl_849;
  assign act_regs_data_and_465_ssc = act_regs_data_2_1_sva_8_mx2c1 & and_dcpl_849;
  assign act_regs_data_or_141_nl = (and_dcpl_929 & and_dcpl_861) | act_regs_data_2_1_sva_8_mx2c1;
  assign act_regs_data_mux_143_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_141_nl, and_dcpl_849);
  assign act_regs_data_and_109_ssc = ActUnitRun_wen & act_regs_data_mux_143_nl &
      mux_215_itm;
  assign act_regs_data_and_466_ssc = (~ act_regs_data_2_0_sva_8_mx2c1) & and_dcpl_849;
  assign act_regs_data_and_467_ssc = act_regs_data_2_0_sva_8_mx2c1 & and_dcpl_849;
  assign act_regs_data_or_142_nl = (and_dcpl_929 & and_dcpl_854) | act_regs_data_2_0_sva_8_mx2c1;
  assign act_regs_data_mux_144_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_142_nl, and_dcpl_849);
  assign act_regs_data_and_110_ssc = ActUnitRun_wen & act_regs_data_mux_144_nl &
      mux_215_itm;
  assign act_regs_data_and_468_ssc = (~ act_regs_data_1_15_sva_8_mx2c1) & and_dcpl_849;
  assign act_regs_data_and_469_ssc = act_regs_data_1_15_sva_8_mx2c1 & and_dcpl_849;
  assign act_regs_data_or_143_nl = (and_dcpl_959 & and_dcpl_877) | act_regs_data_1_15_sva_8_mx2c1;
  assign act_regs_data_mux_145_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_143_nl, and_dcpl_849);
  assign act_regs_data_and_111_ssc = ActUnitRun_wen & act_regs_data_mux_145_nl &
      mux_215_itm;
  assign act_regs_data_and_470_ssc = (~ act_regs_data_1_14_sva_8_mx2c1) & and_dcpl_849;
  assign act_regs_data_and_471_ssc = act_regs_data_1_14_sva_8_mx2c1 & and_dcpl_849;
  assign act_regs_data_or_144_nl = (and_dcpl_959 & and_dcpl_874) | act_regs_data_1_14_sva_8_mx2c1;
  assign act_regs_data_mux_146_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_144_nl, and_dcpl_849);
  assign act_regs_data_and_112_ssc = ActUnitRun_wen & act_regs_data_mux_146_nl &
      mux_215_itm;
  assign act_regs_data_and_472_ssc = (~ act_regs_data_1_13_sva_8_mx2c1) & and_dcpl_849;
  assign act_regs_data_and_473_ssc = act_regs_data_1_13_sva_8_mx2c1 & and_dcpl_849;
  assign act_regs_data_or_145_nl = (and_dcpl_964 & and_dcpl_877) | act_regs_data_1_13_sva_8_mx2c1;
  assign act_regs_data_mux_147_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_145_nl, and_dcpl_849);
  assign act_regs_data_and_113_ssc = ActUnitRun_wen & act_regs_data_mux_147_nl &
      mux_215_itm;
  assign act_regs_data_and_474_ssc = (~ act_regs_data_1_12_sva_8_mx2c1) & and_dcpl_849;
  assign act_regs_data_and_475_ssc = act_regs_data_1_12_sva_8_mx2c1 & and_dcpl_849;
  assign act_regs_data_or_146_nl = (and_dcpl_964 & and_dcpl_874) | act_regs_data_1_12_sva_8_mx2c1;
  assign act_regs_data_mux_148_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_146_nl, and_dcpl_849);
  assign act_regs_data_and_114_ssc = ActUnitRun_wen & act_regs_data_mux_148_nl &
      mux_215_itm;
  assign act_regs_data_and_476_ssc = (~ act_regs_data_1_11_sva_8_mx2c1) & and_dcpl_849;
  assign act_regs_data_and_477_ssc = act_regs_data_1_11_sva_8_mx2c1 & and_dcpl_849;
  assign act_regs_data_or_147_nl = (and_dcpl_959 & and_dcpl_871) | act_regs_data_1_11_sva_8_mx2c1;
  assign act_regs_data_mux_149_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_147_nl, and_dcpl_849);
  assign act_regs_data_and_115_ssc = ActUnitRun_wen & act_regs_data_mux_149_nl &
      mux_215_itm;
  assign act_regs_data_and_478_ssc = (~ act_regs_data_1_10_sva_8_mx2c1) & and_dcpl_849;
  assign act_regs_data_and_479_ssc = act_regs_data_1_10_sva_8_mx2c1 & and_dcpl_849;
  assign act_regs_data_or_148_nl = (and_dcpl_959 & and_dcpl_865) | act_regs_data_1_10_sva_8_mx2c1;
  assign act_regs_data_mux_150_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_148_nl, and_dcpl_849);
  assign act_regs_data_and_116_ssc = ActUnitRun_wen & act_regs_data_mux_150_nl &
      mux_215_itm;
  assign act_regs_data_and_480_ssc = (~ act_regs_data_1_9_sva_8_mx2c1) & and_dcpl_849;
  assign act_regs_data_and_481_ssc = act_regs_data_1_9_sva_8_mx2c1 & and_dcpl_849;
  assign act_regs_data_or_149_nl = (and_dcpl_964 & and_dcpl_871) | act_regs_data_1_9_sva_8_mx2c1;
  assign act_regs_data_mux_151_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_149_nl, and_dcpl_849);
  assign act_regs_data_and_117_ssc = ActUnitRun_wen & act_regs_data_mux_151_nl &
      mux_215_itm;
  assign act_regs_data_and_482_ssc = (~ act_regs_data_1_8_sva_8_mx2c1) & and_dcpl_849;
  assign act_regs_data_and_483_ssc = act_regs_data_1_8_sva_8_mx2c1 & and_dcpl_849;
  assign act_regs_data_or_150_nl = (and_dcpl_964 & and_dcpl_865) | act_regs_data_1_8_sva_8_mx2c1;
  assign act_regs_data_mux_152_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_150_nl, and_dcpl_849);
  assign act_regs_data_and_118_ssc = ActUnitRun_wen & act_regs_data_mux_152_nl &
      mux_215_itm;
  assign act_regs_data_and_484_ssc = (~ act_regs_data_1_7_sva_8_mx2c1) & and_dcpl_849;
  assign act_regs_data_and_485_ssc = act_regs_data_1_7_sva_8_mx2c1 & and_dcpl_849;
  assign act_regs_data_or_151_nl = (and_dcpl_959 & and_dcpl_891) | act_regs_data_1_7_sva_8_mx2c1;
  assign act_regs_data_mux_153_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_151_nl, and_dcpl_849);
  assign act_regs_data_and_119_ssc = ActUnitRun_wen & act_regs_data_mux_153_nl &
      mux_215_itm;
  assign act_regs_data_and_486_ssc = (~ act_regs_data_1_6_sva_8_mx2c1) & and_dcpl_849;
  assign act_regs_data_and_487_ssc = act_regs_data_1_6_sva_8_mx2c1 & and_dcpl_849;
  assign act_regs_data_or_152_nl = (and_dcpl_959 & and_dcpl_888) | act_regs_data_1_6_sva_8_mx2c1;
  assign act_regs_data_mux_154_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_152_nl, and_dcpl_849);
  assign act_regs_data_and_120_ssc = ActUnitRun_wen & act_regs_data_mux_154_nl &
      mux_215_itm;
  assign act_regs_data_and_488_ssc = (~ act_regs_data_1_5_sva_8_mx2c1) & and_dcpl_849;
  assign act_regs_data_and_489_ssc = act_regs_data_1_5_sva_8_mx2c1 & and_dcpl_849;
  assign act_regs_data_or_153_nl = (and_dcpl_964 & and_dcpl_891) | act_regs_data_1_5_sva_8_mx2c1;
  assign act_regs_data_mux_155_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_153_nl, and_dcpl_849);
  assign act_regs_data_and_121_ssc = ActUnitRun_wen & act_regs_data_mux_155_nl &
      mux_215_itm;
  assign act_regs_data_and_490_ssc = (~ act_regs_data_1_4_sva_8_mx2c1) & and_dcpl_849;
  assign act_regs_data_and_491_ssc = act_regs_data_1_4_sva_8_mx2c1 & and_dcpl_849;
  assign act_regs_data_or_154_nl = (and_dcpl_964 & and_dcpl_888) | act_regs_data_1_4_sva_8_mx2c1;
  assign act_regs_data_mux_156_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_154_nl, and_dcpl_849);
  assign act_regs_data_and_122_ssc = ActUnitRun_wen & act_regs_data_mux_156_nl &
      mux_215_itm;
  assign act_regs_data_and_492_ssc = (~ act_regs_data_1_3_sva_8_mx2c1) & and_dcpl_849;
  assign act_regs_data_and_493_ssc = act_regs_data_1_3_sva_8_mx2c1 & and_dcpl_849;
  assign act_regs_data_or_155_nl = (and_dcpl_959 & and_dcpl_861) | act_regs_data_1_3_sva_8_mx2c1;
  assign act_regs_data_mux_157_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_155_nl, and_dcpl_849);
  assign act_regs_data_and_123_ssc = ActUnitRun_wen & act_regs_data_mux_157_nl &
      mux_215_itm;
  assign act_regs_data_and_494_ssc = (~ act_regs_data_1_2_sva_8_mx2c1) & and_dcpl_849;
  assign act_regs_data_and_495_ssc = act_regs_data_1_2_sva_8_mx2c1 & and_dcpl_849;
  assign act_regs_data_or_156_nl = (and_dcpl_959 & and_dcpl_854) | act_regs_data_1_2_sva_8_mx2c1;
  assign act_regs_data_mux_158_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_156_nl, and_dcpl_849);
  assign act_regs_data_and_124_ssc = ActUnitRun_wen & act_regs_data_mux_158_nl &
      mux_215_itm;
  assign act_regs_data_and_496_ssc = (~ act_regs_data_1_1_sva_8_mx2c1) & and_dcpl_849;
  assign act_regs_data_and_497_ssc = act_regs_data_1_1_sva_8_mx2c1 & and_dcpl_849;
  assign act_regs_data_or_157_nl = (and_dcpl_964 & and_dcpl_861) | act_regs_data_1_1_sva_8_mx2c1;
  assign act_regs_data_mux_159_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_157_nl, and_dcpl_849);
  assign act_regs_data_and_125_ssc = ActUnitRun_wen & act_regs_data_mux_159_nl &
      mux_215_itm;
  assign act_regs_data_and_498_ssc = (~ act_regs_data_1_0_sva_8_mx2c1) & and_dcpl_849;
  assign act_regs_data_and_499_ssc = act_regs_data_1_0_sva_8_mx2c1 & and_dcpl_849;
  assign act_regs_data_or_158_nl = (and_dcpl_964 & and_dcpl_854) | act_regs_data_1_0_sva_8_mx2c1;
  assign act_regs_data_mux_160_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_158_nl, and_dcpl_849);
  assign act_regs_data_and_126_ssc = ActUnitRun_wen & act_regs_data_mux_160_nl &
      mux_215_itm;
  assign act_regs_data_and_500_ssc = (~ act_regs_data_0_9_sva_8_mx2c1) & and_dcpl_849;
  assign act_regs_data_and_501_ssc = act_regs_data_0_9_sva_8_mx2c1 & and_dcpl_849;
  assign act_regs_data_or_159_nl = (and_dcpl_857 & and_dcpl_871) | act_regs_data_0_9_sva_8_mx2c1;
  assign act_regs_data_mux_161_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_159_nl, and_dcpl_849);
  assign act_regs_data_and_127_ssc = ActUnitRun_wen & act_regs_data_mux_161_nl &
      mux_215_itm;
  assign nor_333_cse = ~((fsm_output[3:0]!=4'b0001));
  assign and_1108_cse = (fsm_output[2:1]==2'b11);
  assign and_1046_cse = or_992_cse & (fsm_output[2]);
  assign Silu_for_y_and_ssc = ActUnitRun_wen & ((~(and_1046_cse ^ (fsm_output[3])))
      | (fsm_output[4])) & and_dcpl_379;
  assign or_992_cse = (fsm_output[1:0]!=2'b00);
  assign nl_Silu_for_1_else_else_acc_nl = conv_s2s_27_30(ActUnit_RunInst_case_14_nv_scvector_cctor_data_0_sva_30_0[26:0])
      + conv_s2s_29_30(Tanh_for_1_else_else_mul_1_cmp_z[53:25]);
  assign Silu_for_1_else_else_acc_nl = nl_Silu_for_1_else_else_acc_nl[29:0];
  assign Silu_for_1_else_else_acc_itm_29_1 = readslicef_30_29_1(Silu_for_1_else_else_acc_nl);
  assign mux_224_nl = MUX_s_1_2_2(or_tmp_330, mux_tmp_196, fsm_output[1]);
  assign Silu_for_y_and_13_ssc = ActUnitRun_wen & (mux_224_nl | (fsm_output[4]))
      & and_dcpl_379;
  assign mux_225_nl = MUX_s_1_2_2(or_tmp_331, mux_tmp_196, fsm_output[0]);
  assign mux_226_nl = MUX_s_1_2_2(or_tmp_330, mux_225_nl, fsm_output[1]);
  assign Silu_for_y_and_15_ssc = ActUnitRun_wen & (mux_226_nl | (fsm_output[4]))
      & and_dcpl_379;
  assign Gelu_for_else_else_and_1_cse = ActUnitRun_wen & (~ and_dcpl_600);
  assign Silu_for_y_and_17_ssc = ActUnitRun_wen & (~(or_dcpl_290 & and_dcpl_1001))
      & and_dcpl_379;
  assign Silu_for_y_and_7_cse = ActUnitRun_wen & (~((or_992_cse ^ (fsm_output[2]))
      & and_dcpl_1001));
  assign Silu_for_y_and_19_ssc = Silu_for_y_and_7_cse & and_dcpl_379;
  assign and_1451_cse = (fsm_output[0]) & (fsm_output[2]);
  assign mux_329_cse = MUX_s_1_2_2((~ (fsm_output[2])), (fsm_output[2]), fsm_output[0]);
  assign mux_330_cse = MUX_s_1_2_2(mux_329_cse, and_1451_cse, fsm_output[1]);
  assign mux_328_cse = MUX_s_1_2_2((~ (fsm_output[2])), (fsm_output[2]), or_992_cse);
  assign Silu_for_y_and_8_ssc = ActUnitRun_wen & (~((~ mux_205_itm) & and_dcpl_1001))
      & and_dcpl_379;
  assign mux_336_cse = MUX_s_1_2_2((fsm_output[0]), (fsm_output[2]), fsm_output[1]);
  assign mux_337_cse = MUX_s_1_2_2((fsm_output[0]), and_1451_cse, fsm_output[1]);
  assign mux_232_nl = MUX_s_1_2_2(or_tmp_318, or_1077_cse, fsm_output[1]);
  assign Silu_for_y_and_20_ssc = ActUnitRun_wen & (~((~ mux_232_nl) & and_dcpl_1001))
      & and_dcpl_379;
  assign or_1077_cse = (~ (fsm_output[0])) | (fsm_output[2]);
  assign mux_342_cse = MUX_s_1_2_2(and_1451_cse, or_1077_cse, fsm_output[1]);
  assign mux_344_cse = MUX_s_1_2_2(and_1451_cse, mux_329_cse, fsm_output[1]);
  assign Silu_for_y_and_22_ssc = ActUnitRun_wen & (~ and_dcpl_1007) & and_dcpl_379;
  assign and_1249_cse = (fsm_output[0]) & or_dcpl_443;
  assign mux_350_cse = MUX_s_1_2_2(and_1108_cse, or_dcpl_443, fsm_output[0]);
  assign nl_Gelu_for_13_else_else_acc_nl = conv_s2s_26_29(nv_scvector_cctor_nv_scvector_6_for_13_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0])
      + conv_s2s_28_29(Tanh_for_1_else_else_mul_cmp_15_z[72:45]);
  assign Gelu_for_13_else_else_acc_nl = nl_Gelu_for_13_else_else_acc_nl[28:0];
  assign Gelu_for_13_else_else_acc_itm_28_1 = readslicef_29_28_1(Gelu_for_13_else_else_acc_nl);
  assign nl_Gelu_for_8_else_else_acc_nl = conv_s2s_26_29(nv_scvector_cctor_nv_scvector_6_for_8_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0])
      + conv_s2s_28_29(Tanh_for_1_else_else_mul_cmp_14_z[72:45]);
  assign Gelu_for_8_else_else_acc_nl = nl_Gelu_for_8_else_else_acc_nl[28:0];
  assign Gelu_for_8_else_else_acc_itm_28_1 = readslicef_29_28_1(Gelu_for_8_else_else_acc_nl);
  assign act_regs_data_and_299_cse = while_asn_1383 & (~ and_dcpl_849);
  assign act_regs_data_and_300_cse = while_asn_1385 & (~ and_dcpl_849);
  assign act_regs_data_and_301_cse = while_asn_1387 & (~ and_dcpl_849);
  assign act_regs_data_and_302_cse = while_asn_1389 & (~ and_dcpl_849);
  assign act_regs_data_and_303_cse = while_asn_1391 & (~ and_dcpl_849);
  assign act_regs_data_and_304_cse = while_asn_1393 & (~ and_dcpl_849);
  assign act_regs_data_and_305_cse = while_asn_1395 & (~ and_dcpl_849);
  assign nand_297_cse = ~((fsm_output[3:1]==3'b111));
  assign or_1097_cse = (fsm_output[3:1]!=3'b000);
  assign and_1460_nl = nand_297_cse & nand_tmp_13;
  assign mux_354_nl = MUX_s_1_2_2((fsm_output[0]), nand_tmp_13, or_1097_cse);
  assign mux_355_cse = MUX_s_1_2_2(and_1460_nl, mux_354_nl, fsm_output[4]);
  assign nand_298_cse = ~((fsm_output[0]) & nand_tmp_13);
  assign nor_736_cse = ~((fsm_output[4:1]!=4'b0110) | nand_298_cse);
  assign and_1485_cse = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3:2]==2'b11);
  assign and_1488_cse = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]) & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3])
      & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign act_regs_data_and_523_cse = while_asn_1369 & (~ and_dcpl_849);
  assign act_regs_data_and_524_cse = while_asn_1371 & (~ and_dcpl_849);
  assign act_regs_data_and_525_cse = while_asn_1373 & (~ and_dcpl_849);
  assign act_regs_data_and_526_cse = while_asn_1375 & (~ and_dcpl_849);
  assign act_regs_data_and_527_cse = while_asn_1377 & (~ and_dcpl_849);
  assign act_regs_data_and_528_cse = while_asn_1379 & (~ and_dcpl_849);
  assign act_regs_data_and_529_cse = while_asn_1381 & (~ and_dcpl_849);
  assign and_1496_nl = nand_297_cse & or_tmp_518;
  assign mux_410_nl = MUX_s_1_2_2((fsm_output[0]), or_tmp_518, or_1097_cse);
  assign mux_411_cse = MUX_s_1_2_2(and_1496_nl, mux_410_nl, fsm_output[4]);
  assign nand_338_cse = ~((fsm_output[0]) & or_tmp_518);
  assign nor_744_cse = ~((fsm_output[4:1]!=4'b0110) | nand_338_cse);
  assign act_regs_data_and_635_cse = while_asn_1355 & (~ and_dcpl_849);
  assign act_regs_data_and_636_cse = while_asn_1357 & (~ and_dcpl_849);
  assign act_regs_data_and_637_cse = while_asn_1359 & (~ and_dcpl_849);
  assign act_regs_data_and_638_cse = while_asn_1361 & (~ and_dcpl_849);
  assign act_regs_data_and_639_cse = while_asn_1363 & (~ and_dcpl_849);
  assign act_regs_data_and_640_cse = while_asn_1365 & (~ and_dcpl_849);
  assign act_regs_data_and_641_cse = while_asn_1367 & (~ and_dcpl_849);
  assign and_1532_nl = nand_297_cse & nand_tmp_45;
  assign mux_466_nl = MUX_s_1_2_2((fsm_output[0]), nand_tmp_45, or_1097_cse);
  assign mux_467_cse = MUX_s_1_2_2(and_1532_nl, mux_466_nl, fsm_output[4]);
  assign nand_378_cse = ~((fsm_output[0]) & nand_tmp_45);
  assign nor_752_cse = ~((fsm_output[4:1]!=4'b0110) | nand_378_cse);
  assign and_1876_cse = (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]) & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])
      & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]) & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign act_regs_data_and_747_cse = while_asn_1341 & (~ and_dcpl_849);
  assign act_regs_data_and_748_cse = while_asn_1343 & (~ and_dcpl_849);
  assign act_regs_data_and_749_cse = while_asn_1345 & (~ and_dcpl_849);
  assign act_regs_data_and_750_cse = while_asn_1347 & (~ and_dcpl_849);
  assign act_regs_data_and_751_cse = while_asn_1349 & (~ and_dcpl_849);
  assign act_regs_data_and_752_cse = while_asn_1351 & (~ and_dcpl_849);
  assign act_regs_data_and_753_cse = while_asn_1353 & (~ and_dcpl_849);
  assign and_1568_nl = nand_297_cse & or_tmp_726;
  assign mux_522_nl = MUX_s_1_2_2((fsm_output[0]), or_tmp_726, or_1097_cse);
  assign mux_523_cse = MUX_s_1_2_2(and_1568_nl, mux_522_nl, fsm_output[4]);
  assign nand_418_cse = ~((fsm_output[0]) & or_tmp_726);
  assign nor_760_cse = ~((fsm_output[4:1]!=4'b0110) | nand_418_cse);
  assign or_1488_cse = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]);
  assign nor_28_cse = ~((fsm_output[2:0]!=3'b001));
  assign and_1101_cse = (act_config_in_InstFetch_return_sva_7_2[3]) & (act_config_in_InstFetch_return_sva_7_2[5]);
  assign and_1103_cse = (act_config_in_InstFetch_return_sva_7_2[2]) & (act_config_in_InstFetch_return_sva_7_2[3])
      & (act_config_in_InstFetch_return_sva_7_2[5]);
  assign and_1104_cse = (fsm_output[1:0]==2'b11);
  assign ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_mx1
      = MUX_s_1_2_2(rva_in_PopNB_mioi_return_rsc_z_mxwt, ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva,
      is_start_sva);
  assign ActUnit_DecodeAxi_rva_in_reg_rw_sva_mx1 = MUX_s_1_2_2(rva_in_PopNB_mioi_data_rw_rsc_z_mxwt,
      ActUnit_DecodeAxi_rva_in_reg_rw_sva, is_start_sva);
  assign ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0 = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11:8]==4'b1001));
  assign ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_23_4_mx1_tmp_7_0
      = MUX_v_8_2_2((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7:0]), reg_ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_23_4_ftd_12,
      is_start_sva);
  assign act_mem_banks_read_read_data_lpi_1_dfm_1_31_0_mx1 = MUX_v_32_2_2(act_mem_banks_read_for_mux_15_itm,
      act_mem_banks_read_read_data_lpi_1_dfm_1_31_0, ActUnit_CheckStart_start_reg_sva);
  assign act_mem_banks_read_read_data_lpi_1_dfm_1_63_32_mx1 = MUX_v_32_2_2(act_mem_banks_read_for_mux_14_itm,
      act_mem_banks_read_read_data_lpi_1_dfm_1_63_32, ActUnit_CheckStart_start_reg_sva);
  assign act_mem_banks_read_read_data_lpi_1_dfm_1_95_64_mx1 = MUX_v_32_2_2(act_mem_banks_read_for_mux_13_itm,
      act_mem_banks_read_read_data_lpi_1_dfm_1_95_64, ActUnit_CheckStart_start_reg_sva);
  assign act_mem_banks_read_read_data_lpi_1_dfm_1_127_96_mx1 = MUX_v_32_2_2(act_mem_banks_read_for_mux_12_itm,
      act_mem_banks_read_read_data_lpi_1_dfm_1_127_96, ActUnit_CheckStart_start_reg_sva);
  assign act_mem_banks_read_read_data_lpi_1_dfm_1_159_128_mx1 = MUX_v_32_2_2(act_mem_banks_read_for_mux_11_itm,
      act_mem_banks_read_read_data_lpi_1_dfm_1_159_128, ActUnit_CheckStart_start_reg_sva);
  assign act_mem_banks_read_read_data_lpi_1_dfm_1_191_160_mx1 = MUX_v_32_2_2(act_mem_banks_read_for_mux_10_itm,
      act_mem_banks_read_read_data_lpi_1_dfm_1_191_160, ActUnit_CheckStart_start_reg_sva);
  assign act_mem_banks_read_read_data_lpi_1_dfm_1_223_192_mx1 = MUX_v_32_2_2(act_mem_banks_read_for_mux_9_itm,
      act_mem_banks_read_read_data_lpi_1_dfm_1_223_192, ActUnit_CheckStart_start_reg_sva);
  assign act_mem_banks_read_read_data_lpi_1_dfm_1_255_224_mx1 = MUX_v_32_2_2(act_mem_banks_read_for_mux_8_itm,
      act_mem_banks_read_read_data_lpi_1_dfm_1_255_224, ActUnit_CheckStart_start_reg_sva);
  assign act_mem_banks_read_read_data_lpi_1_dfm_1_287_256_mx1 = MUX_v_32_2_2(act_mem_banks_read_for_mux_7_itm,
      act_mem_banks_read_read_data_lpi_1_dfm_1_287_256, ActUnit_CheckStart_start_reg_sva);
  assign act_mem_banks_read_read_data_lpi_1_dfm_1_319_288_mx1 = MUX_v_32_2_2(act_mem_banks_read_for_mux_6_itm,
      act_mem_banks_read_read_data_lpi_1_dfm_1_319_288, ActUnit_CheckStart_start_reg_sva);
  assign act_mem_banks_read_read_data_lpi_1_dfm_1_351_320_mx1 = MUX_v_32_2_2(act_mem_banks_read_for_mux_5_itm,
      act_mem_banks_read_read_data_lpi_1_dfm_1_351_320, ActUnit_CheckStart_start_reg_sva);
  assign act_mem_banks_read_read_data_lpi_1_dfm_1_383_352_mx1 = MUX_v_32_2_2(act_mem_banks_read_for_mux_4_itm,
      act_mem_banks_read_read_data_lpi_1_dfm_1_383_352, ActUnit_CheckStart_start_reg_sva);
  assign act_mem_banks_read_read_data_lpi_1_dfm_1_415_384_mx1 = MUX_v_32_2_2(act_mem_banks_read_for_mux_3_itm,
      act_mem_banks_read_read_data_lpi_1_dfm_1_415_384, ActUnit_CheckStart_start_reg_sva);
  assign act_mem_banks_read_read_data_lpi_1_dfm_1_447_416_mx1 = MUX_v_32_2_2(act_mem_banks_read_for_mux_2_itm,
      act_mem_banks_read_read_data_lpi_1_dfm_1_447_416, ActUnit_CheckStart_start_reg_sva);
  assign act_mem_banks_read_read_data_lpi_1_dfm_1_479_448_mx1 = MUX_v_32_2_2(act_mem_banks_read_for_mux_1_itm,
      act_mem_banks_read_read_data_lpi_1_dfm_1_479_448, ActUnit_CheckStart_start_reg_sva);
  assign act_mem_banks_read_read_data_lpi_1_dfm_1_511_480_mx1 = MUX_v_32_2_2(act_mem_banks_read_for_mux_itm,
      act_mem_banks_read_read_data_lpi_1_dfm_1_511_480, ActUnit_CheckStart_start_reg_sva);
  assign nl_act_read_addrs_sva_2_mx0w0 = (act_config_output_counter_sva[4:0]) + act_config_buffer_addr_base_sva;
  assign act_read_addrs_sva_2_mx0w0 = nl_act_read_addrs_sva_2_mx0w0[4:0];
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_2_mx0w2 = act_read_addrs_lpi_1_dfm_7
      & ({{4{ActUnit_DecodeAxiRead_unequal_tmp_1}}, ActUnit_DecodeAxiRead_unequal_tmp_1})
      & ({{4{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt})
      & ({{4{rva_in_PopNB_mioi_return_rsc_z_mxwt}}, rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign Tanh_for_and_1_cse_sva_mx0w0 = (act_config_in_InstFetch_return_sva_7_2[1:0]==2'b01);
  assign ActUnit_PushOutput_if_for_and_stg_2_7_sva_1 = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2:0]==3'b111);
  assign Tanh_for_and_2_cse_sva_mx0w0 = (act_config_in_InstFetch_return_sva_7_2[1:0]==2'b11);
  assign ActUnit_RunInst_switch_lp_equal_tmp_1_mx0w0 = (act_config_in_InstFetch_mux_tmp[7:4]==4'b0010);
  assign ActUnit_RunInst_switch_lp_equal_tmp_2_mx0w0 = (act_config_in_InstFetch_mux_tmp[7:4]==4'b0011);
  assign ActUnit_RunInst_switch_lp_equal_tmp_3_mx0w0 = (act_config_in_InstFetch_mux_tmp[7:4]==4'b0100);
  assign ActUnit_RunInst_switch_lp_equal_tmp_4_mx0w0 = (act_config_in_InstFetch_mux_tmp[7:4]==4'b0111);
  assign ActUnit_RunInst_switch_lp_equal_tmp_5_mx0w0 = (act_config_in_InstFetch_mux_tmp[7:4]==4'b1011);
  assign ActUnit_RunInst_switch_lp_equal_tmp_6_mx0w0 = (act_config_in_InstFetch_mux_tmp[7:4]==4'b1100);
  assign ActUnit_RunInst_switch_lp_equal_tmp_7_mx0w0 = (act_config_in_InstFetch_mux_tmp[7:4]==4'b1110);
  assign ActUnit_RunInst_switch_lp_equal_tmp_8_mx0w0 = (act_config_in_InstFetch_mux_tmp[7:4]==4'b1111);
  assign ActUnit_RunInst_switch_lp_nor_nl = ~(ActUnit_RunInst_switch_lp_equal_tmp_9
      | ActUnit_RunInst_switch_lp_equal_tmp_1_mx0w0 | ActUnit_RunInst_switch_lp_equal_tmp_2_mx0w0
      | ActUnit_RunInst_switch_lp_equal_tmp_3_mx0w0 | ActUnit_RunInst_switch_lp_equal_tmp_4_mx0w0
      | ActUnit_RunInst_switch_lp_equal_tmp_5_mx0w0 | ActUnit_RunInst_switch_lp_equal_tmp_6_mx0w0
      | ActUnit_RunInst_switch_lp_equal_tmp_7_mx0w0 | ActUnit_RunInst_switch_lp_equal_tmp_8_mx0w0);
  assign ActUnit_RunInst_switch_lp_nor_tmp_mx0 = MUX_s_1_2_2(ActUnit_RunInst_switch_lp_nor_nl,
      ActUnit_RunInst_switch_lp_nor_tmp, or_dcpl_442);
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_less_15_tmp_1 = $signed({1'b0, 25'b1000000000000000000000000})
      < $signed(({ActUnit_RunInst_case_11_nv_scvector_cctor_data_0_sva_1_31 , ActUnit_RunInst_case_11_nv_scvector_cctor_data_0_sva_1_30_0}));
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_less_14_tmp_1 = $signed({1'b0, 25'b1000000000000000000000000})
      < $signed(({nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0}));
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_less_13_tmp_1 = $signed({1'b0, 25'b1000000000000000000000000})
      < $signed(({nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0}));
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_less_12_tmp_1 = $signed({1'b0, 25'b1000000000000000000000000})
      < $signed(({nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0}));
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_less_11_tmp_1 = $signed({1'b0, 25'b1000000000000000000000000})
      < $signed(({nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0}));
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_less_10_tmp_1 = $signed({1'b0, 25'b1000000000000000000000000})
      < $signed(({nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0}));
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_less_9_tmp_1 = $signed({1'b0, 25'b1000000000000000000000000})
      < $signed(({nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0}));
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_less_8_tmp_1 = $signed({1'b0, 25'b1000000000000000000000000})
      < $signed(({nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0}));
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_less_7_tmp_1 = $signed({1'b0, 25'b1000000000000000000000000})
      < $signed(({nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0}));
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_less_6_tmp_1 = $signed({1'b0, 25'b1000000000000000000000000})
      < $signed(({nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0}));
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_less_5_tmp_1 = $signed({1'b0, 25'b1000000000000000000000000})
      < $signed(({nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0}));
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_less_4_tmp_1 = $signed({1'b0, 25'b1000000000000000000000000})
      < $signed(({nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0}));
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_less_3_tmp_1 = $signed({1'b0, 25'b1000000000000000000000000})
      < $signed(({nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0}));
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_less_2_tmp_1 = $signed({1'b0, 25'b1000000000000000000000000})
      < $signed(({nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0}));
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_less_1_tmp_1 = $signed({1'b0, 25'b1000000000000000000000000})
      < $signed(({nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0}));
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_less_tmp_1 = $signed({1'b0, 25'b1000000000000000000000000})
      < $signed(({nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0}));
  assign nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      = MUX_s_1_4_2(act_regs_data_0_2_sva_31, act_regs_data_1_2_sva_31, act_regs_data_2_2_sva_31,
      act_regs_data_3_2_sva_31, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0
      = MUX_v_31_4_2(act_regs_data_0_2_sva_30_0, act_regs_data_1_2_sva_30_0, act_regs_data_2_2_sva_30_0,
      act_regs_data_3_2_sva_30_0, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      = MUX_s_1_4_2(act_regs_data_0_3_sva_31, act_regs_data_1_3_sva_31, act_regs_data_2_3_sva_31,
      act_regs_data_3_3_sva_31, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0
      = MUX_v_31_4_2(act_regs_data_0_3_sva_30_0, act_regs_data_1_3_sva_30_0, act_regs_data_2_3_sva_30_0,
      act_regs_data_3_3_sva_30_0, act_config_in_InstFetch_mux_tmp[3:2]);
  assign ActUnit_RunInst_case_11_nv_scvector_cctor_data_0_sva_1_31 = MUX_s_1_4_2(act_regs_data_0_0_sva_31,
      act_regs_data_1_0_sva_31, act_regs_data_2_0_sva_31, act_regs_data_3_0_sva_31,
      act_config_in_InstFetch_mux_tmp[3:2]);
  assign ActUnit_RunInst_case_11_nv_scvector_cctor_data_0_sva_1_30_0 = MUX_v_31_4_2(act_regs_data_0_0_sva_30_0,
      act_regs_data_1_0_sva_30_0, act_regs_data_2_0_sva_30_0, act_regs_data_3_0_sva_30_0,
      act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      = MUX_s_1_4_2(act_regs_data_0_1_sva_31, act_regs_data_1_1_sva_31, act_regs_data_2_1_sva_31,
      act_regs_data_3_1_sva_31, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0
      = MUX_v_31_4_2(act_regs_data_0_1_sva_30_0, act_regs_data_1_1_sva_30_0, act_regs_data_2_1_sva_30_0,
      act_regs_data_3_1_sva_30_0, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      = MUX_s_1_4_2(act_regs_data_0_4_sva_31, act_regs_data_1_4_sva_31, act_regs_data_2_4_sva_31,
      act_regs_data_3_4_sva_31, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0
      = MUX_v_31_4_2(act_regs_data_0_4_sva_30_0, act_regs_data_1_4_sva_30_0, act_regs_data_2_4_sva_30_0,
      act_regs_data_3_4_sva_30_0, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      = MUX_s_1_4_2(act_regs_data_0_5_sva_31, act_regs_data_1_5_sva_31, act_regs_data_2_5_sva_31,
      act_regs_data_3_5_sva_31, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0
      = MUX_v_31_4_2(act_regs_data_0_5_sva_30_0, act_regs_data_1_5_sva_30_0, act_regs_data_2_5_sva_30_0,
      act_regs_data_3_5_sva_30_0, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      = MUX_s_1_4_2(act_regs_data_0_6_sva_31, act_regs_data_1_6_sva_31, act_regs_data_2_6_sva_31,
      act_regs_data_3_6_sva_31, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0
      = MUX_v_31_4_2(act_regs_data_0_6_sva_30_0, act_regs_data_1_6_sva_30_0, act_regs_data_2_6_sva_30_0,
      act_regs_data_3_6_sva_30_0, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      = MUX_s_1_4_2(act_regs_data_0_7_sva_31, act_regs_data_1_7_sva_31, act_regs_data_2_7_sva_31,
      act_regs_data_3_7_sva_31, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0
      = MUX_v_31_4_2(act_regs_data_0_7_sva_30_0, act_regs_data_1_7_sva_30_0, act_regs_data_2_7_sva_30_0,
      act_regs_data_3_7_sva_30_0, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      = MUX_s_1_4_2(act_regs_data_0_8_sva_31, act_regs_data_1_8_sva_31, act_regs_data_2_8_sva_31,
      act_regs_data_3_8_sva_31, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0
      = MUX_v_31_4_2(act_regs_data_0_8_sva_30_0, act_regs_data_1_8_sva_30_0, act_regs_data_2_8_sva_30_0,
      act_regs_data_3_8_sva_30_0, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      = MUX_s_1_4_2(act_regs_data_0_9_sva_31, act_regs_data_1_9_sva_31, act_regs_data_2_9_sva_31,
      act_regs_data_3_9_sva_31, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0
      = MUX_v_31_4_2(act_regs_data_0_9_sva_30_0, act_regs_data_1_9_sva_30_0, act_regs_data_2_9_sva_30_0,
      act_regs_data_3_9_sva_30_0, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      = MUX_s_1_4_2(act_regs_data_0_10_sva_31, act_regs_data_1_10_sva_31, act_regs_data_2_10_sva_31,
      act_regs_data_3_10_sva_31, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0
      = MUX_v_31_4_2(act_regs_data_0_10_sva_30_0, act_regs_data_1_10_sva_30_0, act_regs_data_2_10_sva_30_0,
      act_regs_data_3_10_sva_30_0, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      = MUX_s_1_4_2(act_regs_data_0_11_sva_31, act_regs_data_1_11_sva_31, act_regs_data_2_11_sva_31,
      act_regs_data_3_11_sva_31, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0
      = MUX_v_31_4_2(act_regs_data_0_11_sva_30_0, act_regs_data_1_11_sva_30_0, act_regs_data_2_11_sva_30_0,
      act_regs_data_3_11_sva_30_0, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      = MUX_s_1_4_2(act_regs_data_0_12_sva_31, act_regs_data_1_12_sva_31, act_regs_data_2_12_sva_31,
      act_regs_data_3_12_sva_31, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0
      = MUX_v_31_4_2(act_regs_data_0_12_sva_30_0, act_regs_data_1_12_sva_30_0, act_regs_data_2_12_sva_30_0,
      act_regs_data_3_12_sva_30_0, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      = MUX_s_1_4_2(act_regs_data_0_13_sva_31, act_regs_data_1_13_sva_31, act_regs_data_2_13_sva_31,
      act_regs_data_3_13_sva_31, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0
      = MUX_v_31_4_2(act_regs_data_0_13_sva_30_0, act_regs_data_1_13_sva_30_0, act_regs_data_2_13_sva_30_0,
      act_regs_data_3_13_sva_30_0, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      = MUX_s_1_4_2(act_regs_data_0_14_sva_31, act_regs_data_1_14_sva_31, act_regs_data_2_14_sva_31,
      act_regs_data_3_14_sva_31, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0
      = MUX_v_31_4_2(act_regs_data_0_14_sva_30_0, act_regs_data_1_14_sva_30_0, act_regs_data_2_14_sva_30_0,
      act_regs_data_3_14_sva_30_0, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      = MUX_s_1_4_2(act_regs_data_0_15_sva_31, act_regs_data_1_15_sva_31, act_regs_data_2_15_sva_31,
      act_regs_data_3_15_sva_31, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0
      = MUX_v_31_4_2(act_regs_data_0_15_sva_30_0, act_regs_data_1_15_sva_30_0, act_regs_data_2_15_sva_30_0,
      act_regs_data_3_15_sva_30_0, act_config_in_InstFetch_mux_tmp[3:2]);
  assign act_config_in_InstFetch_mux_tmp = MUX_v_8_32_2(act_config_inst_regs_0_sva_dfm_5,
      act_config_inst_regs_1_sva_dfm_5, act_config_inst_regs_2_sva_dfm_5, act_config_inst_regs_3_sva_dfm_5,
      act_config_inst_regs_4_sva_dfm_5, act_config_inst_regs_5_sva_dfm_5, act_config_inst_regs_6_sva_dfm_5,
      act_config_inst_regs_7_sva_dfm_5, act_config_inst_regs_8_sva_dfm_5, act_config_inst_regs_9_sva_dfm_5,
      act_config_inst_regs_10_sva_dfm_5, act_config_inst_regs_11_sva_dfm_5, act_config_inst_regs_12_sva_dfm_5,
      act_config_inst_regs_13_sva_dfm_5, act_config_inst_regs_14_sva_dfm_5, act_config_inst_regs_15_sva_dfm_5,
      act_config_inst_regs_16_sva_dfm_6, act_config_inst_regs_17_sva_dfm_6, act_config_inst_regs_18_sva_dfm_6,
      act_config_inst_regs_19_sva_dfm_6, act_config_inst_regs_20_sva_dfm_6, act_config_inst_regs_21_sva_dfm_6,
      act_config_inst_regs_22_sva_dfm_6, act_config_inst_regs_23_sva_dfm_6, act_config_inst_regs_24_sva_dfm_6,
      act_config_inst_regs_25_sva_dfm_6, act_config_inst_regs_26_sva_dfm_6, act_config_inst_regs_27_sva_dfm_6,
      act_config_inst_regs_28_sva_dfm_6, act_config_inst_regs_29_sva_dfm_6, act_config_inst_regs_30_sva_dfm_6,
      act_config_inst_regs_31_sva_dfm_6, act_config_inst_counter_sva);
  assign operator_32_8_true_AC_TRN_AC_WRAP_3_less_tmp = $signed(({nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , (nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[30:24])}))
      < $signed(1'b1);
  assign operator_32_8_true_AC_TRN_AC_WRAP_3_less_1_tmp = $signed(({nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , (nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[30:24])}))
      < $signed(1'b1);
  assign operator_32_8_true_AC_TRN_AC_WRAP_3_less_2_tmp = $signed(({nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , (nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[30:24])}))
      < $signed(1'b1);
  assign operator_32_8_true_AC_TRN_AC_WRAP_3_less_3_tmp = $signed(({nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , (nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[30:24])}))
      < $signed(1'b1);
  assign operator_32_8_true_AC_TRN_AC_WRAP_3_less_4_tmp = $signed(({nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , (nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[30:24])}))
      < $signed(1'b1);
  assign operator_32_8_true_AC_TRN_AC_WRAP_3_less_5_tmp = $signed(({nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , (nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[30:24])}))
      < $signed(1'b1);
  assign operator_32_8_true_AC_TRN_AC_WRAP_3_less_6_tmp = $signed(({nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , (nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[30:24])}))
      < $signed(1'b1);
  assign operator_32_8_true_AC_TRN_AC_WRAP_3_less_7_tmp = $signed(({nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , (nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[30:24])}))
      < $signed(1'b1);
  assign operator_32_8_true_AC_TRN_AC_WRAP_3_less_8_tmp = $signed(({nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , (nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[30:24])}))
      < $signed(1'b1);
  assign operator_32_8_true_AC_TRN_AC_WRAP_3_less_9_tmp = $signed(({nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , (nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[30:24])}))
      < $signed(1'b1);
  assign operator_32_8_true_AC_TRN_AC_WRAP_3_less_10_tmp = $signed(({nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , (nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[30:24])}))
      < $signed(1'b1);
  assign operator_32_8_true_AC_TRN_AC_WRAP_3_less_11_tmp = $signed(({nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , (nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[30:24])}))
      < $signed(1'b1);
  assign operator_32_8_true_AC_TRN_AC_WRAP_3_less_12_tmp = $signed(({nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , (nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[30:24])}))
      < $signed(1'b1);
  assign operator_32_8_true_AC_TRN_AC_WRAP_3_less_13_tmp = $signed(({nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , (nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[30:24])}))
      < $signed(1'b1);
  assign operator_32_8_true_AC_TRN_AC_WRAP_3_less_14_tmp = $signed(({nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , (nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[30:24])}))
      < $signed(1'b1);
  assign operator_32_8_true_AC_TRN_AC_WRAP_3_less_15_tmp = $signed(({ActUnit_RunInst_case_11_nv_scvector_cctor_data_0_sva_1_31
      , (ActUnit_RunInst_case_11_nv_scvector_cctor_data_0_sva_1_30_0[30:24])})) <
      $signed(1'b1);
  assign operator_32_8_true_AC_TRN_AC_WRAP_1_less_15_tmp = $signed({1'b0, 26'b10000000000000000000000000})
      < $signed(({ActUnit_RunInst_case_11_nv_scvector_cctor_data_0_sva_1_31 , ActUnit_RunInst_case_11_nv_scvector_cctor_data_0_sva_1_30_0}));
  assign operator_32_8_true_AC_TRN_AC_WRAP_1_less_14_tmp = $signed({1'b0, 26'b10000000000000000000000000})
      < $signed(({nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0}));
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_less_12_tmp = $signed(({nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , (nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[30:25])}))
      < $signed(1'b1);
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_less_13_tmp = $signed(({nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , (nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[30:25])}))
      < $signed(1'b1);
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_less_14_tmp = $signed(({nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , (nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[30:25])}))
      < $signed(1'b1);
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_less_15_tmp = $signed(({ActUnit_RunInst_case_11_nv_scvector_cctor_data_0_sva_1_31
      , (ActUnit_RunInst_case_11_nv_scvector_cctor_data_0_sva_1_30_0[30:25])})) <
      $signed(1'b1);
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_less_10_tmp = $signed(({nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , (nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[30:25])}))
      < $signed(1'b1);
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_less_11_tmp = $signed(({nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , (nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[30:25])}))
      < $signed(1'b1);
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_less_8_tmp = $signed(({nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , (nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[30:25])}))
      < $signed(1'b1);
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_less_9_tmp = $signed(({nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , (nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[30:25])}))
      < $signed(1'b1);
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_less_6_tmp = $signed(({nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , (nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[30:25])}))
      < $signed(1'b1);
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_less_7_tmp = $signed(({nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , (nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[30:25])}))
      < $signed(1'b1);
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_less_4_tmp = $signed(({nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , (nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[30:25])}))
      < $signed(1'b1);
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_less_5_tmp = $signed(({nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , (nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[30:25])}))
      < $signed(1'b1);
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_less_2_tmp = $signed(({nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , (nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[30:25])}))
      < $signed(1'b1);
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_less_3_tmp = $signed(({nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , (nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[30:25])}))
      < $signed(1'b1);
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_less_tmp = $signed(({nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , (nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[30:25])}))
      < $signed(1'b1);
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_less_1_tmp = $signed(({nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
      , (nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[30:25])}))
      < $signed(1'b1);
  assign ActUnit_RunInst_switch_lp_equal_tmp_9 = (act_config_in_InstFetch_mux_tmp[7:4]==4'b0001);
  assign ActUnit_RunInst_switch_lp_and_16_tmp_mx0w1 = (act_config_in_InstFetch_return_sva_7_2[1:0]==2'b01)
      & act_port_PopNB_mioi_return_rsc_z_mxwt;
  assign ActUnit_RunInst_switch_lp_and_32_tmp_mx0w1 = (act_config_in_InstFetch_return_sva_7_2[1:0]==2'b10)
      & act_port_PopNB_mioi_return_rsc_z_mxwt;
  assign ActUnit_CheckStart_if_ActUnit_CheckStart_if_and_itm_1 = ActUnit_CheckStart_start_reg_sva
      & act_config_is_valid_sva & ActUnit_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva;
  assign act_config_InstIncr_if_equal_1_tmp = act_config_inst_counter_sva_dfm_3 ==
      (operator_6_false_acc_tmp[4:0]);
  assign act_config_InstIncr_act_config_InstIncr_if_and_svs_1 = act_config_InstIncr_if_equal_1_tmp
      & (operator_6_false_acc_tmp[6:5]==2'b00);
  assign ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_31 = MUX_s_1_64_2(act_regs_data_0_0_sva_31,
      act_regs_data_0_1_sva_31, act_regs_data_0_2_sva_31, act_regs_data_0_3_sva_31,
      act_regs_data_0_4_sva_31, act_regs_data_0_5_sva_31, act_regs_data_0_6_sva_31,
      act_regs_data_0_7_sva_31, act_regs_data_0_8_sva_31, act_regs_data_0_9_sva_31,
      act_regs_data_0_10_sva_31, act_regs_data_0_11_sva_31, act_regs_data_0_12_sva_31,
      act_regs_data_0_13_sva_31, act_regs_data_0_14_sva_31, act_regs_data_0_15_sva_31,
      act_regs_data_1_0_sva_31, act_regs_data_1_1_sva_31, act_regs_data_1_2_sva_31,
      act_regs_data_1_3_sva_31, act_regs_data_1_4_sva_31, act_regs_data_1_5_sva_31,
      act_regs_data_1_6_sva_31, act_regs_data_1_7_sva_31, act_regs_data_1_8_sva_31,
      act_regs_data_1_9_sva_31, act_regs_data_1_10_sva_31, act_regs_data_1_11_sva_31,
      act_regs_data_1_12_sva_31, act_regs_data_1_13_sva_31, act_regs_data_1_14_sva_31,
      act_regs_data_1_15_sva_31, act_regs_data_2_0_sva_31, act_regs_data_2_1_sva_31,
      act_regs_data_2_2_sva_31, act_regs_data_2_3_sva_31, act_regs_data_2_4_sva_31,
      act_regs_data_2_5_sva_31, act_regs_data_2_6_sva_31, act_regs_data_2_7_sva_31,
      act_regs_data_2_8_sva_31, act_regs_data_2_9_sva_31, act_regs_data_2_10_sva_31,
      act_regs_data_2_11_sva_31, act_regs_data_2_12_sva_31, act_regs_data_2_13_sva_31,
      act_regs_data_2_14_sva_31, act_regs_data_2_15_sva_31, act_regs_data_3_0_sva_31,
      act_regs_data_3_1_sva_31, act_regs_data_3_2_sva_31, act_regs_data_3_3_sva_31,
      act_regs_data_3_4_sva_31, act_regs_data_3_5_sva_31, act_regs_data_3_6_sva_31,
      act_regs_data_3_7_sva_31, act_regs_data_3_8_sva_31, act_regs_data_3_9_sva_31,
      act_regs_data_3_10_sva_31, act_regs_data_3_11_sva_31, act_regs_data_3_12_sva_31,
      act_regs_data_3_13_sva_31, act_regs_data_3_14_sva_31, act_regs_data_3_15_sva_31,
      {(act_config_in_InstFetch_return_sva_7_2[1:0]) , ActUnit_PushOutput_if_for_i_4_0_sva_3_0});
  assign ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_30_0 =
      MUX_v_31_64_2(act_regs_data_0_0_sva_30_0, act_regs_data_0_1_sva_30_0, act_regs_data_0_2_sva_30_0,
      act_regs_data_0_3_sva_30_0, act_regs_data_0_4_sva_30_0, act_regs_data_0_5_sva_30_0,
      act_regs_data_0_6_sva_30_0, act_regs_data_0_7_sva_30_0, act_regs_data_0_8_sva_30_0,
      act_regs_data_0_9_sva_30_0, act_regs_data_0_10_sva_30_0, act_regs_data_0_11_sva_30_0,
      act_regs_data_0_12_sva_30_0, act_regs_data_0_13_sva_30_0, act_regs_data_0_14_sva_30_0,
      act_regs_data_0_15_sva_30_0, act_regs_data_1_0_sva_30_0, act_regs_data_1_1_sva_30_0,
      act_regs_data_1_2_sva_30_0, act_regs_data_1_3_sva_30_0, act_regs_data_1_4_sva_30_0,
      act_regs_data_1_5_sva_30_0, act_regs_data_1_6_sva_30_0, act_regs_data_1_7_sva_30_0,
      act_regs_data_1_8_sva_30_0, act_regs_data_1_9_sva_30_0, act_regs_data_1_10_sva_30_0,
      act_regs_data_1_11_sva_30_0, act_regs_data_1_12_sva_30_0, act_regs_data_1_13_sva_30_0,
      act_regs_data_1_14_sva_30_0, act_regs_data_1_15_sva_30_0, act_regs_data_2_0_sva_30_0,
      act_regs_data_2_1_sva_30_0, act_regs_data_2_2_sva_30_0, act_regs_data_2_3_sva_30_0,
      act_regs_data_2_4_sva_30_0, act_regs_data_2_5_sva_30_0, act_regs_data_2_6_sva_30_0,
      act_regs_data_2_7_sva_30_0, act_regs_data_2_8_sva_30_0, act_regs_data_2_9_sva_30_0,
      act_regs_data_2_10_sva_30_0, act_regs_data_2_11_sva_30_0, act_regs_data_2_12_sva_30_0,
      act_regs_data_2_13_sva_30_0, act_regs_data_2_14_sva_30_0, act_regs_data_2_15_sva_30_0,
      act_regs_data_3_0_sva_30_0, act_regs_data_3_1_sva_30_0, act_regs_data_3_2_sva_30_0,
      act_regs_data_3_3_sva_30_0, act_regs_data_3_4_sva_30_0, act_regs_data_3_5_sva_30_0,
      act_regs_data_3_6_sva_30_0, act_regs_data_3_7_sva_30_0, act_regs_data_3_8_sva_30_0,
      act_regs_data_3_9_sva_30_0, act_regs_data_3_10_sva_30_0, act_regs_data_3_11_sva_30_0,
      act_regs_data_3_12_sva_30_0, act_regs_data_3_13_sva_30_0, act_regs_data_3_14_sva_30_0,
      act_regs_data_3_15_sva_30_0, {(act_config_in_InstFetch_return_sva_7_2[1:0])
      , ActUnit_PushOutput_if_for_i_4_0_sva_3_0});
  assign act_config_ActConfigRead_else_unequal_tmp_1 = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7:0]==8'b00000010));
  assign act_config_ActConfigRead_unequal_tmp_1 = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7:0]==8'b00000001));
  assign ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_2_tmp
      = ~(act_config_is_zero_first_sva | ActUnit_RunInst_switch_lp_and_32_tmp | ActUnit_RunInst_switch_lp_equal_tmp_2
      | ActUnit_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva
      | ActUnit_RunInst_switch_lp_equal_tmp_4 | ActUnit_RunInst_switch_lp_equal_tmp_5
      | ActUnit_RunInst_switch_lp_equal_tmp_6 | ActUnit_RunInst_switch_lp_equal_tmp_7
      | ActUnit_RunInst_switch_lp_equal_tmp_8 | ActUnit_RunInst_switch_lp_nor_tmp);
  assign ActUnit_DecodeAxiRead_unequal_tmp_1 = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11:8]==4'b1000));
  assign ActUnit_DecodeAxi_if_or_7_tmp_1 = ActUnit_DecodeAxiRead_unequal_tmp_1 |
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_6_nl = act_read_addrs_lpi_1_dfm_7
      & ({{4{ActUnit_DecodeAxiRead_unequal_tmp_1}}, ActUnit_DecodeAxiRead_unequal_tmp_1})
      & (signext_5_1(~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)) & ({{4{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_nl = ~(ActUnit_RunInst_switch_lp_and_32_tmp
      | ActUnit_RunInst_switch_lp_equal_tmp_2 | ActUnit_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva
      | ActUnit_RunInst_switch_lp_equal_tmp_4 | ActUnit_RunInst_switch_lp_equal_tmp_5
      | ActUnit_RunInst_switch_lp_equal_tmp_6 | ActUnit_RunInst_switch_lp_equal_tmp_7
      | ActUnit_RunInst_switch_lp_equal_tmp_8 | ActUnit_RunInst_switch_lp_nor_tmp);
  assign ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_and_18_nl = act_config_inst_counter_sva_dfm_3
      & (signext_5_1(~ act_config_is_zero_first_sva)) & (signext_5_1(ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_nl));
  assign while_mux_53_ssc_mx0 = MUX_v_5_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_6_nl,
      ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_and_18_nl, is_start_sva);
  assign while_and_88_tmp_1 = ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_mx1
      & (~ is_start_sva);
  assign ActUnit_DecodeAxiWrite_else_not_17_nl = ~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0;
  assign act_read_addrs_lpi_1_dfm_7 = MUX_v_5_2_2(5'b00000, (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4:0]),
      ActUnit_DecodeAxiWrite_else_not_17_nl);
  assign Tanh_for_nor_cse_sva_mx0w0 = ~((act_config_in_InstFetch_return_sva_7_2[1:0]!=2'b00));
  assign Tanh_for_and_cse_sva_mx0w0 = (act_config_in_InstFetch_return_sva_7_2[1:0]==2'b10);
  assign ActUnit_RunInst_switch_lp_and_48_tmp_mx0w0 = (act_config_in_InstFetch_return_sva_7_2[1:0]==2'b11)
      & act_port_PopNB_mioi_return_rsc_z_mxwt;
  assign ActUnit_RunInst_switch_lp_and_tmp_mx0w0 = Tanh_for_nor_cse_sva_mx0w0 & act_port_PopNB_mioi_return_rsc_z_mxwt;
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_7_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[31:0])
      & (signext_32_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{31{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{31{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{31{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_0_lpi_1_dfm_7 = MUX_v_32_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_7_nl,
      ({act_regs_data_0_0_sva_8_31 , act_regs_data_0_0_sva_8_30_0}), while_and_1_tmp);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_8_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[63:32])
      & (signext_32_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{31{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{31{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{31{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_1_lpi_1_dfm_7 = MUX_v_32_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_8_nl,
      ({act_regs_data_0_1_sva_8_31 , act_regs_data_0_1_sva_8_30_0}), while_and_1_tmp);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_9_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[95:64])
      & (signext_32_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{31{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{31{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{31{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_2_lpi_1_dfm_7 = MUX_v_32_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_9_nl,
      ({act_regs_data_0_15_sva_8_31 , act_regs_data_0_15_sva_8_30_0}), while_and_1_tmp);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_10_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[127:96])
      & (signext_32_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{31{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{31{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{31{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_3_lpi_1_dfm_7 = MUX_v_32_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_10_nl,
      ({act_regs_data_0_2_sva_8_31 , act_regs_data_0_2_sva_8_30_0}), while_and_1_tmp);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_11_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[159:128])
      & (signext_32_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{31{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{31{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{31{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_4_lpi_1_dfm_7 = MUX_v_32_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_11_nl,
      ({act_regs_data_0_3_sva_8_31 , act_regs_data_0_3_sva_8_30_0}), while_and_1_tmp);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_12_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[191:160])
      & (signext_32_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{31{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{31{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{31{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_5_lpi_1_dfm_7 = MUX_v_32_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_12_nl,
      ({act_regs_data_0_4_sva_8_31 , act_regs_data_0_4_sva_8_30_0}), while_and_1_tmp);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_13_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[223:192])
      & (signext_32_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{31{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{31{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{31{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_6_lpi_1_dfm_7 = MUX_v_32_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_13_nl,
      ({act_regs_data_0_5_sva_8_31 , act_regs_data_0_5_sva_8_30_0}), while_and_1_tmp);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_14_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[255:224])
      & (signext_32_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{31{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{31{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{31{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_7_lpi_1_dfm_7 = MUX_v_32_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_14_nl,
      ({act_regs_data_0_6_sva_8_31 , act_regs_data_0_6_sva_8_30_0}), while_and_1_tmp);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_15_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[287:256])
      & (signext_32_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{31{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{31{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{31{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_8_lpi_1_dfm_7 = MUX_v_32_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_15_nl,
      ({act_regs_data_0_7_sva_8_31 , act_regs_data_0_7_sva_8_30_0}), while_and_1_tmp);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_16_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[319:288])
      & (signext_32_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{31{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{31{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{31{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_9_lpi_1_dfm_7 = MUX_v_32_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_16_nl,
      ({act_regs_data_0_8_sva_8_31 , act_regs_data_0_8_sva_8_30_0}), while_and_1_tmp);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_17_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[351:320])
      & (signext_32_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{31{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{31{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{31{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_10_lpi_1_dfm_7 = MUX_v_32_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_17_nl,
      ({act_regs_data_0_10_sva_8_31 , act_regs_data_0_10_sva_8_30_0}), while_and_1_tmp);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_18_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[383:352])
      & (signext_32_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{31{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{31{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{31{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_11_lpi_1_dfm_7 = MUX_v_32_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_18_nl,
      ({act_regs_data_0_11_sva_8_31 , act_regs_data_0_11_sva_8_30_0}), while_and_1_tmp);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_19_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[415:384])
      & (signext_32_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{31{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{31{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{31{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_12_lpi_1_dfm_7 = MUX_v_32_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_19_nl,
      ({act_regs_data_0_12_sva_8_31 , act_regs_data_0_12_sva_8_30_0}), while_and_1_tmp);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_20_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[447:416])
      & (signext_32_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{31{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{31{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{31{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_13_lpi_1_dfm_7 = MUX_v_32_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_20_nl,
      ({act_regs_data_0_13_sva_8_31 , act_regs_data_0_13_sva_8_30_0}), while_and_1_tmp);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_21_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[479:448])
      & (signext_32_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{31{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{31{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{31{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_14_lpi_1_dfm_7 = MUX_v_32_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_21_nl,
      ({act_regs_data_0_14_sva_8_31 , act_regs_data_0_14_sva_8_30_0}), while_and_1_tmp);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_22_itm = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[511:480])
      & (signext_32_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{31{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{31{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{31{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign while_mux_32_nl = MUX_s_1_2_2((ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_22_itm[31]),
      ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_31, while_and_1_tmp);
  assign while_mux_395_nl = MUX_v_31_2_2((ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_22_itm[30:0]),
      ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_30_0, while_and_1_tmp);
  assign while_while_nand_nl = ~((~ ActUnit_RunInst_switch_lp_and_32_tmp) & is_start_sva);
  assign act_write_data_data_0_15_lpi_1_dfm_7 = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      ({while_mux_32_nl , while_mux_395_nl}), while_while_nand_nl);
  assign while_and_1_tmp = ActUnit_RunInst_switch_lp_and_32_tmp & is_start_sva;
  assign act_config_ActConfigRead_else_else_not_21 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7:0]==8'b00000011);
  assign while_asn_1331 = (~ while_and_88_tmp_1) | ActUnit_DecodeAxi_if_or_7_tmp_1;
  assign while_asn_1333 = (~(act_config_ActConfigRead_unequal_tmp_1 | ActUnit_DecodeAxi_if_or_7_tmp_1))
      & while_and_88_tmp_1;
  assign while_asn_1335 = act_config_ActConfigRead_unequal_tmp_1 & (~ ActUnit_DecodeAxi_if_or_7_tmp_1)
      & while_and_88_tmp_1;
  assign Gelu_for_y_lpi_1_dfm_2_31 = (z_out_28_1[27]) & (~ Tanh_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)
      & (~ Tanh_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs);
  assign Gelu_for_else_mux_15_nl = MUX_v_31_2_2(({{3{z_out_28_1[27]}}, z_out_28_1}),
      nv_scvector_cctor_nv_scvector_6_for_16_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0,
      Tanh_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
  assign operator_32_8_true_AC_TRN_AC_WRAP_3_not_31_nl = ~ Tanh_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs;
  assign Gelu_for_y_lpi_1_dfm_2_30_0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      Gelu_for_else_mux_15_nl, operator_32_8_true_AC_TRN_AC_WRAP_3_not_31_nl);
  assign Gelu_for_y_11_lpi_1_dfm_2_31 = (z_out_2_28_1[27]) & (~ Tanh_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)
      & (~ Tanh_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs);
  assign Gelu_for_else_mux_10_nl = MUX_v_31_2_2(({{3{z_out_2_28_1[27]}}, z_out_2_28_1}),
      nv_scvector_cctor_nv_scvector_6_for_11_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0,
      Tanh_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
  assign operator_32_8_true_AC_TRN_AC_WRAP_3_not_32_nl = ~ Tanh_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs;
  assign Gelu_for_y_11_lpi_1_dfm_2_30_0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      Gelu_for_else_mux_10_nl, operator_32_8_true_AC_TRN_AC_WRAP_3_not_32_nl);
  assign Gelu_for_y_10_lpi_1_dfm_2_31 = (z_out_1_28_1[27]) & (~ Tanh_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)
      & (~ Tanh_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs);
  assign Gelu_for_else_mux_9_nl = MUX_v_31_2_2(({{3{z_out_1_28_1[27]}}, z_out_1_28_1}),
      nv_scvector_cctor_nv_scvector_6_for_10_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0,
      Tanh_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
  assign operator_32_8_true_AC_TRN_AC_WRAP_3_not_33_nl = ~ Tanh_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs;
  assign Gelu_for_y_10_lpi_1_dfm_2_30_0 = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      Gelu_for_else_mux_9_nl, operator_32_8_true_AC_TRN_AC_WRAP_3_not_33_nl);
  assign while_asn_1341 = ~(is_start_sva & while_nor_48_itm);
  assign while_asn_1343 = ActUnit_RunInst_switch_lp_and_48_tmp & ActUnit_RunInst_switch_lp_equal_tmp_2
      & is_start_sva;
  assign while_asn_1345 = reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_2_cse
      & ActUnit_RunInst_switch_lp_equal_tmp_4 & is_start_sva;
  assign while_asn_1347 = reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_2_cse
      & ActUnit_RunInst_switch_lp_equal_tmp_5 & is_start_sva;
  assign while_asn_1349 = reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_2_cse
      & ActUnit_RunInst_switch_lp_equal_tmp_6 & is_start_sva;
  assign while_asn_1351 = reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_2_cse
      & ActUnit_RunInst_switch_lp_equal_tmp_7 & is_start_sva;
  assign while_asn_1353 = Gelu_for_and_2_cse_sva & ActUnit_RunInst_switch_lp_equal_tmp_8
      & is_start_sva;
  assign while_asn_1355 = ~(is_start_sva & while_nor_32_itm);
  assign while_asn_1357 = ActUnit_RunInst_switch_lp_and_32_tmp & ActUnit_RunInst_switch_lp_equal_tmp_2
      & is_start_sva;
  assign while_asn_1359 = reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_cse
      & ActUnit_RunInst_switch_lp_equal_tmp_4 & is_start_sva;
  assign while_asn_1361 = reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_cse
      & ActUnit_RunInst_switch_lp_equal_tmp_5 & is_start_sva;
  assign while_asn_1363 = reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_cse
      & ActUnit_RunInst_switch_lp_equal_tmp_6 & is_start_sva;
  assign while_asn_1365 = reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_cse
      & ActUnit_RunInst_switch_lp_equal_tmp_7 & is_start_sva;
  assign while_asn_1367 = reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_cse
      & ActUnit_RunInst_switch_lp_equal_tmp_8 & is_start_sva;
  assign while_asn_1369 = ~(is_start_sva & while_nor_16_itm);
  assign while_asn_1371 = ActUnit_RunInst_switch_lp_and_16_tmp & ActUnit_RunInst_switch_lp_equal_tmp_2
      & is_start_sva;
  assign while_asn_1373 = reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_1_cse
      & ActUnit_RunInst_switch_lp_equal_tmp_4 & is_start_sva;
  assign while_asn_1375 = reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_1_cse
      & ActUnit_RunInst_switch_lp_equal_tmp_5 & is_start_sva;
  assign while_asn_1377 = reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_1_cse
      & ActUnit_RunInst_switch_lp_equal_tmp_6 & is_start_sva;
  assign while_asn_1379 = reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_1_cse
      & ActUnit_RunInst_switch_lp_equal_tmp_7 & is_start_sva;
  assign while_asn_1381 = ActUnit_PushOutput_if_for_and_stg_2_7_sva & ActUnit_RunInst_switch_lp_equal_tmp_8
      & is_start_sva;
  assign while_asn_1383 = ~(is_start_sva & while_nor_itm);
  assign while_asn_1385 = ActUnit_RunInst_switch_lp_and_tmp & ActUnit_RunInst_switch_lp_equal_tmp_2
      & is_start_sva;
  assign while_asn_1387 = reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_nor_cse
      & ActUnit_RunInst_switch_lp_equal_tmp_4 & is_start_sva;
  assign while_asn_1389 = reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_nor_cse
      & ActUnit_RunInst_switch_lp_equal_tmp_5 & is_start_sva;
  assign while_asn_1391 = reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_nor_cse
      & ActUnit_RunInst_switch_lp_equal_tmp_6 & is_start_sva;
  assign while_asn_1393 = reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_nor_cse
      & ActUnit_RunInst_switch_lp_equal_tmp_7 & is_start_sva;
  assign while_asn_1395 = reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_nor_cse
      & ActUnit_RunInst_switch_lp_equal_tmp_8 & is_start_sva;
  assign nl_ActUnit_RunInst_case_2_for_i_4_0_sva_2 = conv_u2s_4_5(ActUnit_PushOutput_if_for_i_4_0_sva_3_0)
      + 5'b00001;
  assign ActUnit_RunInst_case_2_for_i_4_0_sva_2 = nl_ActUnit_RunInst_case_2_for_i_4_0_sva_2[4:0];
  assign nvhls_get_slc_2U_NVUINT8_return_3_sva_1 = MUX_v_2_32_2((act_config_inst_regs_0_sva_dfm_5[3:2]),
      (act_config_inst_regs_1_sva_dfm_5[3:2]), (act_config_inst_regs_2_sva_dfm_5[3:2]),
      (act_config_inst_regs_3_sva_dfm_5[3:2]), (act_config_inst_regs_4_sva_dfm_5[3:2]),
      (act_config_inst_regs_5_sva_dfm_5[3:2]), (act_config_inst_regs_6_sva_dfm_5[3:2]),
      (act_config_inst_regs_7_sva_dfm_5[3:2]), (act_config_inst_regs_8_sva_dfm_5[3:2]),
      (act_config_inst_regs_9_sva_dfm_5[3:2]), (act_config_inst_regs_10_sva_dfm_5[3:2]),
      (act_config_inst_regs_11_sva_dfm_5[3:2]), (act_config_inst_regs_12_sva_dfm_5[3:2]),
      (act_config_inst_regs_13_sva_dfm_5[3:2]), (act_config_inst_regs_14_sva_dfm_5[3:2]),
      (act_config_inst_regs_15_sva_dfm_5[3:2]), (act_config_inst_regs_16_sva_dfm_6[3:2]),
      (act_config_inst_regs_17_sva_dfm_6[3:2]), (act_config_inst_regs_18_sva_dfm_6[3:2]),
      (act_config_inst_regs_19_sva_dfm_6[3:2]), (act_config_inst_regs_20_sva_dfm_6[3:2]),
      (act_config_inst_regs_21_sva_dfm_6[3:2]), (act_config_inst_regs_22_sva_dfm_6[3:2]),
      (act_config_inst_regs_23_sva_dfm_6[3:2]), (act_config_inst_regs_24_sva_dfm_6[3:2]),
      (act_config_inst_regs_25_sva_dfm_6[3:2]), (act_config_inst_regs_26_sva_dfm_6[3:2]),
      (act_config_inst_regs_27_sva_dfm_6[3:2]), (act_config_inst_regs_28_sva_dfm_6[3:2]),
      (act_config_inst_regs_29_sva_dfm_6[3:2]), (act_config_inst_regs_30_sva_dfm_6[3:2]),
      (act_config_inst_regs_31_sva_dfm_6[3:2]), act_config_inst_counter_sva_dfm_3);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_65_0 = ~((nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b11));
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_67_0 = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1!=2'b00);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_69_0 = ~((nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b10));
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_71_0 = ~((nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b01));
  assign ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1
      = MUX_v_32_16_2(act_port_read_out_data_0_0_sva_dfm, act_port_read_out_data_0_1_sva_dfm,
      act_port_read_out_data_0_2_sva_dfm, act_port_read_out_data_0_3_sva_dfm, act_port_read_out_data_0_4_sva_dfm,
      act_port_read_out_data_0_5_sva_dfm, act_port_read_out_data_0_6_sva_dfm, act_port_read_out_data_0_7_sva_dfm,
      act_port_read_out_data_0_8_sva_dfm, act_port_read_out_data_0_9_sva_dfm, act_port_read_out_data_0_10_sva_dfm,
      act_port_read_out_data_0_11_sva_dfm, act_port_read_out_data_0_12_sva_dfm, act_port_read_out_data_0_13_sva_dfm,
      act_port_read_out_data_0_14_sva_dfm, act_port_read_out_data_0_15_sva_dfm, ActUnit_PushOutput_if_for_i_4_0_sva_3_0);
  assign act_config_InstIncr_if_act_config_InstIncr_if_if_nor_tmp = ~((act_config_output_counter_sva_dfm_3
      != (operator_8_false_acc_sdt_sva_1[7:0])) | (operator_8_false_acc_sdt_sva_1[8]));
  assign nl_operator_8_false_acc_sdt_sva_1 = conv_u2s_8_9(act_config_num_output_sva)
      + 9'b111111111;
  assign operator_8_false_acc_sdt_sva_1 = nl_operator_8_false_acc_sdt_sva_1[8:0];
  assign nl_operator_6_false_acc_tmp = conv_u2s_6_7(act_config_num_inst_sva) + 7'b1111111;
  assign operator_6_false_acc_tmp = nl_operator_6_false_acc_tmp[6:0];
  assign while_asn_1397 = ~(is_start_sva & w_load_lpi_1_dfm_1);
  assign while_asn_1399 = act_config_is_zero_first_sva_dfm_4 & w_load_lpi_1_dfm_1
      & is_start_sva;
  assign while_asn_1401 = (~ act_config_is_zero_first_sva_dfm_4) & w_load_lpi_1_dfm_1
      & is_start_sva;
  assign nl_Tanh_for_16_else_else_acc_nl = conv_s2s_26_31(nv_scvector_cctor_nv_scvector_6_for_16_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0])
      + conv_s2s_30_31(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_1_z[100:71]);
  assign Tanh_for_16_else_else_acc_nl = nl_Tanh_for_16_else_else_acc_nl[30:0];
  assign Tanh_for_Tanh_for_nor_15_nl = ~(Tanh_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | Tanh_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs);
  assign Tanh_for_and_79_nl = Tanh_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      & (~ Tanh_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs);
  assign Tanh_for_16_exs_5_30_0 = MUX1HOT_v_31_3_2(Tanh_for_16_else_else_acc_nl,
      31'b0000001000000000000000000000000, 31'b1111111000000000000000000000000, {Tanh_for_Tanh_for_nor_15_nl
      , Tanh_for_and_79_nl , Tanh_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs});
  assign nl_Tanh_for_15_else_else_acc_nl = conv_s2s_26_31(reg_nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6)
      + conv_s2s_30_31(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_2_z[100:71]);
  assign Tanh_for_15_else_else_acc_nl = nl_Tanh_for_15_else_else_acc_nl[30:0];
  assign Tanh_for_Tanh_for_nor_14_nl = ~(Tanh_for_15_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | Tanh_for_15_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs);
  assign Tanh_for_and_77_nl = Tanh_for_15_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      & (~ Tanh_for_15_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs);
  assign Tanh_for_15_exs_5_30_0 = MUX1HOT_v_31_3_2(Tanh_for_15_else_else_acc_nl,
      31'b0000001000000000000000000000000, 31'b1111111000000000000000000000000, {Tanh_for_Tanh_for_nor_14_nl
      , Tanh_for_and_77_nl , Tanh_for_15_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs});
  assign nl_Tanh_for_14_else_else_acc_nl = conv_s2s_26_31(reg_nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6)
      + conv_s2s_30_31(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_3_z[100:71]);
  assign Tanh_for_14_else_else_acc_nl = nl_Tanh_for_14_else_else_acc_nl[30:0];
  assign Tanh_for_Tanh_for_nor_13_nl = ~(Tanh_for_14_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | Tanh_for_14_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs);
  assign Tanh_for_and_75_nl = Tanh_for_14_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      & (~ Tanh_for_14_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs);
  assign Tanh_for_14_exs_5_30_0 = MUX1HOT_v_31_3_2(Tanh_for_14_else_else_acc_nl,
      31'b0000001000000000000000000000000, 31'b1111111000000000000000000000000, {Tanh_for_Tanh_for_nor_13_nl
      , Tanh_for_and_75_nl , Tanh_for_14_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs});
  assign nl_Tanh_for_13_else_else_acc_nl = conv_s2s_26_31(reg_nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6)
      + conv_s2s_30_31(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_4_z[100:71]);
  assign Tanh_for_13_else_else_acc_nl = nl_Tanh_for_13_else_else_acc_nl[30:0];
  assign Tanh_for_Tanh_for_nor_12_nl = ~(Tanh_for_13_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | Tanh_for_13_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs);
  assign Tanh_for_and_73_nl = Tanh_for_13_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      & (~ Tanh_for_13_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs);
  assign Tanh_for_13_exs_5_30_0 = MUX1HOT_v_31_3_2(Tanh_for_13_else_else_acc_nl,
      31'b0000001000000000000000000000000, 31'b1111111000000000000000000000000, {Tanh_for_Tanh_for_nor_12_nl
      , Tanh_for_and_73_nl , Tanh_for_13_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs});
  assign nl_Tanh_for_12_else_else_acc_nl = conv_s2s_26_31(reg_nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6)
      + conv_s2s_30_31(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_5_z[100:71]);
  assign Tanh_for_12_else_else_acc_nl = nl_Tanh_for_12_else_else_acc_nl[30:0];
  assign Tanh_for_Tanh_for_nor_11_nl = ~(Tanh_for_12_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | Tanh_for_12_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs);
  assign Tanh_for_and_71_nl = Tanh_for_12_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      & (~ Tanh_for_12_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs);
  assign Tanh_for_12_exs_5_30_0 = MUX1HOT_v_31_3_2(Tanh_for_12_else_else_acc_nl,
      31'b0000001000000000000000000000000, 31'b1111111000000000000000000000000, {Tanh_for_Tanh_for_nor_11_nl
      , Tanh_for_and_71_nl , Tanh_for_12_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs});
  assign nl_Tanh_for_11_else_else_acc_nl = conv_s2s_26_31(nv_scvector_cctor_nv_scvector_6_for_11_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0])
      + conv_s2s_30_31(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_6_z[100:71]);
  assign Tanh_for_11_else_else_acc_nl = nl_Tanh_for_11_else_else_acc_nl[30:0];
  assign Tanh_for_Tanh_for_nor_10_nl = ~(Tanh_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | Tanh_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs);
  assign Tanh_for_and_69_nl = Tanh_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      & (~ Tanh_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs);
  assign Tanh_for_11_exs_5_30_0 = MUX1HOT_v_31_3_2(Tanh_for_11_else_else_acc_nl,
      31'b0000001000000000000000000000000, 31'b1111111000000000000000000000000, {Tanh_for_Tanh_for_nor_10_nl
      , Tanh_for_and_69_nl , Tanh_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs});
  assign nl_Tanh_for_10_else_else_acc_nl = conv_s2s_26_31(nv_scvector_cctor_nv_scvector_6_for_10_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0])
      + conv_s2s_30_31(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_7_z[100:71]);
  assign Tanh_for_10_else_else_acc_nl = nl_Tanh_for_10_else_else_acc_nl[30:0];
  assign Tanh_for_Tanh_for_nor_9_nl = ~(Tanh_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | Tanh_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs);
  assign Tanh_for_and_67_nl = Tanh_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      & (~ Tanh_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs);
  assign Tanh_for_10_exs_5_30_0 = MUX1HOT_v_31_3_2(Tanh_for_10_else_else_acc_nl,
      31'b0000001000000000000000000000000, 31'b1111111000000000000000000000000, {Tanh_for_Tanh_for_nor_9_nl
      , Tanh_for_and_67_nl , Tanh_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs});
  assign nl_Tanh_for_9_else_else_acc_nl = conv_s2s_26_31(reg_nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6)
      + conv_s2s_30_31(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_8_z[100:71]);
  assign Tanh_for_9_else_else_acc_nl = nl_Tanh_for_9_else_else_acc_nl[30:0];
  assign Tanh_for_Tanh_for_nor_8_nl = ~(Tanh_for_9_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | Tanh_for_9_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs);
  assign Tanh_for_and_65_nl = Tanh_for_9_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      & (~ Tanh_for_9_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs);
  assign Tanh_for_9_exs_5_30_0 = MUX1HOT_v_31_3_2(Tanh_for_9_else_else_acc_nl, 31'b0000001000000000000000000000000,
      31'b1111111000000000000000000000000, {Tanh_for_Tanh_for_nor_8_nl , Tanh_for_and_65_nl
      , Tanh_for_9_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs});
  assign nl_Tanh_for_8_else_else_acc_nl = conv_s2s_26_31(reg_nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6)
      + conv_s2s_30_31(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_9_z[100:71]);
  assign Tanh_for_8_else_else_acc_nl = nl_Tanh_for_8_else_else_acc_nl[30:0];
  assign Tanh_for_Tanh_for_nor_7_nl = ~(Tanh_for_8_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | Tanh_for_8_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs);
  assign Tanh_for_and_63_nl = Tanh_for_8_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      & (~ Tanh_for_8_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs);
  assign Tanh_for_8_exs_5_30_0 = MUX1HOT_v_31_3_2(Tanh_for_8_else_else_acc_nl, 31'b0000001000000000000000000000000,
      31'b1111111000000000000000000000000, {Tanh_for_Tanh_for_nor_7_nl , Tanh_for_and_63_nl
      , Tanh_for_8_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs});
  assign nl_Tanh_for_7_else_else_acc_nl = conv_s2s_26_31(reg_nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6)
      + conv_s2s_30_31(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_10_z[100:71]);
  assign Tanh_for_7_else_else_acc_nl = nl_Tanh_for_7_else_else_acc_nl[30:0];
  assign Tanh_for_Tanh_for_nor_6_nl = ~(Tanh_for_7_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | Tanh_for_7_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs);
  assign Tanh_for_and_61_nl = Tanh_for_7_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      & (~ Tanh_for_7_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs);
  assign Tanh_for_7_exs_5_30_0 = MUX1HOT_v_31_3_2(Tanh_for_7_else_else_acc_nl, 31'b0000001000000000000000000000000,
      31'b1111111000000000000000000000000, {Tanh_for_Tanh_for_nor_6_nl , Tanh_for_and_61_nl
      , Tanh_for_7_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs});
  assign nl_Tanh_for_6_else_else_acc_nl = conv_s2s_26_31(reg_nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6)
      + conv_s2s_30_31(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_11_z[100:71]);
  assign Tanh_for_6_else_else_acc_nl = nl_Tanh_for_6_else_else_acc_nl[30:0];
  assign Tanh_for_Tanh_for_nor_5_nl = ~(Tanh_for_6_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | Tanh_for_6_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs);
  assign Tanh_for_and_59_nl = Tanh_for_6_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      & (~ Tanh_for_6_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs);
  assign Tanh_for_6_exs_5_30_0 = MUX1HOT_v_31_3_2(Tanh_for_6_else_else_acc_nl, 31'b0000001000000000000000000000000,
      31'b1111111000000000000000000000000, {Tanh_for_Tanh_for_nor_5_nl , Tanh_for_and_59_nl
      , Tanh_for_6_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs});
  assign nl_Tanh_for_5_else_else_acc_nl = conv_s2s_26_31(reg_nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6)
      + conv_s2s_30_31(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_12_z[100:71]);
  assign Tanh_for_5_else_else_acc_nl = nl_Tanh_for_5_else_else_acc_nl[30:0];
  assign Tanh_for_Tanh_for_nor_4_nl = ~(Tanh_for_5_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | Tanh_for_5_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs);
  assign Tanh_for_and_57_nl = Tanh_for_5_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      & (~ Tanh_for_5_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs);
  assign Tanh_for_5_exs_5_30_0 = MUX1HOT_v_31_3_2(Tanh_for_5_else_else_acc_nl, 31'b0000001000000000000000000000000,
      31'b1111111000000000000000000000000, {Tanh_for_Tanh_for_nor_4_nl , Tanh_for_and_57_nl
      , Tanh_for_5_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs});
  assign nl_Tanh_for_4_else_else_acc_nl = conv_s2s_26_31(reg_nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6)
      + conv_s2s_30_31(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_13_z[100:71]);
  assign Tanh_for_4_else_else_acc_nl = nl_Tanh_for_4_else_else_acc_nl[30:0];
  assign Tanh_for_Tanh_for_nor_3_nl = ~(Tanh_for_4_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | Tanh_for_4_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs);
  assign Tanh_for_and_55_nl = Tanh_for_4_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      & (~ Tanh_for_4_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs);
  assign Tanh_for_4_exs_5_30_0 = MUX1HOT_v_31_3_2(Tanh_for_4_else_else_acc_nl, 31'b0000001000000000000000000000000,
      31'b1111111000000000000000000000000, {Tanh_for_Tanh_for_nor_3_nl , Tanh_for_and_55_nl
      , Tanh_for_4_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs});
  assign nl_Tanh_for_3_else_else_acc_nl = conv_s2s_26_31(reg_nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6)
      + conv_s2s_30_31(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_14_z[100:71]);
  assign Tanh_for_3_else_else_acc_nl = nl_Tanh_for_3_else_else_acc_nl[30:0];
  assign Tanh_for_Tanh_for_nor_2_nl = ~(Tanh_for_3_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | Tanh_for_3_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs);
  assign Tanh_for_and_53_nl = Tanh_for_3_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      & (~ Tanh_for_3_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs);
  assign Tanh_for_3_exs_5_30_0 = MUX1HOT_v_31_3_2(Tanh_for_3_else_else_acc_nl, 31'b0000001000000000000000000000000,
      31'b1111111000000000000000000000000, {Tanh_for_Tanh_for_nor_2_nl , Tanh_for_and_53_nl
      , Tanh_for_3_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs});
  assign nl_Tanh_for_2_else_else_acc_nl = conv_s2s_26_31(reg_nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6)
      + conv_s2s_30_31(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_15_z[100:71]);
  assign Tanh_for_2_else_else_acc_nl = nl_Tanh_for_2_else_else_acc_nl[30:0];
  assign Tanh_for_Tanh_for_nor_1_nl = ~(Tanh_for_2_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | Tanh_for_2_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs);
  assign Tanh_for_and_51_nl = Tanh_for_2_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      & (~ Tanh_for_2_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs);
  assign Tanh_for_2_exs_5_30_0 = MUX1HOT_v_31_3_2(Tanh_for_2_else_else_acc_nl, 31'b0000001000000000000000000000000,
      31'b1111111000000000000000000000000, {Tanh_for_Tanh_for_nor_1_nl , Tanh_for_and_51_nl
      , Tanh_for_2_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs});
  assign nl_Tanh_for_1_else_else_acc_nl = conv_s2s_26_31(reg_ActUnit_RunInst_case_11_nv_scvector_cctor_data_0_ftd_6)
      + conv_s2s_30_31(Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_z[100:71]);
  assign Tanh_for_1_else_else_acc_nl = nl_Tanh_for_1_else_else_acc_nl[30:0];
  assign Tanh_for_Tanh_for_nor_nl = ~(Tanh_for_1_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | Tanh_for_1_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs);
  assign Tanh_for_and_49_nl = Tanh_for_1_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      & (~ Tanh_for_1_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs);
  assign Tanh_for_1_exs_5_30_0 = MUX1HOT_v_31_3_2(Tanh_for_1_else_else_acc_nl, 31'b0000001000000000000000000000000,
      31'b1111111000000000000000000000000, {Tanh_for_Tanh_for_nor_nl , Tanh_for_and_49_nl
      , Tanh_for_1_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs});
  assign ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_and_1_nl
      = MUX_v_5_2_2(5'b00000, act_write_addrs_lpi_1_dfm_5, ActUnit_RunInst_switch_lp_and_32_tmp);
  assign while_mux_55_tmp = MUX_v_5_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_2_mx0w2,
      ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_and_1_nl,
      is_start_sva);
  assign nor_57_cse = ~((fsm_output[1]) | (fsm_output[4]));
  assign and_dcpl_9 = is_start_sva & (act_config_in_InstFetch_mux_tmp[5]);
  assign and_dcpl_13 = and_dcpl_9 & (act_config_in_InstFetch_mux_tmp[4]);
  assign and_dcpl_47 = (act_config_in_InstFetch_mux_tmp[6]) & (~ (act_config_in_InstFetch_mux_tmp[4]));
  assign and_dcpl_51 = and_dcpl_9 & (act_config_in_InstFetch_mux_tmp[7]);
  assign and_dcpl_78 = and_dcpl_51 & and_dcpl_47;
  assign and_dcpl_162 = is_start_sva & (act_config_in_InstFetch_return_sva_7_2[5:3]==3'b111);
  assign and_dcpl_366 = (fsm_output[1]) & (~ (fsm_output[4]));
  assign and_dcpl_368 = nor_734_cse & (fsm_output[0]) & and_dcpl_366;
  assign nor_61_cse = ~((~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[8]))
      | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11:9]!=3'b100));
  assign nor_60_nl = ~(is_start_sva | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt) |
      (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[8])) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11:9]!=3'b100));
  assign or_170_nl = is_start_sva | nor_61_cse;
  assign mux_51_cse = MUX_s_1_2_2(nor_60_nl, or_170_nl, ActUnit_RunInst_switch_lp_and_32_tmp);
  assign and_dcpl_369 = mux_51_cse & and_dcpl_368;
  assign and_dcpl_370 = is_start_sva & w_load_lpi_1_dfm_1;
  assign or_tmp_68 = is_start_sva | rva_in_PopNB_mioi_data_rw_rsc_z_mxwt | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[8]))
      | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11:9]!=3'b100);
  assign nor_63_nl = ~(rva_in_PopNB_mioi_data_rw_rsc_z_mxwt | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[8]))
      | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11:9]!=3'b100));
  assign mux_54_nl = MUX_s_1_2_2(nor_63_nl, ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_2_tmp,
      is_start_sva);
  assign mux_tmp_55 = MUX_s_1_2_2((~ mux_54_nl), or_tmp_68, ActUnit_RunInst_switch_lp_and_32_tmp);
  assign and_dcpl_374 = (~ mux_tmp_55) & and_dcpl_368;
  assign and_dcpl_377 = is_start_sva & ActUnit_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva;
  assign nand_nl = ~(act_config_is_zero_first_sva_dfm_4 & w_load_lpi_1_dfm_1);
  assign or_86_nl = act_config_is_zero_first_sva_dfm_4 | (~ w_load_lpi_1_dfm_1);
  assign mux_48_nl = MUX_s_1_2_2(nand_nl, or_86_nl, act_config_is_zero_first_sva);
  assign and_dcpl_379 = (reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_1_cse
      | reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_cse | reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_nor_cse
      | reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_2_cse) &
      (ActUnit_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva
      | mux_48_nl) & is_start_sva & ActUnit_RunInst_switch_lp_equal_tmp_7;
  assign or_tmp_111 = (~ act_config_is_valid_sva) | is_start_sva;
  assign and_dcpl_553 = nor_734_cse & (fsm_output[0]);
  assign and_dcpl_554 = and_dcpl_553 & nor_57_cse;
  assign and_dcpl_556 = nor_734_cse & (~ (fsm_output[0]));
  assign and_dcpl_557 = and_dcpl_556 & and_dcpl_366;
  assign and_dcpl_559 = (fsm_output[0]) & (fsm_output[1]) & (~ (fsm_output[4]));
  assign and_dcpl_560 = ~((act_config_in_InstFetch_return_sva_7_2[2]) | (fsm_output[3]));
  assign and_dcpl_562 = and_dcpl_560 & (~ (fsm_output[2])) & and_dcpl_559;
  assign or_tmp_126 = (fsm_output[3]) | (act_config_in_InstFetch_return_sva_7_2[2]);
  assign and_dcpl_563 = ~((fsm_output[1:0]!=2'b00));
  assign and_dcpl_564 = and_dcpl_563 & (~ (fsm_output[4]));
  assign and_dcpl_565 = and_dcpl_560 & (fsm_output[2]);
  assign and_dcpl_566 = and_dcpl_565 & and_dcpl_564;
  assign and_dcpl_568 = (fsm_output[0]) & (~ (fsm_output[1])) & (~ (fsm_output[4]));
  assign and_dcpl_569 = and_dcpl_565 & and_dcpl_568;
  assign and_dcpl_570 = (fsm_output[1:0]==2'b10);
  assign and_dcpl_571 = and_dcpl_570 & (~ (fsm_output[4]));
  assign and_dcpl_572 = and_dcpl_565 & and_dcpl_571;
  assign and_dcpl_573 = and_dcpl_565 & and_dcpl_559;
  assign and_dcpl_574 = (fsm_output[3:2]==2'b10);
  assign and_dcpl_575 = and_dcpl_574 & (~ (fsm_output[0]));
  assign and_dcpl_576 = and_dcpl_575 & nor_57_cse;
  assign and_dcpl_577 = and_dcpl_574 & (fsm_output[0]);
  assign and_dcpl_578 = and_dcpl_577 & nor_57_cse;
  assign and_dcpl_579 = (act_config_in_InstFetch_return_sva_7_2[2]) & (~ (fsm_output[3]));
  assign and_dcpl_581 = and_dcpl_579 & (~ (fsm_output[2])) & and_dcpl_559;
  assign and_dcpl_582 = and_dcpl_579 & (fsm_output[2]);
  assign and_dcpl_583 = and_dcpl_582 & and_dcpl_564;
  assign and_dcpl_584 = and_dcpl_582 & and_dcpl_568;
  assign and_dcpl_585 = and_dcpl_582 & and_dcpl_571;
  assign and_dcpl_586 = and_dcpl_582 & and_dcpl_559;
  assign and_dcpl_587 = is_start_sva & (~ (fsm_output[4]));
  assign or_tmp_131 = Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
      | Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign or_tmp_133 = Tanh_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
      | Tanh_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  assign or_tmp_134 = Gelu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
      | Gelu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs;
  assign or_tmp_135 = Gelu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
      | Gelu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs;
  assign or_tmp_136 = Gelu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
      | Gelu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs;
  assign and_tmp_9 = or_tmp_136 & or_tmp_135;
  assign or_tmp_139 = Gelu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
      | Gelu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs;
  assign or_tmp_140 = Gelu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
      | Gelu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs;
  assign and_tmp_11 = or_tmp_140 & or_tmp_139;
  assign nand_180_cse = ~((act_config_in_InstFetch_mux_tmp[7:5]==3'b111));
  assign nand_181_cse = ~((act_config_in_InstFetch_mux_tmp[7]) & (act_config_in_InstFetch_mux_tmp[5]));
  assign nor_128_nl = ~(operator_32_8_true_AC_TRN_AC_WRAP_1_less_14_tmp | operator_32_8_true_AC_TRN_AC_WRAP_2_less_14_tmp
      | nand_180_cse);
  assign nor_129_nl = ~(operator_32_8_true_AC_TRN_AC_WRAP_2_less_14_tmp_1 | operator_32_8_true_AC_TRN_AC_WRAP_3_less_14_tmp
      | nand_181_cse);
  assign not_tmp_248 = MUX_s_1_2_2(nor_128_nl, nor_129_nl, act_config_in_InstFetch_mux_tmp[4]);
  assign nand_tmp_3 = ~((fsm_output[0]) & not_tmp_248);
  assign or_tmp_146 = Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
      | Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign or_tmp_147 = Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
      | Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign or_tmp_148 = Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
      | Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign or_tmp_151 = Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
      | Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign or_tmp_159 = Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
      | Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign or_tmp_161 = Tanh_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
      | Tanh_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  assign or_tmp_162 = Gelu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
      | Gelu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs;
  assign or_tmp_163 = Gelu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
      | Gelu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs;
  assign or_tmp_164 = Gelu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
      | Gelu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs;
  assign or_tmp_167 = Gelu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
      | Gelu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs;
  assign or_tmp_168 = Gelu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
      | Gelu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs;
  assign nor_130_nl = ~(operator_32_8_true_AC_TRN_AC_WRAP_1_less_15_tmp | operator_32_8_true_AC_TRN_AC_WRAP_2_less_15_tmp
      | nand_180_cse);
  assign nor_131_nl = ~(operator_32_8_true_AC_TRN_AC_WRAP_2_less_15_tmp_1 | operator_32_8_true_AC_TRN_AC_WRAP_3_less_15_tmp
      | nand_181_cse);
  assign not_tmp_255 = MUX_s_1_2_2(nor_130_nl, nor_131_nl, act_config_in_InstFetch_mux_tmp[4]);
  assign nand_tmp_9 = ~((fsm_output[0]) & not_tmp_255);
  assign or_tmp_174 = Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
      | Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign or_tmp_175 = Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
      | Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign or_tmp_176 = Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
      | Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign or_tmp_179 = Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
      | Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign and_dcpl_590 = (fsm_output[3:2]==2'b01);
  assign and_dcpl_591 = and_dcpl_590 & (~ (fsm_output[0]));
  assign and_dcpl_592 = and_dcpl_591 & nor_57_cse;
  assign or_tmp_184 = (fsm_output[2]) | (~ (fsm_output[0])) | operator_32_8_true_AC_TRN_AC_WRAP_2_less_3_tmp_1
      | operator_32_8_true_AC_TRN_AC_WRAP_3_less_3_tmp | (act_config_in_InstFetch_mux_tmp[7:4]!=4'b1111)
      | (fsm_output[1]) | (fsm_output[3]);
  assign and_dcpl_596 = is_start_sva & (act_config_in_InstFetch_return_sva_7_2[5])
      & (act_config_in_InstFetch_return_sva_7_2[3]);
  assign and_dcpl_599 = and_dcpl_590 & (fsm_output[0]);
  assign and_dcpl_600 = and_dcpl_599 & and_dcpl_366;
  assign not_tmp_262 = ~((act_config_in_InstFetch_mux_tmp[7:4]==4'b1111));
  assign or_tmp_198 = (fsm_output[1:0]!=2'b01) | operator_32_8_true_AC_TRN_AC_WRAP_2_less_tmp_1
      | operator_32_8_true_AC_TRN_AC_WRAP_3_less_tmp | not_tmp_262;
  assign and_dcpl_604 = (~((act_config_in_InstFetch_return_sva_7_2[4]) | (fsm_output[3])))
      & (fsm_output[2]) & and_dcpl_564;
  assign or_tmp_211 = (fsm_output[3:2]!=2'b01);
  assign or_tmp_213 = (~ (fsm_output[0])) | (fsm_output[2]) | (~ (fsm_output[3]));
  assign mux_152_nl = MUX_s_1_2_2(or_tmp_213, or_tmp_211, fsm_output[1]);
  assign and_dcpl_609 = ~(mux_152_nl | (fsm_output[4]));
  assign and_dcpl_612 = (act_config_in_InstFetch_return_sva_7_2[4]) & (fsm_output[3:2]==2'b01)
      & and_dcpl_564;
  assign and_dcpl_613 = and_dcpl_599 & nor_57_cse;
  assign and_dcpl_614 = and_dcpl_591 & and_dcpl_366;
  assign or_tmp_215 = (fsm_output[1:0]!=2'b00) | Tanh_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
      | Tanh_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  assign and_tmp_39 = ((~ (fsm_output[0])) | Gelu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
      | Gelu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & or_tmp_164 & and_tmp_11;
  assign or_tmp_229 = (fsm_output[1:0]!=2'b01) | operator_32_8_true_AC_TRN_AC_WRAP_2_less_1_tmp_1
      | operator_32_8_true_AC_TRN_AC_WRAP_3_less_1_tmp | not_tmp_262;
  assign and_dcpl_616 = (fsm_output[2]) & (~ (fsm_output[4]));
  assign and_dcpl_620 = (~ (act_config_in_InstFetch_return_sva_7_2[4])) & (act_config_in_InstFetch_return_sva_7_2[2]);
  assign and_dcpl_621 = and_dcpl_596 & and_dcpl_620;
  assign or_tmp_237 = (fsm_output[1]) | Tanh_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
      | Tanh_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
      | (fsm_output[0]);
  assign and_710_nl = or_tmp_136 & or_tmp_168;
  assign and_709_nl = or_tmp_136 & or_tmp_135 & or_tmp_168;
  assign mux_tmp_169 = MUX_s_1_2_2(and_710_nl, and_709_nl, fsm_output[0]);
  assign or_tmp_249 = (fsm_output[1:0]!=2'b01) | operator_32_8_true_AC_TRN_AC_WRAP_2_less_2_tmp_1
      | operator_32_8_true_AC_TRN_AC_WRAP_3_less_2_tmp | not_tmp_262;
  assign or_dcpl_290 = and_dcpl_563 | (~ (fsm_output[2]));
  assign and_dcpl_668 = and_dcpl_596 & or_dcpl_290;
  assign and_dcpl_746 = is_start_sva & (~ (fsm_output[3]));
  assign and_dcpl_747 = and_dcpl_746 & (~ (fsm_output[2]));
  assign and_dcpl_748 = and_dcpl_747 & (fsm_output[0]) & (~ (fsm_output[4]));
  assign not_tmp_311 = ~((act_config_in_InstFetch_return_sva_7_2[3]) & (act_config_in_InstFetch_return_sva_7_2[5]));
  assign and_dcpl_767 = and_dcpl_570 & (fsm_output[4]);
  assign and_dcpl_768 = and_dcpl_747 & and_dcpl_767;
  assign and_dcpl_770 = (fsm_output[3:2]==2'b11);
  assign and_dcpl_774 = ~(is_start_sva | (fsm_output[3]));
  assign and_dcpl_775 = and_dcpl_774 & (fsm_output[2]);
  assign and_dcpl_786 = and_dcpl_774 & (~ (fsm_output[2]));
  assign and_dcpl_788 = and_dcpl_553 & and_dcpl_366;
  assign and_dcpl_789 = (fsm_output[1]) & (fsm_output[4]);
  assign and_dcpl_794 = and_dcpl_786 & and_dcpl_767;
  assign or_dcpl_296 = (~((fsm_output[1:0]==2'b11))) | (fsm_output[4]);
  assign or_dcpl_297 = is_start_sva | (fsm_output[3]);
  assign or_dcpl_299 = or_dcpl_297 | (fsm_output[2]) | or_dcpl_296;
  assign or_dcpl_300 = (~ rva_in_PopNB_mioi_return_rsc_z_mxwt) | rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  assign and_dcpl_797 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11:8]==4'b1000);
  assign or_dcpl_301 = and_dcpl_797 | or_dcpl_300;
  assign or_dcpl_303 = ~(rva_in_PopNB_mioi_return_rsc_z_mxwt & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt);
  assign or_dcpl_304 = and_dcpl_797 | or_dcpl_303;
  assign and_dcpl_798 = (~ (fsm_output[1])) & (fsm_output[4]);
  assign and_dcpl_799 = nor_734_cse & and_dcpl_798;
  assign or_dcpl_310 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[8]) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | is_start_sva | or_1033_cse;
  assign or_dcpl_320 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[10]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[9]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt);
  assign or_dcpl_322 = (~ (fsm_output[1])) | (fsm_output[4]);
  assign and_dcpl_802 = nor_734_cse & and_dcpl_570;
  assign and_dcpl_803 = and_dcpl_802 & (fsm_output[4]) & w_axi_rsp_lpi_1_dfm_1 &
      act_read_req_valid_lpi_1_dfm_6;
  assign and_dcpl_805 = and_dcpl_802 & (~(act_read_req_valid_lpi_1_dfm_6 & w_axi_rsp_lpi_1_dfm_1))
      & (fsm_output[4]);
  assign or_dcpl_328 = (while_mux_55_tmp[4]) | (while_mux_55_tmp[1]);
  assign or_dcpl_329 = (while_mux_55_tmp[3:2]!=2'b00);
  assign or_dcpl_330 = or_dcpl_329 | or_dcpl_328;
  assign or_dcpl_332 = or_1077_cse | (~ (fsm_output[1]));
  assign or_dcpl_333 = or_dcpl_332 | (fsm_output[4]) | (while_mux_55_tmp[0]);
  assign or_dcpl_335 = (~ mux_51_cse) | (fsm_output[3]);
  assign or_dcpl_338 = or_dcpl_332 | (fsm_output[4]) | (~ (while_mux_55_tmp[0]));
  assign or_dcpl_341 = (while_mux_55_tmp[4]) | (~ (while_mux_55_tmp[1]));
  assign or_dcpl_342 = or_dcpl_329 | or_dcpl_341;
  assign or_dcpl_347 = (while_mux_55_tmp[3:2]!=2'b01);
  assign or_dcpl_348 = or_dcpl_347 | or_dcpl_328;
  assign or_dcpl_353 = or_dcpl_347 | or_dcpl_341;
  assign or_dcpl_358 = (while_mux_55_tmp[3:2]!=2'b10);
  assign or_dcpl_359 = or_dcpl_358 | or_dcpl_328;
  assign or_dcpl_364 = or_dcpl_358 | or_dcpl_341;
  assign or_dcpl_369 = ~((while_mux_55_tmp[3:2]==2'b11));
  assign or_dcpl_370 = or_dcpl_369 | or_dcpl_328;
  assign or_dcpl_375 = or_dcpl_369 | or_dcpl_341;
  assign or_dcpl_380 = (~ (while_mux_55_tmp[4])) | (while_mux_55_tmp[1]);
  assign or_dcpl_381 = or_dcpl_329 | or_dcpl_380;
  assign or_dcpl_386 = ~((while_mux_55_tmp[4]) & (while_mux_55_tmp[1]));
  assign or_dcpl_387 = or_dcpl_329 | or_dcpl_386;
  assign or_dcpl_392 = or_dcpl_347 | or_dcpl_380;
  assign or_dcpl_397 = or_dcpl_347 | or_dcpl_386;
  assign or_dcpl_402 = or_dcpl_358 | or_dcpl_380;
  assign or_dcpl_407 = or_dcpl_358 | or_dcpl_386;
  assign or_dcpl_412 = or_dcpl_369 | or_dcpl_380;
  assign or_dcpl_417 = or_dcpl_369 | or_dcpl_386;
  assign not_tmp_347 = ~((ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_23_4_mx1_tmp_7_0==8'b00000011)
      & act_config_ActConfigRead_else_unequal_tmp_1 & act_config_ActConfigRead_unequal_tmp_1
      & (~ ActUnit_DecodeAxiRead_unequal_tmp_1) & ActUnit_DecodeAxi_rva_in_reg_rw_sva_mx1
      & ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_mx1
      & (~ is_start_sva));
  assign or_dcpl_423 = or_1033_cse | (~ (fsm_output[0]));
  assign and_dcpl_814 = and_dcpl_556 & and_dcpl_789;
  assign and_dcpl_829 = and_dcpl_786 & and_dcpl_559;
  assign or_tmp_315 = (fsm_output[3:0]!=4'b0011);
  assign mux_tmp_196 = MUX_s_1_2_2((~ (fsm_output[3])), (fsm_output[3]), fsm_output[2]);
  assign mux_tmp_197 = MUX_s_1_2_2(and_dcpl_770, mux_tmp_196, fsm_output[0]);
  assign nor_tmp_46 = (fsm_output[0]) & (fsm_output[2]) & (fsm_output[3]);
  assign and_dcpl_831 = and_dcpl_770 & (~ (fsm_output[0]));
  assign and_dcpl_832 = and_dcpl_831 & and_dcpl_366;
  assign nor_139_cse = ~((fsm_output[1:0]!=2'b10));
  assign or_tmp_317 = nor_139_cse | (fsm_output[3:2]!=2'b00);
  assign or_dcpl_440 = (~((fsm_output[0]) ^ (fsm_output[1]))) | (fsm_output[4:2]!=3'b000);
  assign or_dcpl_442 = or_dcpl_423 | (fsm_output[1]) | (fsm_output[4]);
  assign mux_tmp_203 = MUX_s_1_2_2(nor_734_cse, mux_tmp_196, fsm_output[0]);
  assign and_dcpl_834 = ~((fsm_output[4:3]!=2'b00));
  assign or_tmp_318 = (fsm_output[0]) | (~ (fsm_output[2]));
  assign mux_205_itm = MUX_s_1_2_2(or_tmp_318, (fsm_output[2]), fsm_output[1]);
  assign nand_195_cse = ~((fsm_output[0]) & (fsm_output[2]));
  assign or_dcpl_443 = (fsm_output[2:1]!=2'b00);
  assign and_dcpl_849 = and_dcpl_553 & and_dcpl_798;
  assign or_tmp_322 = (fsm_output[3:0]!=4'b0000);
  assign mux_tmp_214 = MUX_s_1_2_2(nor_734_cse, mux_tmp_196, and_1104_cse);
  assign mux_215_itm = MUX_s_1_2_2(mux_tmp_214, or_tmp_322, fsm_output[4]);
  assign and_dcpl_852 = nor_tmp_46 & and_dcpl_366;
  assign or_dcpl_447 = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3:2]!=2'b00);
  assign or_dcpl_448 = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1:0]!=2'b00);
  assign or_dcpl_449 = or_dcpl_448 | or_dcpl_447;
  assign and_dcpl_853 = ~((ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]));
  assign and_dcpl_854 = and_dcpl_853 & (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]));
  assign and_dcpl_855 = ~((nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b00));
  assign and_dcpl_856 = ~(act_config_is_zero_first_sva_dfm_4 | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]));
  assign and_dcpl_857 = and_dcpl_856 & and_dcpl_855;
  assign or_dcpl_450 = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign or_dcpl_451 = or_dcpl_450 | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign or_dcpl_452 = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]) | (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]);
  assign or_dcpl_453 = or_dcpl_452 | (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]);
  assign or_dcpl_455 = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1:0]!=2'b01);
  assign or_dcpl_456 = or_dcpl_455 | or_dcpl_447;
  assign and_dcpl_860 = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]) & (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]));
  assign and_dcpl_861 = and_dcpl_860 & (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]));
  assign or_dcpl_457 = (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign or_dcpl_458 = or_dcpl_457 | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign or_dcpl_460 = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3:2]!=2'b10);
  assign or_dcpl_461 = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1:0]!=2'b10);
  assign or_dcpl_462 = or_dcpl_461 | or_dcpl_460;
  assign and_dcpl_864 = (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])) & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign and_dcpl_865 = and_dcpl_864 & (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]));
  assign and_dcpl_866 = (~ act_config_is_zero_first_sva_dfm_4) & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]);
  assign and_dcpl_867 = and_dcpl_866 & and_dcpl_855;
  assign or_dcpl_463 = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]));
  assign or_dcpl_464 = or_dcpl_463 | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign or_dcpl_465 = (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])) | (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]);
  assign or_dcpl_466 = or_dcpl_465 | (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]);
  assign or_dcpl_468 = ~((ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1:0]==2'b11));
  assign or_dcpl_469 = or_dcpl_468 | or_dcpl_460;
  assign and_dcpl_870 = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]) & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign and_dcpl_871 = and_dcpl_870 & (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]));
  assign or_dcpl_470 = ~((ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]) & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]));
  assign or_dcpl_471 = or_dcpl_470 | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign or_dcpl_473 = ~((ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3:2]==2'b11));
  assign or_dcpl_474 = or_dcpl_448 | or_dcpl_473;
  assign and_dcpl_874 = and_dcpl_864 & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign or_dcpl_475 = or_dcpl_463 | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]));
  assign or_dcpl_477 = or_dcpl_455 | or_dcpl_473;
  assign and_dcpl_877 = and_dcpl_870 & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign or_dcpl_478 = or_dcpl_470 | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]));
  assign or_dcpl_480 = or_dcpl_461 | or_dcpl_473;
  assign or_dcpl_482 = or_dcpl_461 | or_dcpl_447;
  assign or_dcpl_484 = or_dcpl_468 | or_dcpl_447;
  assign or_dcpl_486 = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3:2]!=2'b01);
  assign or_dcpl_487 = or_dcpl_448 | or_dcpl_486;
  assign or_dcpl_489 = or_dcpl_455 | or_dcpl_486;
  assign and_dcpl_888 = and_dcpl_853 & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign or_dcpl_490 = or_dcpl_450 | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]));
  assign or_dcpl_492 = or_dcpl_461 | or_dcpl_486;
  assign and_dcpl_891 = and_dcpl_860 & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign or_dcpl_493 = or_dcpl_457 | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]));
  assign or_dcpl_495 = or_dcpl_468 | or_dcpl_486;
  assign or_dcpl_497 = or_dcpl_448 | or_dcpl_460;
  assign or_dcpl_499 = or_dcpl_455 | or_dcpl_460;
  assign and_dcpl_900 = and_dcpl_577 & and_dcpl_366;
  assign or_tmp_323 = (fsm_output[0]) | (~ and_dcpl_770);
  assign mux_216_nl = MUX_s_1_2_2(or_tmp_323, or_1033_cse, fsm_output[4]);
  assign and_dcpl_901 = ~(mux_216_nl | (fsm_output[1]));
  assign and_dcpl_903 = (~ (fsm_output[2])) & (fsm_output[0]) & and_dcpl_366;
  assign and_dcpl_906 = rva_in_PopNB_mioi_return_rsc_z_mxwt & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & and_dcpl_774 & and_dcpl_903;
  assign and_dcpl_908 = (~((~(or_dcpl_303 | is_start_sva)) | (fsm_output[3]))) &
      and_dcpl_903;
  assign and_dcpl_909 = and_dcpl_747 & and_dcpl_559;
  assign and_dcpl_916 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7:0]==8'b00000010);
  assign or_dcpl_503 = ~((ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]) & (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]));
  assign or_dcpl_504 = or_dcpl_503 | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]));
  assign or_dcpl_507 = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]) | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]));
  assign or_dcpl_508 = or_dcpl_507 | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]));
  assign and_dcpl_923 = (nvhls_get_slc_2U_NVUINT8_return_3_sva==2'b10);
  assign and_dcpl_924 = and_dcpl_866 & and_dcpl_923;
  assign or_dcpl_523 = or_dcpl_465 | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]));
  assign and_dcpl_929 = and_dcpl_856 & and_dcpl_923;
  assign or_dcpl_526 = or_dcpl_452 | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]));
  assign and_dcpl_958 = (nvhls_get_slc_2U_NVUINT8_return_3_sva==2'b01);
  assign and_dcpl_959 = and_dcpl_866 & and_dcpl_958;
  assign or_dcpl_541 = or_dcpl_503 | (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]);
  assign and_dcpl_964 = and_dcpl_856 & and_dcpl_958;
  assign or_dcpl_544 = or_dcpl_507 | (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]);
  assign and_dcpl_997 = nor_tmp_46 & nor_57_cse;
  assign or_tmp_330 = ~(nand_195_cse & (fsm_output[3]));
  assign or_tmp_331 = (fsm_output[3:2]!=2'b10);
  assign and_dcpl_1001 = (fsm_output[4:3]==2'b01);
  assign mux_228_nl = MUX_s_1_2_2((~ and_dcpl_770), or_tmp_331, or_992_cse);
  assign mux_229_itm = MUX_s_1_2_2(mux_228_nl, or_1097_cse, fsm_output[4]);
  assign mux_230_nl = MUX_s_1_2_2(or_tmp_323, or_tmp_331, fsm_output[1]);
  assign mux_231_itm = MUX_s_1_2_2(mux_230_nl, or_1097_cse, fsm_output[4]);
  assign and_dcpl_1006 = and_dcpl_575 & and_dcpl_366;
  assign mux_233_nl = MUX_s_1_2_2(or_tmp_323, or_tmp_213, fsm_output[1]);
  assign mux_234_itm = MUX_s_1_2_2(mux_233_nl, or_1097_cse, fsm_output[4]);
  assign and_dcpl_1007 = and_dcpl_831 & nor_57_cse;
  assign mux_235_itm = MUX_s_1_2_2(nand_297_cse, or_tmp_322, fsm_output[4]);
  assign or_dcpl_561 = (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b00);
  assign or_dcpl_563 = or_1488_cse | or_dcpl_561;
  assign or_dcpl_566 = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]));
  assign or_dcpl_567 = or_dcpl_566 | or_dcpl_561;
  assign or_dcpl_582 = (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b01);
  assign or_dcpl_583 = or_1488_cse | or_dcpl_582;
  assign or_dcpl_586 = or_dcpl_566 | or_dcpl_582;
  assign or_dcpl_601 = (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b10);
  assign or_dcpl_602 = or_1488_cse | or_dcpl_601;
  assign or_dcpl_605 = or_dcpl_566 | or_dcpl_601;
  assign or_dcpl_620 = ~((nvhls_get_slc_2U_NVUINT8_return_3_sva==2'b11));
  assign or_dcpl_621 = or_1488_cse | or_dcpl_620;
  assign or_dcpl_624 = or_dcpl_566 | or_dcpl_620;
  assign act_config_output_counter_sva_mx0c1 = and_dcpl_553 & and_dcpl_789 & (~ ActUnit_CheckStart_start_reg_sva);
  assign act_config_inst_counter_sva_mx0c1 = and_dcpl_814 & (~(is_start_sva & is_incr_lpi_1_dfm_1));
  assign ActUnit_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva_mx0c2
      = and_dcpl_775 & and_dcpl_568;
  assign ActUnit_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva_mx0c3
      = and_dcpl_556 & and_dcpl_798;
  assign nand_214_nl = ~((fsm_output[0]) & mux_tmp_196);
  assign or_605_nl = or_1033_cse | (fsm_output[0]);
  assign mux_212_nl = MUX_s_1_2_2(nand_214_nl, or_605_nl, fsm_output[4]);
  assign ActUnit_PushOutput_if_for_i_4_0_sva_3_0_mx0c0 = ~(mux_212_nl | (fsm_output[1]));
  assign act_regs_data_0_0_sva_8_mx3c1 = ~((~(or_dcpl_453 | or_dcpl_451)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_0_1_sva_8_mx3c1 = ~((~(or_dcpl_453 | or_dcpl_458)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_0_10_sva_8_mx3c1 = ~((~(or_dcpl_466 | or_dcpl_464)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_0_11_sva_8_mx3c1 = ~((~(or_dcpl_466 | or_dcpl_471)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_0_12_sva_8_mx3c1 = ~((~(or_dcpl_453 | or_dcpl_475)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_0_13_sva_8_mx3c1 = ~((~(or_dcpl_453 | or_dcpl_478)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_0_14_sva_8_mx3c1 = ~((~(or_dcpl_466 | or_dcpl_475)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_0_15_sva_8_mx3c1 = ~((~(or_dcpl_466 | or_dcpl_478)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_0_2_sva_8_mx3c1 = ~((~(or_dcpl_466 | or_dcpl_451)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_0_3_sva_8_mx3c1 = ~((~(or_dcpl_466 | or_dcpl_458)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_0_4_sva_8_mx3c1 = ~((~(or_dcpl_453 | or_dcpl_490)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_0_5_sva_8_mx3c1 = ~((~(or_dcpl_453 | or_dcpl_493)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_0_6_sva_8_mx3c1 = ~((~(or_dcpl_466 | or_dcpl_490)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_0_7_sva_8_mx3c1 = ~((~(or_dcpl_466 | or_dcpl_493)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_0_8_sva_8_mx3c1 = ~((~(or_dcpl_453 | or_dcpl_464)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_3_0_sva_8_mx2c1 = ~((~(or_dcpl_508 | or_dcpl_451)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_2_15_sva_8_mx2c1 = ~((~(or_dcpl_523 | or_dcpl_478)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_2_14_sva_8_mx2c1 = ~((~(or_dcpl_523 | or_dcpl_475)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_2_13_sva_8_mx2c1 = ~((~(or_dcpl_526 | or_dcpl_478)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_2_12_sva_8_mx2c1 = ~((~(or_dcpl_526 | or_dcpl_475)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_2_11_sva_8_mx2c1 = ~((~(or_dcpl_523 | or_dcpl_471)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_2_10_sva_8_mx2c1 = ~((~(or_dcpl_523 | or_dcpl_464)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_2_9_sva_8_mx2c1 = ~((~(or_dcpl_526 | or_dcpl_471)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_2_8_sva_8_mx2c1 = ~((~(or_dcpl_526 | or_dcpl_464)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_2_7_sva_8_mx2c1 = ~((~(or_dcpl_523 | or_dcpl_493)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_2_6_sva_8_mx2c1 = ~((~(or_dcpl_523 | or_dcpl_490)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_2_5_sva_8_mx2c1 = ~((~(or_dcpl_526 | or_dcpl_493)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_2_4_sva_8_mx2c1 = ~((~(or_dcpl_526 | or_dcpl_490)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_2_3_sva_8_mx2c1 = ~((~(or_dcpl_523 | or_dcpl_458)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_2_2_sva_8_mx2c1 = ~((~(or_dcpl_523 | or_dcpl_451)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_2_1_sva_8_mx2c1 = ~((~(or_dcpl_526 | or_dcpl_458)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_2_0_sva_8_mx2c1 = ~((~(or_dcpl_526 | or_dcpl_451)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_1_15_sva_8_mx2c1 = ~((~(or_dcpl_541 | or_dcpl_478)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_1_14_sva_8_mx2c1 = ~((~(or_dcpl_541 | or_dcpl_475)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_1_13_sva_8_mx2c1 = ~((~(or_dcpl_544 | or_dcpl_478)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_1_12_sva_8_mx2c1 = ~((~(or_dcpl_544 | or_dcpl_475)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_1_11_sva_8_mx2c1 = ~((~(or_dcpl_541 | or_dcpl_471)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_1_10_sva_8_mx2c1 = ~((~(or_dcpl_541 | or_dcpl_464)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_1_9_sva_8_mx2c1 = ~((~(or_dcpl_544 | or_dcpl_471)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_1_8_sva_8_mx2c1 = ~((~(or_dcpl_544 | or_dcpl_464)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_1_7_sva_8_mx2c1 = ~((~(or_dcpl_541 | or_dcpl_493)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_1_6_sva_8_mx2c1 = ~((~(or_dcpl_541 | or_dcpl_490)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_1_5_sva_8_mx2c1 = ~((~(or_dcpl_544 | or_dcpl_493)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_1_4_sva_8_mx2c1 = ~((~(or_dcpl_544 | or_dcpl_490)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_1_3_sva_8_mx2c1 = ~((~(or_dcpl_541 | or_dcpl_458)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_1_2_sva_8_mx2c1 = ~((~(or_dcpl_541 | or_dcpl_451)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_1_1_sva_8_mx2c1 = ~((~(or_dcpl_544 | or_dcpl_458)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_1_0_sva_8_mx2c1 = ~((~(or_dcpl_544 | or_dcpl_451)) | act_config_is_zero_first_sva_dfm_4);
  assign act_regs_data_0_9_sva_8_mx2c1 = ~((~(or_dcpl_453 | or_dcpl_471)) | act_config_is_zero_first_sva_dfm_4);
  assign ActUnit_RunInst_switch_lp_and_817_enex5 = ActUnit_RunInst_switch_lp_and_802_cse
      & (reg_act_config_inst_regs_1_sva_dfm_5_enexo_65 | reg_act_config_inst_regs_17_sva_dfm_6_enexo_65
      | reg_act_config_inst_counter_enexo_65 | reg_act_regs_data_0_0_2_enexo_4 |
      reg_act_regs_data_2_0_2_enexo_4 | reg_act_regs_data_1_0_2_enexo_4 | reg_act_regs_data_3_0_2_enexo_4);
  assign nv_scvector_cctor_nv_scvector_3_for_and_enex5 = ActUnit_RunInst_switch_lp_and_802_cse
      & (reg_act_config_inst_regs_1_sva_dfm_5_enexo_66 | reg_act_config_inst_regs_17_sva_dfm_6_enexo_66
      | reg_act_regs_data_0_1_2_enexo_4 | reg_act_regs_data_2_1_2_enexo_4 | reg_act_config_inst_counter_enexo_66
      | reg_act_regs_data_1_1_2_enexo_4 | reg_act_regs_data_3_1_2_enexo_4);
  assign nv_scvector_cctor_nv_scvector_3_for_and_15_enex5 = ActUnit_RunInst_switch_lp_and_802_cse
      & (reg_act_config_inst_regs_17_sva_dfm_6_enexo_67 | reg_act_config_inst_regs_1_sva_dfm_5_enexo_67
      | reg_act_regs_data_2_2_2_enexo_4 | reg_act_regs_data_0_2_2_enexo_4 | reg_act_regs_data_1_2_2_enexo_4
      | reg_act_config_inst_counter_enexo_67 | reg_act_regs_data_3_2_2_enexo_4);
  assign nv_scvector_cctor_nv_scvector_3_for_and_16_enex5 = ActUnit_RunInst_switch_lp_and_802_cse
      & (reg_act_config_inst_regs_1_sva_dfm_5_enexo_68 | reg_act_config_inst_regs_17_sva_dfm_6_enexo_68
      | reg_act_regs_data_3_3_2_enexo_4 | reg_act_regs_data_0_3_2_enexo_4 | reg_act_config_inst_counter_enexo_68
      | reg_act_regs_data_2_3_2_enexo_4 | reg_act_regs_data_1_3_2_enexo_4);
  assign nv_scvector_cctor_nv_scvector_3_for_and_17_enex5 = ActUnit_RunInst_switch_lp_and_802_cse
      & (reg_act_config_inst_regs_17_sva_dfm_6_enexo_69 | reg_act_config_inst_regs_1_sva_dfm_5_enexo_69
      | reg_act_config_inst_counter_enexo_69 | reg_act_regs_data_0_4_2_enexo_4 |
      reg_act_regs_data_3_4_2_enexo_4 | reg_act_regs_data_2_4_2_enexo_4 | reg_act_regs_data_1_4_2_enexo_4);
  assign nv_scvector_cctor_nv_scvector_3_for_and_18_enex5 = ActUnit_RunInst_switch_lp_and_802_cse
      & (reg_act_config_inst_regs_17_sva_dfm_6_enexo_70 | reg_act_config_inst_regs_1_sva_dfm_5_enexo_70
      | reg_act_regs_data_2_5_2_enexo_4 | reg_act_config_inst_counter_enexo_70 |
      reg_act_regs_data_1_5_2_enexo_4 | reg_act_regs_data_3_5_2_enexo_4 | reg_act_regs_data_0_5_2_enexo_4);
  assign nv_scvector_cctor_nv_scvector_3_for_and_19_enex5 = ActUnit_RunInst_switch_lp_and_802_cse
      & (reg_act_config_inst_regs_17_sva_dfm_6_enexo_71 | reg_act_config_inst_regs_1_sva_dfm_5_enexo_71
      | reg_act_regs_data_3_6_2_enexo_4 | reg_act_regs_data_1_6_2_enexo_4 | reg_act_config_inst_counter_enexo_71
      | reg_act_regs_data_2_6_2_enexo_4 | reg_act_regs_data_0_6_2_enexo_4);
  assign nv_scvector_cctor_nv_scvector_3_for_and_20_enex5 = ActUnit_RunInst_switch_lp_and_802_cse
      & (reg_act_config_inst_regs_17_sva_dfm_6_enexo_72 | reg_act_config_inst_regs_1_sva_dfm_5_enexo_72
      | reg_act_regs_data_1_7_2_enexo_4 | reg_act_config_inst_counter_enexo_72 |
      reg_act_regs_data_0_7_2_enexo_4 | reg_act_regs_data_2_7_2_enexo_4 | reg_act_regs_data_3_7_2_enexo_4);
  assign nv_scvector_cctor_nv_scvector_3_for_and_21_enex5 = ActUnit_RunInst_switch_lp_and_802_cse
      & (reg_act_config_inst_regs_1_sva_dfm_5_enexo_73 | reg_act_config_inst_regs_17_sva_dfm_6_enexo_73
      | reg_act_regs_data_2_8_2_enexo_4 | reg_act_config_inst_counter_enexo_73 |
      reg_act_regs_data_1_8_2_enexo_4 | reg_act_regs_data_3_8_2_enexo_4 | reg_act_regs_data_0_8_2_enexo_4);
  assign nv_scvector_cctor_nv_scvector_3_for_and_22_enex5 = ActUnit_RunInst_switch_lp_and_802_cse
      & (reg_act_config_inst_regs_1_sva_dfm_5_enexo_74 | reg_act_config_inst_regs_17_sva_dfm_6_enexo_74
      | reg_act_regs_data_0_11_2_enexo_4 | reg_act_regs_data_1_11_2_enexo_4 | reg_act_regs_data_3_11_2_enexo_4
      | reg_act_config_inst_counter_enexo_74 | reg_act_regs_data_2_11_2_enexo_4);
  assign nv_scvector_cctor_nv_scvector_3_for_and_23_enex5 = ActUnit_RunInst_switch_lp_and_802_cse
      & (reg_act_config_inst_regs_1_sva_dfm_5_enexo_75 | reg_act_config_inst_regs_17_sva_dfm_6_enexo_75
      | reg_act_config_inst_counter_enexo_75 | reg_act_regs_data_3_12_2_enexo_4 |
      reg_act_regs_data_1_12_2_enexo_4 | reg_act_regs_data_2_12_2_enexo_4 | reg_act_regs_data_0_12_2_enexo_4);
  assign nv_scvector_cctor_nv_scvector_3_for_and_24_enex5 = ActUnit_RunInst_switch_lp_and_802_cse
      & (reg_act_config_inst_regs_1_sva_dfm_5_enexo_76 | reg_act_config_inst_regs_17_sva_dfm_6_enexo_76
      | reg_act_config_inst_counter_enexo_76 | reg_act_regs_data_1_13_2_enexo_4 |
      reg_act_regs_data_2_13_2_enexo_4 | reg_act_regs_data_0_13_2_enexo_4 | reg_act_regs_data_3_13_2_enexo_4);
  assign nv_scvector_cctor_nv_scvector_3_for_and_25_enex5 = ActUnit_RunInst_switch_lp_and_802_cse
      & (reg_act_config_inst_regs_1_sva_dfm_5_enexo_77 | reg_act_config_inst_regs_17_sva_dfm_6_enexo_77
      | reg_act_regs_data_2_14_2_enexo_4 | reg_act_regs_data_3_14_2_enexo_4 | reg_act_regs_data_0_14_2_enexo_4
      | reg_act_regs_data_1_14_2_enexo_4 | reg_act_config_inst_counter_enexo_77);
  assign or_dcpl_639 = ~(and_dcpl_916 | act_config_ActConfigRead_else_else_not_21);
  assign and_dcpl_1013 = and_dcpl_1001 & (fsm_output[2]);
  assign and_dcpl_1019 = (fsm_output[4:2]==3'b010);
  assign and_dcpl_1021 = (fsm_output[1:0]==2'b01);
  assign and_dcpl_1028 = (fsm_output[4:2]==3'b011);
  assign and_dcpl_1046 = (fsm_output[4:2]==3'b001);
  assign and_1152_cse = and_dcpl_1019 & and_dcpl_563;
  assign and_1156_cse = and_dcpl_1019 & (fsm_output[1:0]==2'b10);
  assign and_1158_cse = and_dcpl_1019 & (fsm_output[1:0]==2'b11);
  assign and_1161_cse = and_dcpl_1028 & and_dcpl_563;
  assign and_1154_cse = and_dcpl_1019 & and_dcpl_1021;
  assign and_1181_cse = and_dcpl_1046 & and_dcpl_1021;
  assign and_1183_cse = and_dcpl_1046 & and_dcpl_570;
  assign and_1185_cse = and_dcpl_1046 & and_1104_cse;
  assign and_1190_cse = and_dcpl_1019 & and_dcpl_570;
  assign and_1191_cse = and_dcpl_1019 & and_1104_cse;
  assign Tanh_for_else_else_and_2_cse = (~ (act_config_in_InstFetch_mux_tmp[6]))
      & and_dcpl_554;
  assign Tanh_for_else_else_and_3_cse = and_dcpl_47 & and_dcpl_554;
  assign mux_92_nl = MUX_s_1_2_2((~ (fsm_output[3])), or_tmp_126, fsm_output[2]);
  assign and_568_nl = (fsm_output[2]) & or_tmp_126;
  assign mux_93_nl = MUX_s_1_2_2(mux_92_nl, and_568_nl, fsm_output[0]);
  assign mux_91_nl = MUX_s_1_2_2((fsm_output[3]), or_tmp_126, or_1071_cse);
  assign mux_94_nl = MUX_s_1_2_2(mux_93_nl, mux_91_nl, fsm_output[1]);
  assign Tanh_for_else_else_or_cse = ((act_config_in_InstFetch_mux_tmp[6]) & (act_config_in_InstFetch_mux_tmp[4])
      & and_dcpl_554) | mux_94_nl | (fsm_output[4]);
  assign or_tmp_421 = ActUnit_RunInst_switch_lp_equal_tmp_4 | ActUnit_RunInst_switch_lp_equal_tmp_5
      | ActUnit_RunInst_switch_lp_equal_tmp_6 | ActUnit_RunInst_switch_lp_equal_tmp_7
      | ActUnit_RunInst_switch_lp_equal_tmp_8;
  assign nand_tmp_13 = ~((~(ActUnit_RunInst_switch_lp_and_tmp & ActUnit_RunInst_switch_lp_equal_tmp_2))
      & is_start_sva & while_nor_itm & (~(or_tmp_421 & reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_nor_cse)));
  assign or_tmp_446 = (fsm_output[4:1]!=4'b0110) | nand_298_cse;
  assign or_tmp_517 = ActUnit_RunInst_switch_lp_equal_tmp_4 | ActUnit_RunInst_switch_lp_equal_tmp_5
      | ActUnit_RunInst_switch_lp_equal_tmp_6 | ActUnit_RunInst_switch_lp_equal_tmp_7;
  assign or_tmp_518 = (ActUnit_PushOutput_if_for_and_stg_2_7_sva & ActUnit_RunInst_switch_lp_equal_tmp_8)
      | (~((~(ActUnit_RunInst_switch_lp_and_16_tmp & ActUnit_RunInst_switch_lp_equal_tmp_2))
      & is_start_sva & while_nor_16_itm & (~(or_tmp_517 & reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_1_cse))));
  assign or_tmp_547 = (fsm_output[4:1]!=4'b0110) | nand_338_cse;
  assign nand_tmp_45 = ~((~(ActUnit_RunInst_switch_lp_and_32_tmp & ActUnit_RunInst_switch_lp_equal_tmp_2))
      & is_start_sva & while_nor_32_itm & (~(or_tmp_421 & reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_cse)));
  assign or_tmp_654 = (fsm_output[4:1]!=4'b0110) | nand_378_cse;
  assign or_tmp_726 = (Gelu_for_and_2_cse_sva & ActUnit_RunInst_switch_lp_equal_tmp_8)
      | (~((~(ActUnit_RunInst_switch_lp_and_48_tmp & ActUnit_RunInst_switch_lp_equal_tmp_2))
      & is_start_sva & while_nor_48_itm & (~(or_tmp_517 & reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_2_cse))));
  assign or_tmp_755 = (fsm_output[4:1]!=4'b0110) | nand_418_cse;
  assign or_dcpl_652 = (and_dcpl_852 & (~ nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_71_0))
      | and_dcpl_554;
  assign and_dcpl_1229 = and_dcpl_852 & (~ nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_67_0);
  assign or_dcpl_655 = and_dcpl_1229 | and_dcpl_997;
  assign w_load_and_tmp = ActUnitRun_wen & ((is_start_sva & (~ or_dcpl_440)) | and_dcpl_554)
      & or_71_cse;
  assign is_start_and_tmp = ActUnitRun_wen & (and_dcpl_768 | and_dcpl_794);
  assign and_1602_nl = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]) & (nvhls_get_slc_2U_NVUINT8_return_3_sva==2'b11)
      & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]) & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3])
      & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign mux_576_nl = MUX_s_1_2_2(or_tmp_755, (~ mux_523_cse), and_1602_nl);
  assign mux_577_nl = MUX_s_1_2_2(mux_576_nl, or_tmp_755, ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]);
  assign and_1417_tmp = (~ mux_577_nl) & ActUnitRun_wen;
  assign mux_564_nl = MUX_s_1_2_2(or_tmp_755, (~ mux_523_cse), and_1485_cse);
  assign or_1495_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b11) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]);
  assign mux_573_nl = MUX_s_1_2_2(mux_564_nl, or_tmp_755, or_1495_nl);
  assign and_1415_tmp = (~ mux_573_nl) & ActUnitRun_wen;
  assign and_1596_nl = (nvhls_get_slc_2U_NVUINT8_return_3_sva==2'b11) & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])
      & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]) & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign mux_568_nl = MUX_s_1_2_2(or_tmp_755, (~ mux_523_cse), and_1596_nl);
  assign mux_569_nl = MUX_s_1_2_2(mux_568_nl, or_tmp_755, or_1488_cse);
  assign and_1413_tmp = (~ mux_569_nl) & ActUnitRun_wen;
  assign mux_622_nl = MUX_s_1_2_2(or_tmp_755, (~ mux_523_cse), and_1485_cse);
  assign or_1481_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b11) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]);
  assign mux_565_nl = MUX_s_1_2_2(mux_622_nl, or_tmp_755, or_1481_nl);
  assign and_1411_tmp = (~ mux_565_nl) & ActUnitRun_wen;
  assign nand_448_nl = ~((~ (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4])) & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      & (nvhls_get_slc_2U_NVUINT8_return_3_sva==2'b11) & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])
      & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]) & (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2])));
  assign mux_561_nl = MUX_s_1_2_2(mux_523_cse, nor_760_cse, nand_448_nl);
  assign and_1409_tmp = mux_561_nl & ActUnitRun_wen;
  assign or_1467_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b11) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])
      | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign mux_558_nl = MUX_s_1_2_2(mux_523_cse, nor_760_cse, or_1467_nl);
  assign and_1407_tmp = mux_558_nl & ActUnitRun_wen;
  assign or_1460_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b11) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]))
      | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign mux_555_nl = MUX_s_1_2_2(mux_523_cse, nor_760_cse, or_1460_nl);
  assign and_1405_tmp = mux_555_nl & ActUnitRun_wen;
  assign or_1453_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b11) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])
      | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign mux_552_nl = MUX_s_1_2_2(mux_523_cse, nor_760_cse, or_1453_nl);
  assign and_1403_tmp = mux_552_nl & ActUnitRun_wen;
  assign mux_540_nl = MUX_s_1_2_2(or_tmp_755, (~ mux_523_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign or_1446_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b11) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_549_nl = MUX_s_1_2_2(mux_540_nl, or_tmp_755, or_1446_nl);
  assign and_1401_tmp = (~ mux_549_nl) & ActUnitRun_wen;
  assign mux_621_nl = MUX_s_1_2_2(or_tmp_755, (~ mux_523_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign or_1439_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b11) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_545_nl = MUX_s_1_2_2(mux_621_nl, or_tmp_755, or_1439_nl);
  assign and_1399_tmp = (~ mux_545_nl) & ActUnitRun_wen;
  assign mux_620_nl = MUX_s_1_2_2(or_tmp_755, (~ mux_523_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign or_1432_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b11) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_541_nl = MUX_s_1_2_2(mux_620_nl, or_tmp_755, or_1432_nl);
  assign and_1397_tmp = (~ mux_541_nl) & ActUnitRun_wen;
  assign mux_536_nl = MUX_s_1_2_2(or_tmp_755, (~ mux_523_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign or_1425_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b11) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_537_nl = MUX_s_1_2_2(mux_536_nl, or_tmp_755, or_1425_nl);
  assign and_1395_tmp = (~ mux_537_nl) & ActUnitRun_wen;
  assign or_1418_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b11) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign mux_533_nl = MUX_s_1_2_2(mux_523_cse, nor_760_cse, or_1418_nl);
  assign and_1393_tmp = mux_533_nl & ActUnitRun_wen;
  assign or_1411_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b11) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign mux_530_nl = MUX_s_1_2_2(mux_523_cse, nor_760_cse, or_1411_nl);
  assign and_1391_tmp = mux_530_nl & ActUnitRun_wen;
  assign or_1404_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b11) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign mux_527_nl = MUX_s_1_2_2(mux_523_cse, nor_760_cse, or_1404_nl);
  assign and_1389_tmp = mux_527_nl & ActUnitRun_wen;
  assign or_1397_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b11) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign mux_524_nl = MUX_s_1_2_2(mux_523_cse, nor_760_cse, or_1397_nl);
  assign and_1387_tmp = mux_524_nl & ActUnitRun_wen;
  assign mux_512_nl = MUX_s_1_2_2(or_tmp_654, (~ mux_467_cse), and_1876_cse);
  assign or_1391_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]);
  assign mux_521_nl = MUX_s_1_2_2(mux_512_nl, or_tmp_654, or_1391_nl);
  assign and_1385_tmp = (~ mux_521_nl) & ActUnitRun_wen;
  assign mux_508_nl = MUX_s_1_2_2(or_tmp_654, (~ mux_467_cse), and_1485_cse);
  assign or_1385_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b10) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]);
  assign mux_517_nl = MUX_s_1_2_2(mux_508_nl, or_tmp_654, or_1385_nl);
  assign and_1383_tmp = (~ mux_517_nl) & ActUnitRun_wen;
  assign mux_619_nl = MUX_s_1_2_2(or_tmp_654, (~ mux_467_cse), and_1876_cse);
  assign or_1379_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]);
  assign mux_513_nl = MUX_s_1_2_2(mux_619_nl, or_tmp_654, or_1379_nl);
  assign and_1381_tmp = (~ mux_513_nl) & ActUnitRun_wen;
  assign mux_618_nl = MUX_s_1_2_2(or_tmp_654, (~ mux_467_cse), and_1485_cse);
  assign or_1373_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b10) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]);
  assign mux_509_nl = MUX_s_1_2_2(mux_618_nl, or_tmp_654, or_1373_nl);
  assign and_1379_tmp = (~ mux_509_nl) & ActUnitRun_wen;
  assign or_1367_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b10) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]))
      | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign mux_505_nl = MUX_s_1_2_2(mux_467_cse, nor_752_cse, or_1367_nl);
  assign and_1377_tmp = mux_505_nl & ActUnitRun_wen;
  assign or_1361_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b10) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])
      | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign mux_502_nl = MUX_s_1_2_2(mux_467_cse, nor_752_cse, or_1361_nl);
  assign and_1375_tmp = mux_502_nl & ActUnitRun_wen;
  assign or_1355_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b10) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]))
      | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign mux_499_nl = MUX_s_1_2_2(mux_467_cse, nor_752_cse, or_1355_nl);
  assign and_1373_tmp = mux_499_nl & ActUnitRun_wen;
  assign or_1349_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b10) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])
      | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign mux_496_nl = MUX_s_1_2_2(mux_467_cse, nor_752_cse, or_1349_nl);
  assign and_1371_tmp = mux_496_nl & ActUnitRun_wen;
  assign mux_484_nl = MUX_s_1_2_2(or_tmp_654, (~ mux_467_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign or_1343_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b10) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_493_nl = MUX_s_1_2_2(mux_484_nl, or_tmp_654, or_1343_nl);
  assign and_1369_tmp = (~ mux_493_nl) & ActUnitRun_wen;
  assign mux_617_nl = MUX_s_1_2_2(or_tmp_654, (~ mux_467_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign or_1337_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b10) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_489_nl = MUX_s_1_2_2(mux_617_nl, or_tmp_654, or_1337_nl);
  assign and_1367_tmp = (~ mux_489_nl) & ActUnitRun_wen;
  assign mux_616_nl = MUX_s_1_2_2(or_tmp_654, (~ mux_467_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign or_1331_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b10) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_485_nl = MUX_s_1_2_2(mux_616_nl, or_tmp_654, or_1331_nl);
  assign and_1365_tmp = (~ mux_485_nl) & ActUnitRun_wen;
  assign mux_480_nl = MUX_s_1_2_2(or_tmp_654, (~ mux_467_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign or_1325_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b10) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_481_nl = MUX_s_1_2_2(mux_480_nl, or_tmp_654, or_1325_nl);
  assign and_1363_tmp = (~ mux_481_nl) & ActUnitRun_wen;
  assign or_1319_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b10) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign mux_477_nl = MUX_s_1_2_2(mux_467_cse, nor_752_cse, or_1319_nl);
  assign and_1361_tmp = mux_477_nl & ActUnitRun_wen;
  assign or_1313_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b10) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign mux_474_nl = MUX_s_1_2_2(mux_467_cse, nor_752_cse, or_1313_nl);
  assign and_1359_tmp = mux_474_nl & ActUnitRun_wen;
  assign or_1307_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b10) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign mux_471_nl = MUX_s_1_2_2(mux_467_cse, nor_752_cse, or_1307_nl);
  assign and_1357_tmp = mux_471_nl & ActUnitRun_wen;
  assign or_1301_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b10) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign mux_468_nl = MUX_s_1_2_2(mux_467_cse, nor_752_cse, or_1301_nl);
  assign and_1355_tmp = mux_468_nl & ActUnitRun_wen;
  assign mux_456_nl = MUX_s_1_2_2(or_tmp_547, (~ mux_411_cse), and_1488_cse);
  assign or_1294_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b01);
  assign mux_465_nl = MUX_s_1_2_2(mux_456_nl, or_tmp_547, or_1294_nl);
  assign and_1353_tmp = (~ mux_465_nl) & ActUnitRun_wen;
  assign mux_452_nl = MUX_s_1_2_2(or_tmp_547, (~ mux_411_cse), and_1485_cse);
  assign or_1287_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b01) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]);
  assign mux_461_nl = MUX_s_1_2_2(mux_452_nl, or_tmp_547, or_1287_nl);
  assign and_1351_tmp = (~ mux_461_nl) & ActUnitRun_wen;
  assign mux_615_nl = MUX_s_1_2_2(or_tmp_547, (~ mux_411_cse), and_1488_cse);
  assign or_1280_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b01);
  assign mux_457_nl = MUX_s_1_2_2(mux_615_nl, or_tmp_547, or_1280_nl);
  assign and_1349_tmp = (~ mux_457_nl) & ActUnitRun_wen;
  assign mux_614_nl = MUX_s_1_2_2(or_tmp_547, (~ mux_411_cse), and_1485_cse);
  assign or_1273_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b01) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]);
  assign mux_453_nl = MUX_s_1_2_2(mux_614_nl, or_tmp_547, or_1273_nl);
  assign and_1347_tmp = (~ mux_453_nl) & ActUnitRun_wen;
  assign or_1266_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b01) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]))
      | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign mux_449_nl = MUX_s_1_2_2(mux_411_cse, nor_744_cse, or_1266_nl);
  assign and_1345_tmp = mux_449_nl & ActUnitRun_wen;
  assign or_1259_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b01) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])
      | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign mux_446_nl = MUX_s_1_2_2(mux_411_cse, nor_744_cse, or_1259_nl);
  assign and_1343_tmp = mux_446_nl & ActUnitRun_wen;
  assign or_1252_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b01) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]))
      | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign mux_443_nl = MUX_s_1_2_2(mux_411_cse, nor_744_cse, or_1252_nl);
  assign and_1341_tmp = mux_443_nl & ActUnitRun_wen;
  assign or_1245_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b01) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])
      | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign mux_440_nl = MUX_s_1_2_2(mux_411_cse, nor_744_cse, or_1245_nl);
  assign and_1339_tmp = mux_440_nl & ActUnitRun_wen;
  assign mux_428_nl = MUX_s_1_2_2(or_tmp_547, (~ mux_411_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign or_1238_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b01) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_437_nl = MUX_s_1_2_2(mux_428_nl, or_tmp_547, or_1238_nl);
  assign and_1337_tmp = (~ mux_437_nl) & ActUnitRun_wen;
  assign mux_613_nl = MUX_s_1_2_2(or_tmp_547, (~ mux_411_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign or_1231_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b01) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_433_nl = MUX_s_1_2_2(mux_613_nl, or_tmp_547, or_1231_nl);
  assign and_1335_tmp = (~ mux_433_nl) & ActUnitRun_wen;
  assign mux_612_nl = MUX_s_1_2_2(or_tmp_547, (~ mux_411_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign or_1224_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b01) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_429_nl = MUX_s_1_2_2(mux_612_nl, or_tmp_547, or_1224_nl);
  assign and_1333_tmp = (~ mux_429_nl) & ActUnitRun_wen;
  assign mux_424_nl = MUX_s_1_2_2(or_tmp_547, (~ mux_411_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign or_1217_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b01) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_425_nl = MUX_s_1_2_2(mux_424_nl, or_tmp_547, or_1217_nl);
  assign and_1331_tmp = (~ mux_425_nl) & ActUnitRun_wen;
  assign or_1210_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b01) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign mux_421_nl = MUX_s_1_2_2(mux_411_cse, nor_744_cse, or_1210_nl);
  assign and_1329_tmp = mux_421_nl & ActUnitRun_wen;
  assign or_1203_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b01) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign mux_418_nl = MUX_s_1_2_2(mux_411_cse, nor_744_cse, or_1203_nl);
  assign and_1327_tmp = mux_418_nl & ActUnitRun_wen;
  assign or_1196_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b01) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign mux_415_nl = MUX_s_1_2_2(mux_411_cse, nor_744_cse, or_1196_nl);
  assign and_1325_tmp = mux_415_nl & ActUnitRun_wen;
  assign or_1189_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b01) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign mux_412_nl = MUX_s_1_2_2(mux_411_cse, nor_744_cse, or_1189_nl);
  assign and_1323_tmp = mux_412_nl & ActUnitRun_wen;
  assign or_1078_nl = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0!=4'b0010);
  assign mux_349_nl = MUX_s_1_2_2(mux_342_cse, mux_344_cse, or_1078_nl);
  assign and_1246_tmp = mux_349_nl & (fsm_output[4:3]==2'b01) & ActUnitRun_wen;
  assign mux_400_nl = MUX_s_1_2_2(or_tmp_446, (~ mux_355_cse), and_1488_cse);
  assign or_1183_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b00);
  assign mux_409_nl = MUX_s_1_2_2(mux_400_nl, or_tmp_446, or_1183_nl);
  assign and_1321_tmp = (~ mux_409_nl) & ActUnitRun_wen;
  assign and_1456_nl = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0==4'b1110);
  assign mux_345_nl = MUX_s_1_2_2(mux_344_cse, mux_342_cse, and_1456_nl);
  assign and_1243_tmp = mux_345_nl & (fsm_output[4:3]==2'b01) & ActUnitRun_wen;
  assign mux_396_nl = MUX_s_1_2_2(or_tmp_446, (~ mux_355_cse), and_1485_cse);
  assign or_1177_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b00) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]);
  assign mux_405_nl = MUX_s_1_2_2(mux_396_nl, or_tmp_446, or_1177_nl);
  assign and_1319_tmp = (~ mux_405_nl) & ActUnitRun_wen;
  assign and_1454_nl = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0==4'b1101);
  assign mux_338_nl = MUX_s_1_2_2(mux_337_cse, mux_336_cse, and_1454_nl);
  assign and_1237_tmp = mux_338_nl & (fsm_output[4:3]==2'b01) & ActUnitRun_wen;
  assign mux_611_nl = MUX_s_1_2_2(or_tmp_446, (~ mux_355_cse), and_1488_cse);
  assign or_1171_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b00);
  assign mux_401_nl = MUX_s_1_2_2(mux_611_nl, or_tmp_446, or_1171_nl);
  assign and_1317_tmp = (~ mux_401_nl) & ActUnitRun_wen;
  assign nor_362_nl = ~((ActUnit_PushOutput_if_for_i_4_0_sva_3_0!=4'b1100));
  assign mux_331_nl = MUX_s_1_2_2(mux_330_cse, mux_328_cse, nor_362_nl);
  assign and_1231_tmp = mux_331_nl & (fsm_output[4:3]==2'b01) & ActUnitRun_wen;
  assign mux_610_nl = MUX_s_1_2_2(or_tmp_446, (~ mux_355_cse), and_1485_cse);
  assign or_1165_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b00) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]);
  assign mux_397_nl = MUX_s_1_2_2(mux_610_nl, or_tmp_446, or_1165_nl);
  assign and_1315_tmp = (~ mux_397_nl) & ActUnitRun_wen;
  assign and_1275_tmp = (((ActUnit_PushOutput_if_for_i_4_0_sva_3_0==4'b1011)) | (fsm_output[1:0]!=2'b10))
      & (fsm_output[4:2]==3'b011) & ActUnitRun_wen;
  assign or_1159_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b00) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]))
      | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign mux_393_nl = MUX_s_1_2_2(mux_355_cse, nor_736_cse, or_1159_nl);
  assign and_1313_tmp = mux_393_nl & ActUnitRun_wen;
  assign and_1268_tmp = (((ActUnit_PushOutput_if_for_i_4_0_sva_3_0==4'b1010)) | (fsm_output[1:0]!=2'b10))
      & (fsm_output[4:2]==3'b011) & ActUnitRun_wen;
  assign or_1153_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b00) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])
      | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign mux_390_nl = MUX_s_1_2_2(mux_355_cse, nor_736_cse, or_1153_nl);
  assign and_1311_tmp = mux_390_nl & ActUnitRun_wen;
  assign or_1147_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b00) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]))
      | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign mux_387_nl = MUX_s_1_2_2(mux_355_cse, nor_736_cse, or_1147_nl);
  assign and_1309_tmp = mux_387_nl & ActUnitRun_wen;
  assign or_1076_nl = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0!=4'b1001);
  assign mux_341_nl = MUX_s_1_2_2(mux_336_cse, mux_337_cse, or_1076_nl);
  assign and_1240_tmp = mux_341_nl & (fsm_output[4:3]==2'b01) & ActUnitRun_wen;
  assign or_1141_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b00) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])
      | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign mux_384_nl = MUX_s_1_2_2(mux_355_cse, nor_736_cse, or_1141_nl);
  assign and_1307_tmp = mux_384_nl & ActUnitRun_wen;
  assign or_1074_nl = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0!=4'b1000);
  assign mux_335_nl = MUX_s_1_2_2(mux_328_cse, mux_330_cse, or_1074_nl);
  assign and_1234_tmp = mux_335_nl & (fsm_output[4:3]==2'b01) & ActUnitRun_wen;
  assign mux_372_nl = MUX_s_1_2_2(or_tmp_446, (~ mux_355_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign or_1135_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b00) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_381_nl = MUX_s_1_2_2(mux_372_nl, or_tmp_446, or_1135_nl);
  assign and_1305_tmp = (~ mux_381_nl) & ActUnitRun_wen;
  assign mux_325_nl = MUX_s_1_2_2((~ (fsm_output[3])), (fsm_output[3]), fsm_output[0]);
  assign and_1449_nl = (fsm_output[0]) & (fsm_output[3]);
  assign mux_326_nl = MUX_s_1_2_2(mux_325_nl, and_1449_nl, fsm_output[1]);
  assign mux_324_nl = MUX_s_1_2_2((~ (fsm_output[3])), (fsm_output[3]), or_992_cse);
  assign and_1450_nl = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0==4'b0111);
  assign mux_327_nl = MUX_s_1_2_2(mux_326_nl, mux_324_nl, and_1450_nl);
  assign and_1228_tmp = mux_327_nl & (fsm_output[2]) & (~ (fsm_output[4])) & ActUnitRun_wen;
  assign mux_609_nl = MUX_s_1_2_2(or_tmp_446, (~ mux_355_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign or_1129_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b00) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_377_nl = MUX_s_1_2_2(mux_609_nl, or_tmp_446, or_1129_nl);
  assign and_1303_tmp = (~ mux_377_nl) & ActUnitRun_wen;
  assign and_1289_tmp = (((ActUnit_PushOutput_if_for_i_4_0_sva_3_0==4'b0110)) | (fsm_output[1:0]!=2'b10))
      & (fsm_output[4:2]==3'b011) & ActUnitRun_wen;
  assign mux_608_nl = MUX_s_1_2_2(or_tmp_446, (~ mux_355_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign or_1123_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b00) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_373_nl = MUX_s_1_2_2(mux_608_nl, or_tmp_446, or_1123_nl);
  assign and_1301_tmp = (~ mux_373_nl) & ActUnitRun_wen;
  assign and_1282_tmp = (((ActUnit_PushOutput_if_for_i_4_0_sva_3_0==4'b0101)) | (fsm_output[1:0]!=2'b10))
      & (fsm_output[4:2]==3'b011) & ActUnitRun_wen;
  assign mux_368_nl = MUX_s_1_2_2(or_tmp_446, (~ mux_355_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign or_1117_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b00) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_369_nl = MUX_s_1_2_2(mux_368_nl, or_tmp_446, or_1117_nl);
  assign and_1299_tmp = (~ mux_369_nl) & ActUnitRun_wen;
  assign nor_372_nl = ~((ActUnit_PushOutput_if_for_i_4_0_sva_3_0!=4'b0100));
  assign mux_353_nl = MUX_s_1_2_2(and_1249_cse, mux_350_cse, nor_372_nl);
  assign and_1254_tmp = mux_353_nl & (fsm_output[4:3]==2'b01) & ActUnitRun_wen;
  assign or_1111_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b00) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign mux_365_nl = MUX_s_1_2_2(mux_355_cse, nor_736_cse, or_1111_nl);
  assign and_1297_tmp = mux_365_nl & ActUnitRun_wen;
  assign or_1080_nl = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0!=4'b0011);
  assign mux_351_nl = MUX_s_1_2_2(mux_350_cse, and_1249_cse, or_1080_nl);
  assign and_1250_tmp = mux_351_nl & (fsm_output[4:3]==2'b01) & ActUnitRun_wen;
  assign or_1105_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b00) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign mux_362_nl = MUX_s_1_2_2(mux_355_cse, nor_736_cse, or_1105_nl);
  assign and_1295_tmp = mux_362_nl & ActUnitRun_wen;
  assign and_1261_tmp = (((ActUnit_PushOutput_if_for_i_4_0_sva_3_0==4'b0001)) | (fsm_output[1:0]!=2'b10))
      & (fsm_output[4:2]==3'b011) & ActUnitRun_wen;
  assign or_1099_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b00) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign mux_359_nl = MUX_s_1_2_2(mux_355_cse, nor_736_cse, or_1099_nl);
  assign and_1293_tmp = mux_359_nl & ActUnitRun_wen;
  assign mux_322_nl = MUX_s_1_2_2((~ (fsm_output[3])), (fsm_output[3]), or_1071_cse);
  assign mux_321_nl = MUX_s_1_2_2(nor_734_cse, (fsm_output[3]), fsm_output[0]);
  assign or_1069_nl = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0!=4'b0000);
  assign mux_323_nl = MUX_s_1_2_2(mux_322_nl, mux_321_nl, or_1069_nl);
  assign and_1225_tmp = mux_323_nl & (fsm_output[1]) & (~ (fsm_output[4])) & ActUnitRun_wen;
  assign or_1093_nl = (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b00) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign mux_356_nl = MUX_s_1_2_2(mux_355_cse, nor_736_cse, or_1093_nl);
  assign and_1291_tmp = mux_356_nl & ActUnitRun_wen;
  assign or_991_nl = and_1108_cse | (fsm_output[3]);
  assign mux_221_nl = MUX_s_1_2_2(or_991_nl, nor_333_cse, fsm_output[4]);
  assign ActUnit_CheckStart_start_reg_and_tmp = ActUnitRun_wen & (~ mux_221_nl);
  assign act_config_inst_counter_and_tmp = ActUnitRun_wen & ((and_dcpl_746 & (~((fsm_output[2])
      | (fsm_output[0]))) & and_dcpl_789 & is_incr_lpi_1_dfm_1) | act_config_inst_counter_sva_mx0c1);
  assign ActUnit_PushOutput_if_for_and_27_itm = ActUnit_PushOutput_if_for_and_stg_2_7_sva
      & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign Tanh_for_else_else_and_8_cse = (~ (act_config_in_InstFetch_mux_tmp[4]))
      & and_dcpl_554;
  assign Tanh_for_else_else_and_9_cse = (act_config_in_InstFetch_mux_tmp[4]) & and_dcpl_554;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Tanh_for_1_else_else_mul_1_cmp_cgo_ir_1_cse <= 1'b0;
      reg_Tanh_for_1_else_else_mul_1_cmp_cgo_ir_cse <= 1'b0;
      reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_15_cse <= 1'b0;
      reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_14_cse <= 1'b0;
      reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_13_cse <= 1'b0;
      reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_12_cse <= 1'b0;
      reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_11_cse <= 1'b0;
      reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_10_cse <= 1'b0;
      reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_9_cse <= 1'b0;
      reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_8_cse <= 1'b0;
      reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_7_cse <= 1'b0;
      reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_6_cse <= 1'b0;
      reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_5_cse <= 1'b0;
      reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_4_cse <= 1'b0;
      reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_3_cse <= 1'b0;
      reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_2_cse <= 1'b0;
      reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_1_cse <= 1'b0;
      reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_cse <= 1'b0;
      reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_15_cse <= 1'b0;
      reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_14_cse <= 1'b0;
      reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_13_cse <= 1'b0;
      reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_12_cse <= 1'b0;
      reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_11_cse <= 1'b0;
      reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_10_cse <= 1'b0;
      reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_9_cse <= 1'b0;
      reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_8_cse <= 1'b0;
      reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_7_cse <= 1'b0;
      reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_6_cse <= 1'b0;
      reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_5_cse <= 1'b0;
      reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_4_cse <= 1'b0;
      reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_3_cse <= 1'b0;
      reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_2_cse <= 1'b0;
      reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_1_cse <= 1'b0;
      reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_cse <= 1'b0;
      reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_13_cse <= 1'b0;
      reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_12_cse <= 1'b0;
      reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_11_cse <= 1'b0;
      reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_10_cse <= 1'b0;
      reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_9_cse <= 1'b0;
      reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_8_cse <= 1'b0;
      reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_7_cse <= 1'b0;
      reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_6_cse <= 1'b0;
      reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_5_cse <= 1'b0;
      reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_4_cse <= 1'b0;
      reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_3_cse <= 1'b0;
      reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_2_cse <= 1'b0;
      reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_1_cse <= 1'b0;
      reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_cse <= 1'b0;
      reg_done_Push_mioi_iswt0_cse <= 1'b0;
      reg_output_port_Push_mioi_iswt0_cse <= 1'b0;
      reg_start_PopNB_mioi_iswt0_cse <= 1'b0;
      reg_rva_out_Push_mioi_iswt0_cse <= 1'b0;
      reg_act_port_PopNB_mioi_iswt0_cse <= 1'b0;
      reg_rva_in_PopNB_mioi_iswt0_cse <= 1'b0;
      ActUnit_RunInst_switch_lp_nor_tmp <= 1'b0;
    end
    else if ( ActUnitRun_wen ) begin
      reg_Tanh_for_1_else_else_mul_1_cmp_cgo_ir_1_cse <= and_605_rmff;
      reg_Tanh_for_1_else_else_mul_1_cmp_cgo_ir_cse <= and_617_rmff;
      reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_15_cse <= and_621_rmff;
      reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_14_cse <= and_626_rmff;
      reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_13_cse <= and_633_rmff;
      reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_12_cse <= and_658_rmff;
      reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_11_cse <= and_665_rmff;
      reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_10_cse <= and_669_rmff;
      reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_9_cse <= and_673_rmff;
      reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_8_cse <= and_677_rmff;
      reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_7_cse <= and_681_rmff;
      reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_6_cse <= and_685_rmff;
      reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_5_cse <= and_689_rmff;
      reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_4_cse <= and_693_rmff;
      reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_3_cse <= and_697_rmff;
      reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_2_cse <= and_701_rmff;
      reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_1_cse <= and_705_rmff;
      reg_Tanh_for_1_else_else_mul_cmp_cgo_ir_cse <= and_713_rmff;
      reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_15_cse <= and_719_rmff;
      reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_14_cse <= and_724_rmff;
      reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_13_cse <= and_729_rmff;
      reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_12_cse <= and_734_rmff;
      reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_11_cse <= and_739_rmff;
      reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_10_cse <= and_744_rmff;
      reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_9_cse <= and_749_rmff;
      reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_8_cse <= and_754_rmff;
      reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_7_cse <= and_759_rmff;
      reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_6_cse <= and_764_rmff;
      reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_5_cse <= and_769_rmff;
      reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_4_cse <= and_774_rmff;
      reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_3_cse <= and_779_rmff;
      reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_2_cse <= and_784_rmff;
      reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_1_cse <= and_789_rmff;
      reg_Tanh_for_1_else_else_Tanh_for_else_else_mul_cmp_cgo_ir_cse <= and_794_rmff;
      reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_13_cse <= and_799_rmff;
      reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_12_cse <= and_800_rmff;
      reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_11_cse <= and_801_rmff;
      reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_10_cse <= and_802_rmff;
      reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_9_cse <= and_803_rmff;
      reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_8_cse <= and_804_rmff;
      reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_7_cse <= and_805_rmff;
      reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_6_cse <= and_806_rmff;
      reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_5_cse <= and_807_rmff;
      reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_4_cse <= and_808_rmff;
      reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_3_cse <= and_809_rmff;
      reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_2_cse <= and_810_rmff;
      reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_1_cse <= and_811_rmff;
      reg_Tanh_for_3_else_else_mul_1_cmp_cgo_ir_cse <= and_812_rmff;
      reg_done_Push_mioi_iswt0_cse <= and_819_rmff;
      reg_output_port_Push_mioi_iswt0_cse <= and_823_rmff;
      reg_start_PopNB_mioi_iswt0_cse <= and_826_rmff;
      reg_rva_out_Push_mioi_iswt0_cse <= and_830_rmff;
      reg_act_port_PopNB_mioi_iswt0_cse <= and_835_rmff;
      reg_rva_in_PopNB_mioi_iswt0_cse <= and_837_rmff;
      ActUnit_RunInst_switch_lp_nor_tmp <= ActUnit_RunInst_switch_lp_nor_tmp_mx0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_config_is_zero_first_sva <= 1'b0;
    end
    else if ( ActUnitRun_wen & (fsm_output[4]) ) begin
      act_config_is_zero_first_sva <= MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
          while_else_1_mux_1_itm, and_843_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva
          <= 1'b0;
      ActUnit_DecodeAxi_rva_in_reg_rw_sva <= 1'b0;
    end
    else if ( ActUnit_DecodeAxi_if_and_37_cse ) begin
      ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva
          <= ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_mx1;
      ActUnit_DecodeAxi_rva_in_reg_rw_sva <= ActUnit_DecodeAxi_rva_in_reg_rw_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      is_start_sva <= 1'b0;
    end
    else if ( is_start_and_tmp ) begin
      is_start_sva <= MUX_s_1_2_2(while_else_1_while_else_1_nand_1_nl, ActUnit_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva,
          and_dcpl_794);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_DecodeAxiRead_else_unequal_tmp <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_301 | or_dcpl_299)) ) begin
      ActUnit_DecodeAxiRead_else_unequal_tmp <= ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_DecodeAxiWrite_else_unequal_tmp <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_304 | or_dcpl_299)) ) begin
      ActUnit_DecodeAxiWrite_else_unequal_tmp <= ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_config_inst_regs_0_sva_0 <= 1'b0;
      act_config_inst_regs_16_sva_0 <= 1'b0;
      act_config_inst_regs_1_sva_0 <= 1'b0;
      act_config_inst_regs_17_sva_0 <= 1'b0;
    end
    else if ( act_config_inst_regs_and_36_cse ) begin
      act_config_inst_regs_0_sva_0 <= act_config_inst_regs_0_sva_dfm_5[0];
      act_config_inst_regs_16_sva_0 <= act_config_inst_regs_16_sva_dfm_6[0];
      act_config_inst_regs_1_sva_0 <= act_config_inst_regs_1_sva_dfm_5[0];
      act_config_inst_regs_17_sva_0 <= act_config_inst_regs_17_sva_dfm_6[0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_config_num_inst_sva <= 6'b000001;
      act_config_num_output_sva <= 8'b00000001;
      act_config_buffer_addr_base_sva <= 5'b00000;
      act_config_output_addr_base_sva <= 8'b00000000;
    end
    else if ( act_config_num_inst_and_cse ) begin
      act_config_num_inst_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[29:24];
      act_config_num_output_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[39:32];
      act_config_buffer_addr_base_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[52:48];
      act_config_output_addr_base_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[71:64];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_config_is_valid_sva <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~(act_config_ActConfigRead_unequal_tmp_1 | ActUnit_DecodeAxiRead_unequal_tmp_1
        | or_dcpl_303 | or_dcpl_297 | or_1077_cse | or_dcpl_322)) ) begin
      act_config_is_valid_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_29_24_sva_dfm_6 <= 6'b000000;
      rva_out_reg_data_39_32_sva_dfm_6 <= 8'b00000000;
      rva_out_reg_data_52_48_sva_dfm_6 <= 5'b00000;
      rva_out_reg_data_71_64_sva_dfm_6 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_cse ) begin
      rva_out_reg_data_29_24_sva_dfm_6 <= MUX_v_6_2_2((act_mem_banks_read_read_data_lpi_1_dfm_1_31_0[29:24]),
          rva_out_reg_data_29_24_sva_dfm_3, and_dcpl_805);
      rva_out_reg_data_39_32_sva_dfm_6 <= MUX_v_8_2_2((act_mem_banks_read_read_data_lpi_1_dfm_1_63_32[7:0]),
          rva_out_reg_data_39_32_sva_dfm_3, and_dcpl_805);
      rva_out_reg_data_52_48_sva_dfm_6 <= MUX_v_5_2_2((act_mem_banks_read_read_data_lpi_1_dfm_1_63_32[20:16]),
          rva_out_reg_data_52_48_sva_dfm_3, and_dcpl_805);
      rva_out_reg_data_71_64_sva_dfm_6 <= MUX_v_8_2_2((act_mem_banks_read_read_data_lpi_1_dfm_1_95_64[7:0]),
          rva_out_reg_data_71_64_sva_dfm_3, and_dcpl_805);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_0_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_0_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_0_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_0_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_0_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_0_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_0_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_0_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_0_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_0_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_0_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_0_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_0_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_0_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_0_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_0_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_cse ) begin
      act_mem_banks_bank_a_0_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_0_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_0_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_0_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_0_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_0_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_0_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_0_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_0_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_0_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_0_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_0_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_0_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_0_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_0_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_0_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_1_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_1_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_1_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_1_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_1_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_1_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_1_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_1_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_1_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_1_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_1_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_1_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_1_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_1_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_1_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_1_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_1_cse ) begin
      act_mem_banks_bank_a_1_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_1_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_1_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_1_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_1_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_1_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_1_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_1_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_1_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_1_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_1_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_1_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_1_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_1_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_1_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_1_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_2_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_2_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_2_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_2_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_2_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_2_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_2_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_2_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_2_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_2_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_2_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_2_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_2_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_2_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_2_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_2_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_2_cse ) begin
      act_mem_banks_bank_a_2_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_2_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_2_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_2_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_2_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_2_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_2_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_2_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_2_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_2_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_2_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_2_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_2_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_2_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_2_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_2_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_3_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_3_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_3_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_3_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_3_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_3_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_3_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_3_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_3_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_3_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_3_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_3_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_3_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_3_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_3_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_3_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_3_cse ) begin
      act_mem_banks_bank_a_3_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_3_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_3_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_3_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_3_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_3_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_3_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_3_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_3_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_3_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_3_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_3_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_3_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_3_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_3_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_3_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_4_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_4_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_4_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_4_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_4_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_4_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_4_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_4_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_4_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_4_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_4_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_4_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_4_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_4_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_4_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_4_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_4_cse ) begin
      act_mem_banks_bank_a_4_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_4_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_4_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_4_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_4_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_4_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_4_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_4_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_4_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_4_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_4_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_4_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_4_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_4_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_4_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_4_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_5_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_5_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_5_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_5_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_5_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_5_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_5_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_5_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_5_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_5_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_5_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_5_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_5_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_5_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_5_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_5_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_5_cse ) begin
      act_mem_banks_bank_a_5_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_5_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_5_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_5_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_5_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_5_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_5_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_5_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_5_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_5_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_5_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_5_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_5_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_5_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_5_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_5_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_6_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_6_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_6_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_6_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_6_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_6_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_6_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_6_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_6_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_6_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_6_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_6_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_6_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_6_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_6_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_6_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_6_cse ) begin
      act_mem_banks_bank_a_6_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_6_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_6_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_6_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_6_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_6_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_6_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_6_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_6_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_6_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_6_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_6_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_6_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_6_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_6_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_6_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_7_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_7_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_7_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_7_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_7_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_7_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_7_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_7_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_7_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_7_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_7_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_7_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_7_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_7_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_7_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_7_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_7_cse ) begin
      act_mem_banks_bank_a_7_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_7_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_7_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_7_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_7_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_7_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_7_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_7_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_7_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_7_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_7_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_7_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_7_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_7_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_7_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_7_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_8_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_8_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_8_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_8_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_8_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_8_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_8_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_8_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_8_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_8_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_8_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_8_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_8_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_8_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_8_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_8_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_8_cse ) begin
      act_mem_banks_bank_a_8_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_8_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_8_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_8_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_8_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_8_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_8_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_8_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_8_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_8_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_8_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_8_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_8_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_8_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_8_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_8_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_9_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_9_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_9_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_9_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_9_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_9_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_9_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_9_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_9_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_9_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_9_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_9_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_9_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_9_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_9_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_9_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_9_cse ) begin
      act_mem_banks_bank_a_9_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_9_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_9_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_9_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_9_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_9_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_9_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_9_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_9_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_9_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_9_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_9_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_9_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_9_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_9_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_9_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_10_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_10_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_10_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_10_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_10_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_10_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_10_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_10_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_10_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_10_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_10_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_10_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_10_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_10_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_10_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_10_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_10_cse ) begin
      act_mem_banks_bank_a_10_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_10_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_10_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_10_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_10_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_10_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_10_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_10_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_10_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_10_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_10_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_10_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_10_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_10_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_10_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_10_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_11_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_11_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_11_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_11_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_11_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_11_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_11_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_11_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_11_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_11_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_11_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_11_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_11_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_11_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_11_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_11_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_11_cse ) begin
      act_mem_banks_bank_a_11_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_11_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_11_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_11_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_11_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_11_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_11_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_11_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_11_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_11_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_11_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_11_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_11_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_11_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_11_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_11_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_12_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_12_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_12_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_12_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_12_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_12_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_12_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_12_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_12_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_12_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_12_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_12_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_12_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_12_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_12_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_12_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_12_cse ) begin
      act_mem_banks_bank_a_12_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_12_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_12_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_12_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_12_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_12_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_12_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_12_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_12_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_12_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_12_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_12_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_12_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_12_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_12_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_12_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_13_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_13_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_13_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_13_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_13_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_13_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_13_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_13_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_13_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_13_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_13_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_13_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_13_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_13_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_13_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_13_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_13_cse ) begin
      act_mem_banks_bank_a_13_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_13_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_13_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_13_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_13_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_13_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_13_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_13_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_13_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_13_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_13_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_13_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_13_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_13_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_13_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_13_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_14_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_14_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_14_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_14_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_14_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_14_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_14_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_14_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_14_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_14_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_14_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_14_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_14_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_14_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_14_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_14_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_14_cse ) begin
      act_mem_banks_bank_a_14_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_14_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_14_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_14_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_14_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_14_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_14_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_14_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_14_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_14_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_14_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_14_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_14_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_14_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_14_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_14_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_15_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_15_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_15_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_15_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_15_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_15_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_15_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_15_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_15_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_15_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_15_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_15_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_15_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_15_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_15_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_15_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_15_cse ) begin
      act_mem_banks_bank_a_15_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_15_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_15_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_15_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_15_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_15_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_15_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_15_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_15_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_15_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_15_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_15_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_15_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_15_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_15_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_15_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_16_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_16_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_16_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_16_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_16_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_16_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_16_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_16_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_16_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_16_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_16_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_16_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_16_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_16_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_16_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_16_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_16_cse ) begin
      act_mem_banks_bank_a_16_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_16_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_16_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_16_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_16_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_16_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_16_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_16_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_16_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_16_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_16_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_16_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_16_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_16_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_16_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_16_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_17_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_17_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_17_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_17_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_17_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_17_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_17_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_17_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_17_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_17_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_17_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_17_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_17_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_17_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_17_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_17_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_17_cse ) begin
      act_mem_banks_bank_a_17_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_17_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_17_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_17_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_17_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_17_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_17_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_17_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_17_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_17_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_17_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_17_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_17_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_17_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_17_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_17_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_18_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_18_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_18_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_18_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_18_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_18_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_18_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_18_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_18_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_18_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_18_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_18_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_18_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_18_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_18_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_18_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_18_cse ) begin
      act_mem_banks_bank_a_18_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_18_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_18_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_18_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_18_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_18_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_18_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_18_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_18_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_18_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_18_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_18_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_18_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_18_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_18_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_18_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_19_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_19_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_19_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_19_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_19_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_19_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_19_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_19_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_19_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_19_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_19_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_19_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_19_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_19_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_19_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_19_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_19_cse ) begin
      act_mem_banks_bank_a_19_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_19_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_19_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_19_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_19_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_19_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_19_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_19_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_19_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_19_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_19_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_19_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_19_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_19_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_19_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_19_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_20_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_20_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_20_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_20_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_20_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_20_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_20_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_20_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_20_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_20_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_20_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_20_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_20_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_20_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_20_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_20_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_20_cse ) begin
      act_mem_banks_bank_a_20_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_20_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_20_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_20_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_20_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_20_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_20_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_20_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_20_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_20_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_20_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_20_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_20_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_20_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_20_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_20_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_21_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_21_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_21_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_21_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_21_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_21_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_21_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_21_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_21_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_21_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_21_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_21_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_21_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_21_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_21_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_21_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_21_cse ) begin
      act_mem_banks_bank_a_21_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_21_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_21_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_21_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_21_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_21_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_21_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_21_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_21_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_21_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_21_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_21_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_21_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_21_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_21_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_21_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_22_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_22_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_22_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_22_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_22_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_22_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_22_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_22_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_22_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_22_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_22_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_22_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_22_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_22_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_22_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_22_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_22_cse ) begin
      act_mem_banks_bank_a_22_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_22_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_22_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_22_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_22_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_22_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_22_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_22_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_22_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_22_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_22_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_22_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_22_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_22_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_22_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_22_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_23_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_23_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_23_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_23_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_23_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_23_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_23_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_23_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_23_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_23_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_23_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_23_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_23_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_23_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_23_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_23_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_23_cse ) begin
      act_mem_banks_bank_a_23_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_23_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_23_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_23_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_23_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_23_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_23_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_23_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_23_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_23_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_23_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_23_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_23_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_23_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_23_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_23_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_24_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_24_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_24_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_24_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_24_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_24_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_24_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_24_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_24_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_24_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_24_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_24_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_24_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_24_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_24_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_24_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_24_cse ) begin
      act_mem_banks_bank_a_24_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_24_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_24_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_24_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_24_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_24_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_24_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_24_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_24_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_24_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_24_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_24_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_24_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_24_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_24_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_24_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_25_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_25_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_25_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_25_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_25_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_25_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_25_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_25_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_25_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_25_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_25_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_25_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_25_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_25_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_25_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_25_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_25_cse ) begin
      act_mem_banks_bank_a_25_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_25_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_25_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_25_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_25_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_25_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_25_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_25_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_25_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_25_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_25_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_25_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_25_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_25_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_25_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_25_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_26_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_26_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_26_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_26_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_26_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_26_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_26_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_26_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_26_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_26_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_26_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_26_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_26_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_26_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_26_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_26_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_26_cse ) begin
      act_mem_banks_bank_a_26_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_26_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_26_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_26_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_26_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_26_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_26_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_26_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_26_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_26_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_26_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_26_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_26_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_26_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_26_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_26_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_27_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_27_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_27_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_27_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_27_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_27_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_27_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_27_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_27_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_27_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_27_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_27_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_27_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_27_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_27_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_27_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_27_cse ) begin
      act_mem_banks_bank_a_27_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_27_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_27_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_27_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_27_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_27_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_27_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_27_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_27_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_27_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_27_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_27_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_27_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_27_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_27_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_27_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_28_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_28_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_28_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_28_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_28_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_28_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_28_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_28_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_28_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_28_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_28_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_28_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_28_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_28_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_28_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_28_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_28_cse ) begin
      act_mem_banks_bank_a_28_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_28_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_28_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_28_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_28_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_28_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_28_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_28_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_28_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_28_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_28_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_28_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_28_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_28_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_28_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_28_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_29_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_29_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_29_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_29_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_29_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_29_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_29_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_29_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_29_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_29_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_29_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_29_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_29_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_29_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_29_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_29_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_29_cse ) begin
      act_mem_banks_bank_a_29_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_29_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_29_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_29_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_29_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_29_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_29_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_29_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_29_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_29_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_29_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_29_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_29_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_29_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_29_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_29_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_30_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_30_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_30_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_30_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_30_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_30_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_30_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_30_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_30_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_30_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_30_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_30_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_30_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_30_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_30_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_30_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_30_cse ) begin
      act_mem_banks_bank_a_30_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_30_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_30_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_30_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_30_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_30_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_30_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_30_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_30_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_30_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_30_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_30_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_30_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_30_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_30_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_30_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_31_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_31_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_31_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_31_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_31_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_31_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_31_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_31_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_31_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_31_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_31_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_31_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_31_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_31_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_31_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_31_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_31_cse ) begin
      act_mem_banks_bank_a_31_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_31_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_31_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_31_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_31_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_31_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_31_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_31_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_31_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_31_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_31_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_31_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_31_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_31_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_31_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_31_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_config_inst_regs_16_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_17_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_18_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_19_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_20_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_21_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_22_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_23_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_24_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_25_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_26_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_27_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_28_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_29_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_30_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_31_sva_dfm_6 <= 8'b00000000;
    end
    else if ( act_config_inst_regs_and_4_cse ) begin
      act_config_inst_regs_16_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[7:0];
      act_config_inst_regs_17_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[15:8];
      act_config_inst_regs_18_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[23:16];
      act_config_inst_regs_19_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[31:24];
      act_config_inst_regs_20_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[39:32];
      act_config_inst_regs_21_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[47:40];
      act_config_inst_regs_22_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[55:48];
      act_config_inst_regs_23_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[63:56];
      act_config_inst_regs_24_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[71:64];
      act_config_inst_regs_25_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[79:72];
      act_config_inst_regs_26_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[87:80];
      act_config_inst_regs_27_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[95:88];
      act_config_inst_regs_28_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[103:96];
      act_config_inst_regs_29_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[111:104];
      act_config_inst_regs_30_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[119:112];
      act_config_inst_regs_31_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[127:120];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_config_inst_regs_0_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_1_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_2_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_3_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_4_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_5_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_6_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_7_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_8_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_9_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_10_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_11_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_12_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_13_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_14_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_15_sva_dfm_5 <= 8'b00000000;
    end
    else if ( act_config_inst_regs_and_20_cse ) begin
      act_config_inst_regs_0_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[7:0];
      act_config_inst_regs_1_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[15:8];
      act_config_inst_regs_2_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[23:16];
      act_config_inst_regs_3_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[31:24];
      act_config_inst_regs_4_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[39:32];
      act_config_inst_regs_5_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[47:40];
      act_config_inst_regs_6_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[55:48];
      act_config_inst_regs_7_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[63:56];
      act_config_inst_regs_8_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[71:64];
      act_config_inst_regs_9_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[79:72];
      act_config_inst_regs_10_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[87:80];
      act_config_inst_regs_11_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[95:88];
      act_config_inst_regs_12_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[103:96];
      act_config_inst_regs_13_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[111:104];
      act_config_inst_regs_14_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[119:112];
      act_config_inst_regs_15_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[127:120];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_config_output_counter_sva <= 8'b00000000;
    end
    else if ( ActUnitRun_wen & ((and_dcpl_553 & and_dcpl_789 & ActUnit_CheckStart_start_reg_sva)
        | act_config_output_counter_sva_mx0c1) ) begin
      act_config_output_counter_sva <= MUX_v_8_2_2(act_config_InstIncr_if_act_config_InstIncr_if_and_1_nl,
          act_config_output_counter_sva_dfm_3, act_config_output_counter_sva_mx0c1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_config_inst_counter_sva <= 5'b00000;
    end
    else if ( act_config_inst_counter_and_tmp ) begin
      act_config_inst_counter_sva <= MUX_v_5_2_2(act_config_InstIncr_act_config_InstIncr_and_1_nl,
          act_config_inst_counter_sva_dfm_3, act_config_inst_counter_sva_mx0c1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_15_sva_31 <= 1'b0;
      act_regs_data_3_14_sva_31 <= 1'b0;
      act_regs_data_3_13_sva_31 <= 1'b0;
      act_regs_data_3_12_sva_31 <= 1'b0;
      act_regs_data_3_11_sva_31 <= 1'b0;
      act_regs_data_3_10_sva_31 <= 1'b0;
      act_regs_data_3_9_sva_31 <= 1'b0;
      act_regs_data_3_8_sva_31 <= 1'b0;
      act_regs_data_3_7_sva_31 <= 1'b0;
      act_regs_data_3_6_sva_31 <= 1'b0;
      act_regs_data_3_5_sva_31 <= 1'b0;
      act_regs_data_3_4_sva_31 <= 1'b0;
      act_regs_data_3_3_sva_31 <= 1'b0;
      act_regs_data_3_2_sva_31 <= 1'b0;
      act_regs_data_3_1_sva_31 <= 1'b0;
      act_regs_data_3_0_sva_31 <= 1'b0;
      act_regs_data_2_15_sva_31 <= 1'b0;
      act_regs_data_2_14_sva_31 <= 1'b0;
      act_regs_data_2_13_sva_31 <= 1'b0;
      act_regs_data_2_12_sva_31 <= 1'b0;
      act_regs_data_2_11_sva_31 <= 1'b0;
      act_regs_data_2_10_sva_31 <= 1'b0;
      act_regs_data_2_9_sva_31 <= 1'b0;
      act_regs_data_2_8_sva_31 <= 1'b0;
      act_regs_data_2_7_sva_31 <= 1'b0;
      act_regs_data_2_6_sva_31 <= 1'b0;
      act_regs_data_2_5_sva_31 <= 1'b0;
      act_regs_data_2_4_sva_31 <= 1'b0;
      act_regs_data_2_3_sva_31 <= 1'b0;
      act_regs_data_2_2_sva_31 <= 1'b0;
      act_regs_data_2_1_sva_31 <= 1'b0;
      act_regs_data_2_0_sva_31 <= 1'b0;
      act_regs_data_1_15_sva_31 <= 1'b0;
      act_regs_data_1_14_sva_31 <= 1'b0;
      act_regs_data_1_13_sva_31 <= 1'b0;
      act_regs_data_1_12_sva_31 <= 1'b0;
      act_regs_data_1_11_sva_31 <= 1'b0;
      act_regs_data_1_10_sva_31 <= 1'b0;
      act_regs_data_1_9_sva_31 <= 1'b0;
      act_regs_data_1_8_sva_31 <= 1'b0;
      act_regs_data_1_7_sva_31 <= 1'b0;
      act_regs_data_1_6_sva_31 <= 1'b0;
      act_regs_data_1_5_sva_31 <= 1'b0;
      act_regs_data_1_4_sva_31 <= 1'b0;
      act_regs_data_1_3_sva_31 <= 1'b0;
      act_regs_data_1_2_sva_31 <= 1'b0;
      act_regs_data_1_1_sva_31 <= 1'b0;
      act_regs_data_1_0_sva_31 <= 1'b0;
      act_regs_data_0_15_sva_31 <= 1'b0;
      act_regs_data_0_14_sva_31 <= 1'b0;
      act_regs_data_0_13_sva_31 <= 1'b0;
      act_regs_data_0_12_sva_31 <= 1'b0;
      act_regs_data_0_11_sva_31 <= 1'b0;
      act_regs_data_0_10_sva_31 <= 1'b0;
      act_regs_data_0_9_sva_31 <= 1'b0;
      act_regs_data_0_8_sva_31 <= 1'b0;
      act_regs_data_0_7_sva_31 <= 1'b0;
      act_regs_data_0_6_sva_31 <= 1'b0;
      act_regs_data_0_5_sva_31 <= 1'b0;
      act_regs_data_0_4_sva_31 <= 1'b0;
      act_regs_data_0_3_sva_31 <= 1'b0;
      act_regs_data_0_2_sva_31 <= 1'b0;
      act_regs_data_0_1_sva_31 <= 1'b0;
      act_regs_data_0_0_sva_31 <= 1'b0;
    end
    else if ( act_regs_data_and_cse ) begin
      act_regs_data_3_15_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_3_15_sva_dfm_2_31,
          act_regs_data_2_2_sva_8_31, act_regs_data_3_15_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_3_14_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_3_14_sva_dfm_2_31,
          act_regs_data_2_15_sva_8_31, act_regs_data_3_14_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_3_13_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_3_13_sva_dfm_2_31,
          act_regs_data_2_14_sva_8_31, act_regs_data_3_13_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_3_12_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_3_12_sva_dfm_2_31,
          act_regs_data_2_13_sva_8_31, act_regs_data_3_12_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_3_11_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_3_11_sva_dfm_2_31,
          act_regs_data_2_12_sva_8_31, act_regs_data_3_11_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_3_10_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_3_10_sva_dfm_2_31,
          act_regs_data_2_11_sva_8_31, act_regs_data_3_10_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_3_9_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_3_9_sva_dfm_2_31,
          act_regs_data_3_0_sva_8_31, act_regs_data_3_9_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_3_8_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_3_8_sva_dfm_2_31,
          act_regs_data_2_9_sva_8_31, act_regs_data_3_8_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_3_7_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_3_7_sva_dfm_2_31,
          act_regs_data_2_8_sva_8_31, act_regs_data_3_7_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_3_6_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_3_6_sva_dfm_2_31,
          act_regs_data_2_7_sva_8_31, act_regs_data_3_6_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_3_5_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_3_5_sva_dfm_2_31,
          act_regs_data_2_6_sva_8_31, act_regs_data_3_5_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_3_4_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_3_4_sva_dfm_2_31,
          act_regs_data_2_5_sva_8_31, act_regs_data_3_4_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_3_3_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_3_3_sva_dfm_2_31,
          act_regs_data_2_4_sva_8_31, act_regs_data_3_3_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_3_2_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_3_2_sva_dfm_2_31,
          act_regs_data_2_3_sva_8_31, act_regs_data_3_2_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_3_1_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_3_1_sva_dfm_2_31,
          act_regs_data_2_10_sva_8_31, act_regs_data_3_1_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_3_0_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_3_0_sva_dfm_2_31,
          act_regs_data_2_1_sva_8_31, act_regs_data_3_0_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_2_15_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_2_15_sva_dfm_2_31,
          act_regs_data_1_2_sva_8_31, act_regs_data_2_15_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_2_14_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_2_14_sva_dfm_2_31,
          act_regs_data_1_15_sva_8_31, act_regs_data_2_14_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_2_13_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_2_13_sva_dfm_2_31,
          act_regs_data_1_14_sva_8_31, act_regs_data_2_13_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_2_12_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_2_12_sva_dfm_2_31,
          act_regs_data_1_13_sva_8_31, act_regs_data_2_12_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_2_11_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_2_11_sva_dfm_2_31,
          act_regs_data_1_12_sva_8_31, act_regs_data_2_11_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_2_10_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_2_10_sva_dfm_2_31,
          act_regs_data_1_11_sva_8_31, act_regs_data_2_10_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_2_9_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_2_9_sva_dfm_2_31,
          act_regs_data_2_0_sva_8_31, act_regs_data_2_9_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_2_8_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_2_8_sva_dfm_2_31,
          act_regs_data_1_9_sva_8_31, act_regs_data_2_8_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_2_7_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_2_7_sva_dfm_2_31,
          act_regs_data_1_8_sva_8_31, act_regs_data_2_7_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_2_6_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_2_6_sva_dfm_2_31,
          act_regs_data_1_7_sva_8_31, act_regs_data_2_6_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_2_5_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_2_5_sva_dfm_2_31,
          act_regs_data_1_6_sva_8_31, act_regs_data_2_5_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_2_4_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_2_4_sva_dfm_2_31,
          act_regs_data_1_5_sva_8_31, act_regs_data_2_4_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_2_3_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_2_3_sva_dfm_2_31,
          act_regs_data_1_4_sva_8_31, act_regs_data_2_3_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_2_2_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_2_2_sva_dfm_2_31,
          act_regs_data_1_3_sva_8_31, act_regs_data_2_2_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_2_1_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_2_1_sva_dfm_2_31,
          act_regs_data_1_10_sva_8_31, act_regs_data_2_1_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_2_0_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_2_0_sva_dfm_2_31,
          act_regs_data_1_1_sva_8_31, act_regs_data_2_0_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_1_15_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_1_15_sva_dfm_2_31,
          act_regs_data_0_2_sva_8_31, act_regs_data_1_15_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_1_14_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_1_14_sva_dfm_2_31,
          act_regs_data_0_15_sva_8_31, act_regs_data_1_14_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_1_13_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_1_13_sva_dfm_2_31,
          act_regs_data_0_14_sva_8_31, act_regs_data_1_13_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_1_12_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_1_12_sva_dfm_2_31,
          act_regs_data_0_13_sva_8_31, act_regs_data_1_12_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_1_11_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_1_11_sva_dfm_2_31,
          act_regs_data_0_12_sva_8_31, act_regs_data_1_11_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_1_10_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_1_10_sva_dfm_2_31,
          act_regs_data_0_11_sva_8_31, act_regs_data_1_10_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_1_9_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_1_9_sva_dfm_2_31,
          act_regs_data_1_0_sva_8_31, act_regs_data_1_9_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_1_8_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_1_8_sva_dfm_2_31,
          act_regs_data_0_9_sva_8_31, act_regs_data_1_8_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_1_7_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_1_7_sva_dfm_2_31,
          act_regs_data_0_8_sva_8_31, act_regs_data_1_7_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_1_6_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_1_6_sva_dfm_2_31,
          act_regs_data_0_7_sva_8_31, act_regs_data_1_6_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_1_5_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_1_5_sva_dfm_2_31,
          act_regs_data_0_6_sva_8_31, act_regs_data_1_5_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_1_4_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_1_4_sva_dfm_2_31,
          act_regs_data_0_5_sva_8_31, act_regs_data_1_4_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_1_3_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_1_3_sva_dfm_2_31,
          act_regs_data_0_4_sva_8_31, act_regs_data_1_3_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_1_2_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_1_2_sva_dfm_2_31,
          act_regs_data_0_3_sva_8_31, act_regs_data_1_2_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_1_1_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_1_1_sva_dfm_2_31,
          act_regs_data_0_10_sva_8_31, act_regs_data_1_1_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_1_0_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_1_0_sva_dfm_2_31,
          act_regs_data_0_1_sva_8_31, act_regs_data_1_0_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_0_15_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_0_15_sva_dfm_2_31,
          ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_31, act_regs_data_0_15_sva_8_31,
          {while_asn_1397 , while_asn_1399 , while_asn_1401});
      act_regs_data_0_14_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_0_14_sva_dfm_2_31,
          ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_31, act_regs_data_0_14_sva_8_31,
          {while_asn_1397 , while_asn_1399 , while_asn_1401});
      act_regs_data_0_13_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_0_13_sva_dfm_2_31,
          ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_31, act_regs_data_0_13_sva_8_31,
          {while_asn_1397 , while_asn_1399 , while_asn_1401});
      act_regs_data_0_12_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_0_12_sva_dfm_2_31,
          ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_31, act_regs_data_0_12_sva_8_31,
          {while_asn_1397 , while_asn_1399 , while_asn_1401});
      act_regs_data_0_11_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_0_11_sva_dfm_2_31,
          ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_31, act_regs_data_0_11_sva_8_31,
          {while_asn_1397 , while_asn_1399 , while_asn_1401});
      act_regs_data_0_10_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_0_10_sva_dfm_2_31,
          ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_31, act_regs_data_0_10_sva_8_31,
          {while_asn_1397 , while_asn_1399 , while_asn_1401});
      act_regs_data_0_9_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_0_9_sva_dfm_2_31,
          act_regs_data_0_0_sva_8_31, act_regs_data_0_9_sva_8_31, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
      act_regs_data_0_8_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_0_8_sva_dfm_2_31,
          ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_31, act_regs_data_0_8_sva_8_31,
          {while_asn_1397 , while_asn_1399 , while_asn_1401});
      act_regs_data_0_7_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_0_7_sva_dfm_2_31,
          ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_31, act_regs_data_0_7_sva_8_31,
          {while_asn_1397 , while_asn_1399 , while_asn_1401});
      act_regs_data_0_6_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_0_6_sva_dfm_2_31,
          ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_31, act_regs_data_0_6_sva_8_31,
          {while_asn_1397 , while_asn_1399 , while_asn_1401});
      act_regs_data_0_5_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_0_5_sva_dfm_2_31,
          ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_31, act_regs_data_0_5_sva_8_31,
          {while_asn_1397 , while_asn_1399 , while_asn_1401});
      act_regs_data_0_4_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_0_4_sva_dfm_2_31,
          ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_31, act_regs_data_0_4_sva_8_31,
          {while_asn_1397 , while_asn_1399 , while_asn_1401});
      act_regs_data_0_3_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_0_3_sva_dfm_2_31,
          ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_31, act_regs_data_0_3_sva_8_31,
          {while_asn_1397 , while_asn_1399 , while_asn_1401});
      act_regs_data_0_2_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_0_2_sva_dfm_2_31,
          ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_31, act_regs_data_0_2_sva_8_31,
          {while_asn_1397 , while_asn_1399 , while_asn_1401});
      act_regs_data_0_1_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_0_1_sva_dfm_2_31,
          ActUnit_PushOutput_if_output_port_reg_data_data_1_sva_31, act_regs_data_0_1_sva_8_31,
          {while_asn_1397 , while_asn_1399 , while_asn_1401});
      act_regs_data_0_0_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_0_0_sva_dfm_2_31,
          ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_31, act_regs_data_0_0_sva_8_31,
          {while_asn_1397 , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_15_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_859_enex5 ) begin
      act_regs_data_3_15_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_3_15_sva_dfm_2_30_0,
          act_regs_data_2_2_sva_8_30_0, act_regs_data_3_15_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_14_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_860_enex5 ) begin
      act_regs_data_3_14_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_3_14_sva_dfm_2_30_0,
          act_regs_data_2_15_sva_8_30_0, act_regs_data_3_14_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_13_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_861_enex5 ) begin
      act_regs_data_3_13_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_3_13_sva_dfm_2_30_0,
          act_regs_data_2_14_sva_8_30_0, act_regs_data_3_13_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_12_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_862_enex5 ) begin
      act_regs_data_3_12_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_3_12_sva_dfm_2_30_0,
          act_regs_data_2_13_sva_8_30_0, act_regs_data_3_12_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_11_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_863_enex5 ) begin
      act_regs_data_3_11_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_3_11_sva_dfm_2_30_0,
          act_regs_data_2_12_sva_8_30_0, act_regs_data_3_11_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_10_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_864_enex5 ) begin
      act_regs_data_3_10_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_3_10_sva_dfm_2_30_0,
          act_regs_data_2_11_sva_8_30_0, act_regs_data_3_10_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_9_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_865_enex5 ) begin
      act_regs_data_3_9_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_3_9_sva_dfm_2_30_0,
          act_regs_data_3_0_sva_8_30_0, act_regs_data_3_9_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_8_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_866_enex5 ) begin
      act_regs_data_3_8_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_3_8_sva_dfm_2_30_0,
          act_regs_data_2_9_sva_8_30_0, act_regs_data_3_8_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_7_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_867_enex5 ) begin
      act_regs_data_3_7_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_3_7_sva_dfm_2_30_0,
          act_regs_data_2_8_sva_8_30_0, act_regs_data_3_7_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_6_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_868_enex5 ) begin
      act_regs_data_3_6_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_3_6_sva_dfm_2_30_0,
          act_regs_data_2_7_sva_8_30_0, act_regs_data_3_6_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_5_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_869_enex5 ) begin
      act_regs_data_3_5_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_3_5_sva_dfm_2_30_0,
          act_regs_data_2_6_sva_8_30_0, act_regs_data_3_5_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_4_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_870_enex5 ) begin
      act_regs_data_3_4_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_3_4_sva_dfm_2_30_0,
          act_regs_data_2_5_sva_8_30_0, act_regs_data_3_4_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_3_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_871_enex5 ) begin
      act_regs_data_3_3_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_3_3_sva_dfm_2_30_0,
          act_regs_data_2_4_sva_8_30_0, act_regs_data_3_3_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_2_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_872_enex5 ) begin
      act_regs_data_3_2_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_3_2_sva_dfm_2_30_0,
          act_regs_data_2_3_sva_8_30_0, act_regs_data_3_2_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_1_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_873_enex5 ) begin
      act_regs_data_3_1_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_3_1_sva_dfm_2_30_0,
          act_regs_data_2_10_sva_8_30_0, act_regs_data_3_1_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_0_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_874_enex5 ) begin
      act_regs_data_3_0_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_3_0_sva_dfm_2_30_0,
          act_regs_data_2_1_sva_8_30_0, act_regs_data_3_0_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_15_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_875_enex5 ) begin
      act_regs_data_2_15_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_2_15_sva_dfm_2_30_0,
          act_regs_data_1_2_sva_8_30_0, act_regs_data_2_15_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_14_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_876_enex5 ) begin
      act_regs_data_2_14_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_2_14_sva_dfm_2_30_0,
          act_regs_data_1_15_sva_8_30_0, act_regs_data_2_14_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_13_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_877_enex5 ) begin
      act_regs_data_2_13_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_2_13_sva_dfm_2_30_0,
          act_regs_data_1_14_sva_8_30_0, act_regs_data_2_13_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_12_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_878_enex5 ) begin
      act_regs_data_2_12_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_2_12_sva_dfm_2_30_0,
          act_regs_data_1_13_sva_8_30_0, act_regs_data_2_12_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_11_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_879_enex5 ) begin
      act_regs_data_2_11_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_2_11_sva_dfm_2_30_0,
          act_regs_data_1_12_sva_8_30_0, act_regs_data_2_11_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_10_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_880_enex5 ) begin
      act_regs_data_2_10_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_2_10_sva_dfm_2_30_0,
          act_regs_data_1_11_sva_8_30_0, act_regs_data_2_10_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_9_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_881_enex5 ) begin
      act_regs_data_2_9_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_2_9_sva_dfm_2_30_0,
          act_regs_data_2_0_sva_8_30_0, act_regs_data_2_9_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_8_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_882_enex5 ) begin
      act_regs_data_2_8_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_2_8_sva_dfm_2_30_0,
          act_regs_data_1_9_sva_8_30_0, act_regs_data_2_8_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_7_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_883_enex5 ) begin
      act_regs_data_2_7_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_2_7_sva_dfm_2_30_0,
          act_regs_data_1_8_sva_8_30_0, act_regs_data_2_7_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_6_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_884_enex5 ) begin
      act_regs_data_2_6_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_2_6_sva_dfm_2_30_0,
          act_regs_data_1_7_sva_8_30_0, act_regs_data_2_6_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_5_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_885_enex5 ) begin
      act_regs_data_2_5_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_2_5_sva_dfm_2_30_0,
          act_regs_data_1_6_sva_8_30_0, act_regs_data_2_5_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_4_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_886_enex5 ) begin
      act_regs_data_2_4_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_2_4_sva_dfm_2_30_0,
          act_regs_data_1_5_sva_8_30_0, act_regs_data_2_4_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_3_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_887_enex5 ) begin
      act_regs_data_2_3_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_2_3_sva_dfm_2_30_0,
          act_regs_data_1_4_sva_8_30_0, act_regs_data_2_3_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_2_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_888_enex5 ) begin
      act_regs_data_2_2_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_2_2_sva_dfm_2_30_0,
          act_regs_data_1_3_sva_8_30_0, act_regs_data_2_2_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_1_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_889_enex5 ) begin
      act_regs_data_2_1_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_2_1_sva_dfm_2_30_0,
          act_regs_data_1_10_sva_8_30_0, act_regs_data_2_1_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_0_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_890_enex5 ) begin
      act_regs_data_2_0_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_2_0_sva_dfm_2_30_0,
          act_regs_data_1_1_sva_8_30_0, act_regs_data_2_0_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_15_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_891_enex5 ) begin
      act_regs_data_1_15_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_1_15_sva_dfm_2_30_0,
          act_regs_data_0_2_sva_8_30_0, act_regs_data_1_15_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_14_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_892_enex5 ) begin
      act_regs_data_1_14_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_1_14_sva_dfm_2_30_0,
          act_regs_data_0_15_sva_8_30_0, act_regs_data_1_14_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_13_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_893_enex5 ) begin
      act_regs_data_1_13_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_1_13_sva_dfm_2_30_0,
          act_regs_data_0_14_sva_8_30_0, act_regs_data_1_13_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_12_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_894_enex5 ) begin
      act_regs_data_1_12_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_1_12_sva_dfm_2_30_0,
          act_regs_data_0_13_sva_8_30_0, act_regs_data_1_12_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_11_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_895_enex5 ) begin
      act_regs_data_1_11_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_1_11_sva_dfm_2_30_0,
          act_regs_data_0_12_sva_8_30_0, act_regs_data_1_11_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_10_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_896_enex5 ) begin
      act_regs_data_1_10_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_1_10_sva_dfm_2_30_0,
          act_regs_data_0_11_sva_8_30_0, act_regs_data_1_10_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_9_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_897_enex5 ) begin
      act_regs_data_1_9_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_1_9_sva_dfm_2_30_0,
          act_regs_data_1_0_sva_8_30_0, act_regs_data_1_9_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_8_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_898_enex5 ) begin
      act_regs_data_1_8_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_1_8_sva_dfm_2_30_0,
          act_regs_data_0_9_sva_8_30_0, act_regs_data_1_8_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_7_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_899_enex5 ) begin
      act_regs_data_1_7_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_1_7_sva_dfm_2_30_0,
          act_regs_data_0_8_sva_8_30_0, act_regs_data_1_7_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_6_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_900_enex5 ) begin
      act_regs_data_1_6_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_1_6_sva_dfm_2_30_0,
          act_regs_data_0_7_sva_8_30_0, act_regs_data_1_6_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_5_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_901_enex5 ) begin
      act_regs_data_1_5_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_1_5_sva_dfm_2_30_0,
          act_regs_data_0_6_sva_8_30_0, act_regs_data_1_5_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_4_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_902_enex5 ) begin
      act_regs_data_1_4_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_1_4_sva_dfm_2_30_0,
          act_regs_data_0_5_sva_8_30_0, act_regs_data_1_4_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_3_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_903_enex5 ) begin
      act_regs_data_1_3_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_1_3_sva_dfm_2_30_0,
          act_regs_data_0_4_sva_8_30_0, act_regs_data_1_3_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_2_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_904_enex5 ) begin
      act_regs_data_1_2_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_1_2_sva_dfm_2_30_0,
          act_regs_data_0_3_sva_8_30_0, act_regs_data_1_2_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_1_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_905_enex5 ) begin
      act_regs_data_1_1_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_1_1_sva_dfm_2_30_0,
          act_regs_data_0_10_sva_8_30_0, act_regs_data_1_1_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_0_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_906_enex5 ) begin
      act_regs_data_1_0_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_1_0_sva_dfm_2_30_0,
          act_regs_data_0_1_sva_8_30_0, act_regs_data_1_0_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_15_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_907_enex5 ) begin
      act_regs_data_0_15_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_0_15_sva_dfm_2_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_30_0, act_regs_data_0_15_sva_8_30_0,
          {while_asn_1397 , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_14_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_908_enex5 ) begin
      act_regs_data_0_14_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_0_14_sva_dfm_2_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_30_0, act_regs_data_0_14_sva_8_30_0,
          {while_asn_1397 , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_13_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_909_enex5 ) begin
      act_regs_data_0_13_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_0_13_sva_dfm_2_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_30_0, act_regs_data_0_13_sva_8_30_0,
          {while_asn_1397 , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_12_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_910_enex5 ) begin
      act_regs_data_0_12_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_0_12_sva_dfm_2_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_30_0, act_regs_data_0_12_sva_8_30_0,
          {while_asn_1397 , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_11_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_911_enex5 ) begin
      act_regs_data_0_11_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_0_11_sva_dfm_2_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_30_0, act_regs_data_0_11_sva_8_30_0,
          {while_asn_1397 , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_10_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_912_enex5 ) begin
      act_regs_data_0_10_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_0_10_sva_dfm_2_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_30_0, act_regs_data_0_10_sva_8_30_0,
          {while_asn_1397 , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_9_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_913_enex5 ) begin
      act_regs_data_0_9_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_0_9_sva_dfm_2_30_0,
          act_regs_data_0_0_sva_8_30_0, act_regs_data_0_9_sva_8_30_0, {while_asn_1397
          , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_8_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_914_enex5 ) begin
      act_regs_data_0_8_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_0_8_sva_dfm_2_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_30_0, act_regs_data_0_8_sva_8_30_0,
          {while_asn_1397 , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_7_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_915_enex5 ) begin
      act_regs_data_0_7_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_0_7_sva_dfm_2_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_30_0, act_regs_data_0_7_sva_8_30_0,
          {while_asn_1397 , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_6_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_916_enex5 ) begin
      act_regs_data_0_6_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_0_6_sva_dfm_2_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_30_0, act_regs_data_0_6_sva_8_30_0,
          {while_asn_1397 , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_5_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_917_enex5 ) begin
      act_regs_data_0_5_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_0_5_sva_dfm_2_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_30_0, act_regs_data_0_5_sva_8_30_0,
          {while_asn_1397 , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_4_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_918_enex5 ) begin
      act_regs_data_0_4_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_0_4_sva_dfm_2_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_30_0, act_regs_data_0_4_sva_8_30_0,
          {while_asn_1397 , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_3_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_919_enex5 ) begin
      act_regs_data_0_3_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_0_3_sva_dfm_2_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_30_0, act_regs_data_0_3_sva_8_30_0,
          {while_asn_1397 , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_2_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_920_enex5 ) begin
      act_regs_data_0_2_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_0_2_sva_dfm_2_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_30_0, act_regs_data_0_2_sva_8_30_0,
          {while_asn_1397 , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_1_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_921_enex5 ) begin
      act_regs_data_0_1_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_0_1_sva_dfm_2_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_1_sva_30_0, act_regs_data_0_1_sva_8_30_0,
          {while_asn_1397 , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_0_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_922_enex5 ) begin
      act_regs_data_0_0_sva_30_0 <= MUX1HOT_v_31_3_2(act_regs_data_0_0_sva_dfm_2_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_30_0, act_regs_data_0_0_sva_8_30_0,
          {while_asn_1397 , while_asn_1399 , while_asn_1401});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_31_0 <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_read_read_data_and_16_enex5 ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_31_0 <= act_mem_banks_read_for_mux_15_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_63_32 <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_read_read_data_and_17_enex5 ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_63_32 <= act_mem_banks_read_for_mux_14_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_95_64 <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_read_read_data_and_18_enex5 ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_95_64 <= act_mem_banks_read_for_mux_13_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_127_96 <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_read_read_data_and_19_enex5 ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_127_96 <= act_mem_banks_read_for_mux_12_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_159_128 <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_read_read_data_and_20_enex5 ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_159_128 <= act_mem_banks_read_for_mux_11_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_191_160 <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_read_read_data_and_21_enex5 ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_191_160 <= act_mem_banks_read_for_mux_10_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_223_192 <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_read_read_data_and_22_enex5 ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_223_192 <= act_mem_banks_read_for_mux_9_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_255_224 <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_read_read_data_and_23_enex5 ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_255_224 <= act_mem_banks_read_for_mux_8_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_287_256 <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_read_read_data_and_24_enex5 ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_287_256 <= act_mem_banks_read_for_mux_7_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_319_288 <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_read_read_data_and_25_enex5 ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_319_288 <= act_mem_banks_read_for_mux_6_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_351_320 <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_read_read_data_and_26_enex5 ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_351_320 <= act_mem_banks_read_for_mux_5_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_383_352 <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_read_read_data_and_27_enex5 ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_383_352 <= act_mem_banks_read_for_mux_4_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_415_384 <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_read_read_data_and_28_enex5 ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_415_384 <= act_mem_banks_read_for_mux_3_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_447_416 <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_read_read_data_and_29_enex5 ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_447_416 <= act_mem_banks_read_for_mux_2_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_479_448 <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_read_read_data_and_30_enex5 ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_479_448 <= act_mem_banks_read_for_mux_1_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_511_480 <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_read_read_data_and_31_enex5 ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_511_480 <= act_mem_banks_read_for_mux_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_read_out_data_0_0_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_port_read_out_data_and_16_enex5 ) begin
      act_port_read_out_data_0_0_sva_dfm <= act_mem_banks_read_read_data_lpi_1_dfm_1_31_0_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_read_out_data_0_1_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_port_read_out_data_and_17_enex5 ) begin
      act_port_read_out_data_0_1_sva_dfm <= act_mem_banks_read_read_data_lpi_1_dfm_1_63_32_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_read_out_data_0_2_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_port_read_out_data_and_18_enex5 ) begin
      act_port_read_out_data_0_2_sva_dfm <= act_mem_banks_read_read_data_lpi_1_dfm_1_95_64_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_read_out_data_0_3_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_port_read_out_data_and_19_enex5 ) begin
      act_port_read_out_data_0_3_sva_dfm <= act_mem_banks_read_read_data_lpi_1_dfm_1_127_96_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_read_out_data_0_4_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_port_read_out_data_and_20_enex5 ) begin
      act_port_read_out_data_0_4_sva_dfm <= act_mem_banks_read_read_data_lpi_1_dfm_1_159_128_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_read_out_data_0_5_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_port_read_out_data_and_21_enex5 ) begin
      act_port_read_out_data_0_5_sva_dfm <= act_mem_banks_read_read_data_lpi_1_dfm_1_191_160_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_read_out_data_0_6_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_port_read_out_data_and_22_enex5 ) begin
      act_port_read_out_data_0_6_sva_dfm <= act_mem_banks_read_read_data_lpi_1_dfm_1_223_192_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_read_out_data_0_7_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_port_read_out_data_and_23_enex5 ) begin
      act_port_read_out_data_0_7_sva_dfm <= act_mem_banks_read_read_data_lpi_1_dfm_1_255_224_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_read_out_data_0_8_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_port_read_out_data_and_24_enex5 ) begin
      act_port_read_out_data_0_8_sva_dfm <= act_mem_banks_read_read_data_lpi_1_dfm_1_287_256_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_read_out_data_0_9_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_port_read_out_data_and_25_enex5 ) begin
      act_port_read_out_data_0_9_sva_dfm <= act_mem_banks_read_read_data_lpi_1_dfm_1_319_288_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_read_out_data_0_10_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_port_read_out_data_and_26_enex5 ) begin
      act_port_read_out_data_0_10_sva_dfm <= act_mem_banks_read_read_data_lpi_1_dfm_1_351_320_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_read_out_data_0_11_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_port_read_out_data_and_27_enex5 ) begin
      act_port_read_out_data_0_11_sva_dfm <= act_mem_banks_read_read_data_lpi_1_dfm_1_383_352_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_read_out_data_0_12_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_port_read_out_data_and_28_enex5 ) begin
      act_port_read_out_data_0_12_sva_dfm <= act_mem_banks_read_read_data_lpi_1_dfm_1_415_384_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_read_out_data_0_13_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_port_read_out_data_and_29_enex5 ) begin
      act_port_read_out_data_0_13_sva_dfm <= act_mem_banks_read_read_data_lpi_1_dfm_1_447_416_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_read_out_data_0_14_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_port_read_out_data_and_30_enex5 ) begin
      act_port_read_out_data_0_14_sva_dfm <= act_mem_banks_read_read_data_lpi_1_dfm_1_479_448_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_read_out_data_0_15_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_port_read_out_data_and_31_enex5 ) begin
      act_port_read_out_data_0_15_sva_dfm <= act_mem_banks_read_read_data_lpi_1_dfm_1_511_480_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_write_addrs_lpi_1_dfm_5 <= 5'b00000;
    end
    else if ( mux_296_nl & (fsm_output[0]) & (~ (fsm_output[3])) & (~ (fsm_output[2]))
        & (~ (fsm_output[4])) & ActUnitRun_wen ) begin
      act_write_addrs_lpi_1_dfm_5 <= MUX_v_5_2_2(act_read_addrs_sva_2_mx0w0, ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_2_mx0w2,
          and_880_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_for_and_stg_2_7_sva <= 1'b0;
      Gelu_for_and_2_cse_sva <= 1'b0;
    end
    else if ( ActUnit_PushOutput_if_for_and_28_cse ) begin
      ActUnit_PushOutput_if_for_and_stg_2_7_sva <= MUX1HOT_s_1_4_2(Tanh_for_and_1_cse_sva_mx0w0,
          ActUnit_PushOutput_if_for_and_stg_2_7_sva_1, rva_out_reg_data_0_sva_dfm_3,
          (act_mem_banks_read_read_data_lpi_1_dfm_1_31_0[0]), {and_dcpl_788 , and_dcpl_832
          , Tanh_for_or_cse , Tanh_for_and_87_cse});
      Gelu_for_and_2_cse_sva <= MUX1HOT_s_1_3_2(Tanh_for_and_2_cse_sva_mx0w0, rva_out_reg_data_8_sva_dfm_3,
          (act_mem_banks_read_read_data_lpi_1_dfm_1_31_0[8]), {and_dcpl_788 , Tanh_for_or_cse
          , Tanh_for_and_87_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_159_128_sva_dfm_3 <= 32'b00000000000000000000000000000000;
      rva_out_reg_data_191_160_sva_dfm_3 <= 32'b00000000000000000000000000000000;
      rva_out_reg_data_223_192_sva_dfm_3 <= 32'b00000000000000000000000000000000;
      rva_out_reg_data_255_224_sva_dfm_3 <= 32'b00000000000000000000000000000000;
      rva_out_reg_data_287_256_sva_dfm_3 <= 32'b00000000000000000000000000000000;
      rva_out_reg_data_319_288_sva_dfm_3 <= 32'b00000000000000000000000000000000;
      rva_out_reg_data_351_320_sva_dfm_3 <= 32'b00000000000000000000000000000000;
      rva_out_reg_data_383_352_sva_dfm_3 <= 32'b00000000000000000000000000000000;
      rva_out_reg_data_415_384_sva_dfm_3 <= 32'b00000000000000000000000000000000;
      rva_out_reg_data_447_416_sva_dfm_3 <= 32'b00000000000000000000000000000000;
      rva_out_reg_data_479_448_sva_dfm_3 <= 32'b00000000000000000000000000000000;
      rva_out_reg_data_511_480_sva_dfm_3 <= 32'b00000000000000000000000000000000;
    end
    else if ( and_1211_cse ) begin
      rva_out_reg_data_159_128_sva_dfm_3 <= MUX_v_32_2_2(ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_13_nl,
          act_mem_banks_read_read_data_lpi_1_dfm_1_159_128, and_dcpl_803);
      rva_out_reg_data_191_160_sva_dfm_3 <= MUX_v_32_2_2(ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_12_nl,
          act_mem_banks_read_read_data_lpi_1_dfm_1_191_160, and_dcpl_803);
      rva_out_reg_data_223_192_sva_dfm_3 <= MUX_v_32_2_2(ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_11_nl,
          act_mem_banks_read_read_data_lpi_1_dfm_1_223_192, and_dcpl_803);
      rva_out_reg_data_255_224_sva_dfm_3 <= MUX_v_32_2_2(ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_10_nl,
          act_mem_banks_read_read_data_lpi_1_dfm_1_255_224, and_dcpl_803);
      rva_out_reg_data_287_256_sva_dfm_3 <= MUX_v_32_2_2(ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_9_nl,
          act_mem_banks_read_read_data_lpi_1_dfm_1_287_256, and_dcpl_803);
      rva_out_reg_data_319_288_sva_dfm_3 <= MUX_v_32_2_2(ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_8_nl,
          act_mem_banks_read_read_data_lpi_1_dfm_1_319_288, and_dcpl_803);
      rva_out_reg_data_351_320_sva_dfm_3 <= MUX_v_32_2_2(ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_7_nl,
          act_mem_banks_read_read_data_lpi_1_dfm_1_351_320, and_dcpl_803);
      rva_out_reg_data_383_352_sva_dfm_3 <= MUX_v_32_2_2(ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_6_nl,
          act_mem_banks_read_read_data_lpi_1_dfm_1_383_352, and_dcpl_803);
      rva_out_reg_data_415_384_sva_dfm_3 <= MUX_v_32_2_2(ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_5_nl,
          act_mem_banks_read_read_data_lpi_1_dfm_1_415_384, and_dcpl_803);
      rva_out_reg_data_447_416_sva_dfm_3 <= MUX_v_32_2_2(ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_4_nl,
          act_mem_banks_read_read_data_lpi_1_dfm_1_447_416, and_dcpl_803);
      rva_out_reg_data_479_448_sva_dfm_3 <= MUX_v_32_2_2(ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_3_nl,
          act_mem_banks_read_read_data_lpi_1_dfm_1_479_448, and_dcpl_803);
      rva_out_reg_data_511_480_sva_dfm_3 <= MUX_v_32_2_2(ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_nl,
          act_mem_banks_read_read_data_lpi_1_dfm_1_511_480, and_dcpl_803);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_103_96_sva_dfm_3 <= 8'b00000000;
      rva_out_reg_data_111_104_sva_dfm_3 <= 8'b00000000;
      rva_out_reg_data_119_112_sva_dfm_3 <= 8'b00000000;
      rva_out_reg_data_127_120_sva_dfm_3 <= 8'b00000000;
      rva_out_reg_data_23_16_sva_dfm_3 <= 8'b00000000;
      rva_out_reg_data_47_40_sva_dfm_3 <= 8'b00000000;
      rva_out_reg_data_63_56_sva_dfm_3 <= 8'b00000000;
      rva_out_reg_data_79_72_sva_dfm_3 <= 8'b00000000;
      rva_out_reg_data_87_80_sva_dfm_3 <= 8'b00000000;
      rva_out_reg_data_95_88_sva_dfm_3 <= 8'b00000000;
      rva_out_reg_data_31_30_sva_dfm_3 <= 2'b00;
      rva_out_reg_data_15_9_sva_dfm_3 <= 7'b0000000;
      rva_out_reg_data_7_1_sva_dfm_3 <= 7'b0000000;
      rva_out_reg_data_55_53_sva_dfm_3 <= 3'b000;
    end
    else if ( rva_out_reg_data_and_16_cse ) begin
      rva_out_reg_data_103_96_sva_dfm_3 <= MUX_v_8_2_2(and_1111_nl, (act_mem_banks_read_read_data_lpi_1_dfm_1_127_96[7:0]),
          and_dcpl_803);
      rva_out_reg_data_111_104_sva_dfm_3 <= MUX_v_8_2_2(and_1113_nl, (act_mem_banks_read_read_data_lpi_1_dfm_1_127_96[15:8]),
          and_dcpl_803);
      rva_out_reg_data_119_112_sva_dfm_3 <= MUX_v_8_2_2(and_1115_nl, (act_mem_banks_read_read_data_lpi_1_dfm_1_127_96[23:16]),
          and_dcpl_803);
      rva_out_reg_data_127_120_sva_dfm_3 <= MUX_v_8_2_2(and_1117_nl, (act_mem_banks_read_read_data_lpi_1_dfm_1_127_96[31:24]),
          and_dcpl_803);
      rva_out_reg_data_23_16_sva_dfm_3 <= MUX_v_8_2_2(and_1119_nl, (act_mem_banks_read_read_data_lpi_1_dfm_1_31_0[23:16]),
          and_dcpl_803);
      rva_out_reg_data_47_40_sva_dfm_3 <= MUX_v_8_2_2(and_1121_nl, (act_mem_banks_read_read_data_lpi_1_dfm_1_63_32[15:8]),
          and_dcpl_803);
      rva_out_reg_data_63_56_sva_dfm_3 <= MUX_v_8_2_2(and_1123_nl, (act_mem_banks_read_read_data_lpi_1_dfm_1_63_32[31:24]),
          and_dcpl_803);
      rva_out_reg_data_79_72_sva_dfm_3 <= MUX_v_8_2_2(and_1125_nl, (act_mem_banks_read_read_data_lpi_1_dfm_1_95_64[15:8]),
          and_dcpl_803);
      rva_out_reg_data_87_80_sva_dfm_3 <= MUX_v_8_2_2(and_1127_nl, (act_mem_banks_read_read_data_lpi_1_dfm_1_95_64[23:16]),
          and_dcpl_803);
      rva_out_reg_data_95_88_sva_dfm_3 <= MUX_v_8_2_2(and_1129_nl, (act_mem_banks_read_read_data_lpi_1_dfm_1_95_64[31:24]),
          and_dcpl_803);
      rva_out_reg_data_31_30_sva_dfm_3 <= MUX_v_2_2_2(and_1131_nl, (act_mem_banks_read_read_data_lpi_1_dfm_1_31_0[31:30]),
          and_dcpl_803);
      rva_out_reg_data_15_9_sva_dfm_3 <= MUX_v_7_2_2(and_1133_nl, (act_mem_banks_read_read_data_lpi_1_dfm_1_31_0[15:9]),
          and_dcpl_803);
      rva_out_reg_data_7_1_sva_dfm_3 <= MUX_v_7_2_2(and_1135_nl, (act_mem_banks_read_read_data_lpi_1_dfm_1_31_0[7:1]),
          and_dcpl_803);
      rva_out_reg_data_55_53_sva_dfm_3 <= MUX_v_3_2_2(and_1137_nl, (act_mem_banks_read_read_data_lpi_1_dfm_1_63_32[23:21]),
          and_dcpl_803);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      w_load_lpi_1_dfm_1 <= 1'b0;
    end
    else if ( w_load_and_tmp ) begin
      w_load_lpi_1_dfm_1 <= ~(ActUnit_RunInst_switch_lp_mux_1_nl | ActUnit_RunInst_switch_lp_mux_2_nl
          | ActUnit_RunInst_switch_lp_mux_4_nl | ActUnit_RunInst_switch_lp_mux_5_nl
          | ActUnit_RunInst_switch_lp_mux_7_nl | ActUnit_RunInst_switch_lp_mux_9_nl
          | ActUnit_RunInst_switch_lp_mux_11_nl | ActUnit_RunInst_switch_lp_mux_13_nl
          | ActUnit_RunInst_switch_lp_nor_tmp_mx0);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_RunInst_switch_lp_equal_tmp_2 <= 1'b0;
      ActUnit_RunInst_switch_lp_equal_tmp_4 <= 1'b0;
      ActUnit_RunInst_switch_lp_equal_tmp_5 <= 1'b0;
      ActUnit_RunInst_switch_lp_equal_tmp_6 <= 1'b0;
      ActUnit_RunInst_switch_lp_equal_tmp_7 <= 1'b0;
      ActUnit_RunInst_switch_lp_equal_tmp_8 <= 1'b0;
      Tanh_for_1_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= 1'b0;
      Tanh_for_2_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= 1'b0;
      Tanh_for_3_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= 1'b0;
      Tanh_for_4_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= 1'b0;
      Tanh_for_5_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= 1'b0;
      Tanh_for_6_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= 1'b0;
      Tanh_for_7_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= 1'b0;
      Tanh_for_8_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= 1'b0;
      Tanh_for_9_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= 1'b0;
      Tanh_for_12_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= 1'b0;
      Tanh_for_13_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= 1'b0;
      Tanh_for_14_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= 1'b0;
      Tanh_for_15_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= 1'b0;
      Tanh_for_15_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
          <= 1'b0;
      Tanh_for_14_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
          <= 1'b0;
      Tanh_for_13_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
          <= 1'b0;
      Tanh_for_12_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
          <= 1'b0;
      Tanh_for_9_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
          <= 1'b0;
      Tanh_for_8_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
          <= 1'b0;
      Tanh_for_7_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
          <= 1'b0;
      Tanh_for_6_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
          <= 1'b0;
      Tanh_for_5_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
          <= 1'b0;
      Tanh_for_4_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
          <= 1'b0;
      Tanh_for_3_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
          <= 1'b0;
      Tanh_for_2_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
          <= 1'b0;
      Tanh_for_1_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
          <= 1'b0;
    end
    else if ( ActUnit_RunInst_switch_lp_and_802_cse ) begin
      ActUnit_RunInst_switch_lp_equal_tmp_2 <= ActUnit_RunInst_switch_lp_equal_tmp_2_mx0w0;
      ActUnit_RunInst_switch_lp_equal_tmp_4 <= ActUnit_RunInst_switch_lp_equal_tmp_4_mx0w0;
      ActUnit_RunInst_switch_lp_equal_tmp_5 <= ActUnit_RunInst_switch_lp_equal_tmp_5_mx0w0;
      ActUnit_RunInst_switch_lp_equal_tmp_6 <= ActUnit_RunInst_switch_lp_equal_tmp_6_mx0w0;
      ActUnit_RunInst_switch_lp_equal_tmp_7 <= ActUnit_RunInst_switch_lp_equal_tmp_7_mx0w0;
      ActUnit_RunInst_switch_lp_equal_tmp_8 <= ActUnit_RunInst_switch_lp_equal_tmp_8_mx0w0;
      Tanh_for_1_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_15_tmp_1;
      Tanh_for_2_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_14_tmp_1;
      Tanh_for_3_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_13_tmp_1;
      Tanh_for_4_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_12_tmp_1;
      Tanh_for_5_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_11_tmp_1;
      Tanh_for_6_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_10_tmp_1;
      Tanh_for_7_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_9_tmp_1;
      Tanh_for_8_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_8_tmp_1;
      Tanh_for_9_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_7_tmp_1;
      Tanh_for_12_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_4_tmp_1;
      Tanh_for_13_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_3_tmp_1;
      Tanh_for_14_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_2_tmp_1;
      Tanh_for_15_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_1_tmp_1;
      Tanh_for_15_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_3_less_1_tmp;
      Tanh_for_14_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_3_less_2_tmp;
      Tanh_for_13_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_3_less_3_tmp;
      Tanh_for_12_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_3_less_4_tmp;
      Tanh_for_9_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_3_less_7_tmp;
      Tanh_for_8_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_3_less_8_tmp;
      Tanh_for_7_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_3_less_9_tmp;
      Tanh_for_6_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_3_less_10_tmp;
      Tanh_for_5_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_3_less_11_tmp;
      Tanh_for_4_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_3_less_12_tmp;
      Tanh_for_3_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_3_less_13_tmp;
      Tanh_for_2_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_3_less_14_tmp;
      Tanh_for_1_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_3_less_15_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= 1'b0;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= MUX_s_1_4_2(act_regs_data_0_15_sva_31, act_regs_data_1_15_sva_31, act_regs_data_2_15_sva_31,
          act_regs_data_3_15_sva_31, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= MUX_s_1_4_2(act_regs_data_0_14_sva_31, act_regs_data_1_14_sva_31, act_regs_data_2_14_sva_31,
          act_regs_data_3_14_sva_31, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= MUX_s_1_4_2(act_regs_data_0_13_sva_31, act_regs_data_1_13_sva_31, act_regs_data_2_13_sva_31,
          act_regs_data_3_13_sva_31, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= MUX_s_1_4_2(act_regs_data_0_12_sva_31, act_regs_data_1_12_sva_31, act_regs_data_2_12_sva_31,
          act_regs_data_3_12_sva_31, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= MUX_s_1_4_2(act_regs_data_0_11_sva_31, act_regs_data_1_11_sva_31, act_regs_data_2_11_sva_31,
          act_regs_data_3_11_sva_31, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= MUX_s_1_4_2(act_regs_data_0_10_sva_31, act_regs_data_1_10_sva_31, act_regs_data_2_10_sva_31,
          act_regs_data_3_10_sva_31, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= MUX_s_1_4_2(act_regs_data_0_9_sva_31, act_regs_data_1_9_sva_31, act_regs_data_2_9_sva_31,
          act_regs_data_3_9_sva_31, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= MUX_s_1_4_2(act_regs_data_0_8_sva_31, act_regs_data_1_8_sva_31, act_regs_data_2_8_sva_31,
          act_regs_data_3_8_sva_31, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= MUX_s_1_4_2(act_regs_data_0_7_sva_31, act_regs_data_1_7_sva_31, act_regs_data_2_7_sva_31,
          act_regs_data_3_7_sva_31, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= MUX_s_1_4_2(act_regs_data_0_6_sva_31, act_regs_data_1_6_sva_31, act_regs_data_2_6_sva_31,
          act_regs_data_3_6_sva_31, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= MUX_s_1_4_2(act_regs_data_0_5_sva_31, act_regs_data_1_5_sva_31, act_regs_data_2_5_sva_31,
          act_regs_data_3_5_sva_31, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= MUX_s_1_4_2(act_regs_data_0_4_sva_31, act_regs_data_1_4_sva_31, act_regs_data_2_4_sva_31,
          act_regs_data_3_4_sva_31, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= MUX_s_1_4_2(act_regs_data_0_3_sva_31, act_regs_data_1_3_sva_31, act_regs_data_2_3_sva_31,
          act_regs_data_3_3_sva_31, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= MUX_s_1_4_2(act_regs_data_0_2_sva_31, act_regs_data_1_2_sva_31, act_regs_data_2_2_sva_31,
          act_regs_data_3_2_sva_31, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= MUX_s_1_4_2(act_regs_data_0_1_sva_31, act_regs_data_1_1_sva_31, act_regs_data_2_1_sva_31,
          act_regs_data_3_1_sva_31, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= MUX_s_1_4_2(act_regs_data_0_0_sva_31, act_regs_data_1_0_sva_31, act_regs_data_2_0_sva_31,
          act_regs_data_3_0_sva_31, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_37_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0
          <= MUX_v_31_4_2(act_regs_data_0_15_sva_30_0, act_regs_data_1_15_sva_30_0,
          act_regs_data_2_15_sva_30_0, act_regs_data_3_15_sva_30_0, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_38_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0
          <= MUX_v_31_4_2(act_regs_data_0_14_sva_30_0, act_regs_data_1_14_sva_30_0,
          act_regs_data_2_14_sva_30_0, act_regs_data_3_14_sva_30_0, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_39_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0
          <= MUX_v_31_4_2(act_regs_data_0_13_sva_30_0, act_regs_data_1_13_sva_30_0,
          act_regs_data_2_13_sva_30_0, act_regs_data_3_13_sva_30_0, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_40_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0
          <= MUX_v_31_4_2(act_regs_data_0_12_sva_30_0, act_regs_data_1_12_sva_30_0,
          act_regs_data_2_12_sva_30_0, act_regs_data_3_12_sva_30_0, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_41_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0
          <= MUX_v_31_4_2(act_regs_data_0_11_sva_30_0, act_regs_data_1_11_sva_30_0,
          act_regs_data_2_11_sva_30_0, act_regs_data_3_11_sva_30_0, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_42_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0
          <= MUX_v_31_4_2(act_regs_data_0_10_sva_30_0, act_regs_data_1_10_sva_30_0,
          act_regs_data_2_10_sva_30_0, act_regs_data_3_10_sva_30_0, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_43_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0
          <= MUX_v_31_4_2(act_regs_data_0_9_sva_30_0, act_regs_data_1_9_sva_30_0,
          act_regs_data_2_9_sva_30_0, act_regs_data_3_9_sva_30_0, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_44_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0
          <= MUX_v_31_4_2(act_regs_data_0_8_sva_30_0, act_regs_data_1_8_sva_30_0,
          act_regs_data_2_8_sva_30_0, act_regs_data_3_8_sva_30_0, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_45_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0
          <= MUX_v_31_4_2(act_regs_data_0_7_sva_30_0, act_regs_data_1_7_sva_30_0,
          act_regs_data_2_7_sva_30_0, act_regs_data_3_7_sva_30_0, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_46_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0
          <= MUX_v_31_4_2(act_regs_data_0_6_sva_30_0, act_regs_data_1_6_sva_30_0,
          act_regs_data_2_6_sva_30_0, act_regs_data_3_6_sva_30_0, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_47_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0
          <= MUX_v_31_4_2(act_regs_data_0_5_sva_30_0, act_regs_data_1_5_sva_30_0,
          act_regs_data_2_5_sva_30_0, act_regs_data_3_5_sva_30_0, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_48_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0
          <= MUX_v_31_4_2(act_regs_data_0_4_sva_30_0, act_regs_data_1_4_sva_30_0,
          act_regs_data_2_4_sva_30_0, act_regs_data_3_4_sva_30_0, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_49_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0
          <= MUX_v_31_4_2(act_regs_data_0_3_sva_30_0, act_regs_data_1_3_sva_30_0,
          act_regs_data_2_3_sva_30_0, act_regs_data_3_3_sva_30_0, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_50_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0
          <= MUX_v_31_4_2(act_regs_data_0_2_sva_30_0, act_regs_data_1_2_sva_30_0,
          act_regs_data_2_2_sva_30_0, act_regs_data_3_2_sva_30_0, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_51_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0
          <= MUX_v_31_4_2(act_regs_data_0_1_sva_30_0, act_regs_data_1_1_sva_30_0,
          act_regs_data_2_1_sva_30_0, act_regs_data_3_1_sva_30_0, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_52_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0
          <= MUX_v_31_4_2(act_regs_data_0_0_sva_30_0, act_regs_data_1_0_sva_30_0,
          act_regs_data_2_0_sva_30_0, act_regs_data_3_0_sva_30_0, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Tanh_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= 1'b0;
    end
    else if ( ActUnit_RunInst_switch_lp_and_802_cse & and_dcpl_13 & (~((act_config_in_InstFetch_mux_tmp[6])
        & operator_32_8_true_AC_TRN_AC_WRAP_3_less_6_tmp)) & (act_config_in_InstFetch_mux_tmp[7])
        ) begin
      Tanh_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_6_tmp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Tanh_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= 1'b0;
    end
    else if ( ActUnit_RunInst_switch_lp_and_802_cse & and_dcpl_13 & (~((act_config_in_InstFetch_mux_tmp[6])
        & operator_32_8_true_AC_TRN_AC_WRAP_3_less_5_tmp)) & (act_config_in_InstFetch_mux_tmp[7])
        ) begin
      Tanh_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_5_tmp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Tanh_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= 1'b0;
    end
    else if ( ActUnit_RunInst_switch_lp_and_802_cse & and_dcpl_13 & (~((act_config_in_InstFetch_mux_tmp[6])
        & operator_32_8_true_AC_TRN_AC_WRAP_3_less_tmp)) & (act_config_in_InstFetch_mux_tmp[7])
        ) begin
      Tanh_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_tmp_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_lpi_1_dfm <= 31'b0000000000000000000000000000000;
    end
    else if ( Relu_for_y_qelse_and_31_enex5 ) begin
      Relu_for_y_qr_30_0_lpi_1_dfm <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0,
          nv_scvector_cctor_nv_scvector_4_for_not_14_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_15_lpi_1_dfm <= 31'b0000000000000000000000000000000;
    end
    else if ( Relu_for_y_qelse_and_32_enex5 ) begin
      Relu_for_y_qr_30_0_15_lpi_1_dfm <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0,
          nv_scvector_cctor_nv_scvector_4_for_not_13_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_14_lpi_1_dfm <= 31'b0000000000000000000000000000000;
    end
    else if ( Relu_for_y_qelse_and_33_enex5 ) begin
      Relu_for_y_qr_30_0_14_lpi_1_dfm <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0,
          nv_scvector_cctor_nv_scvector_4_for_not_12_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_13_lpi_1_dfm <= 31'b0000000000000000000000000000000;
    end
    else if ( Relu_for_y_qelse_and_34_enex5 ) begin
      Relu_for_y_qr_30_0_13_lpi_1_dfm <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0,
          nv_scvector_cctor_nv_scvector_4_for_not_11_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_12_lpi_1_dfm <= 31'b0000000000000000000000000000000;
    end
    else if ( Relu_for_y_qelse_and_35_enex5 ) begin
      Relu_for_y_qr_30_0_12_lpi_1_dfm <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0,
          nv_scvector_cctor_nv_scvector_4_for_not_10_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_11_lpi_1_dfm <= 31'b0000000000000000000000000000000;
    end
    else if ( Relu_for_y_qelse_and_36_enex5 ) begin
      Relu_for_y_qr_30_0_11_lpi_1_dfm <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0,
          nv_scvector_cctor_nv_scvector_4_for_not_9_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_10_lpi_1_dfm <= 31'b0000000000000000000000000000000;
    end
    else if ( Relu_for_y_qelse_and_37_enex5 ) begin
      Relu_for_y_qr_30_0_10_lpi_1_dfm <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0,
          nv_scvector_cctor_nv_scvector_4_for_not_8_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_9_lpi_1_dfm <= 31'b0000000000000000000000000000000;
    end
    else if ( Relu_for_y_qelse_and_38_enex5 ) begin
      Relu_for_y_qr_30_0_9_lpi_1_dfm <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0,
          nv_scvector_cctor_nv_scvector_4_for_not_7_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_8_lpi_1_dfm <= 31'b0000000000000000000000000000000;
    end
    else if ( Relu_for_y_qelse_and_39_enex5 ) begin
      Relu_for_y_qr_30_0_8_lpi_1_dfm <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0,
          nv_scvector_cctor_nv_scvector_4_for_not_6_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_7_lpi_1_dfm <= 31'b0000000000000000000000000000000;
    end
    else if ( Relu_for_y_qelse_and_40_enex5 ) begin
      Relu_for_y_qr_30_0_7_lpi_1_dfm <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0,
          nv_scvector_cctor_nv_scvector_4_for_not_5_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_6_lpi_1_dfm <= 31'b0000000000000000000000000000000;
    end
    else if ( Relu_for_y_qelse_and_41_enex5 ) begin
      Relu_for_y_qr_30_0_6_lpi_1_dfm <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0,
          nv_scvector_cctor_nv_scvector_4_for_not_4_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_5_lpi_1_dfm <= 31'b0000000000000000000000000000000;
    end
    else if ( Relu_for_y_qelse_and_42_enex5 ) begin
      Relu_for_y_qr_30_0_5_lpi_1_dfm <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0,
          nv_scvector_cctor_nv_scvector_4_for_not_3_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_4_lpi_1_dfm <= 31'b0000000000000000000000000000000;
    end
    else if ( Relu_for_y_qelse_and_43_enex5 ) begin
      Relu_for_y_qr_30_0_4_lpi_1_dfm <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0,
          nv_scvector_cctor_nv_scvector_4_for_not_2_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_3_lpi_1_dfm <= 31'b0000000000000000000000000000000;
    end
    else if ( Relu_for_y_qelse_and_44_enex5 ) begin
      Relu_for_y_qr_30_0_3_lpi_1_dfm <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0,
          nv_scvector_cctor_nv_scvector_4_for_not_1_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_2_lpi_1_dfm <= 31'b0000000000000000000000000000000;
    end
    else if ( Relu_for_y_qelse_and_45_enex5 ) begin
      Relu_for_y_qr_30_0_2_lpi_1_dfm <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0,
          nv_scvector_cctor_nv_scvector_4_for_not_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_1_lpi_1_dfm <= 31'b0000000000000000000000000000000;
    end
    else if ( Relu_for_y_qelse_and_46_enex5 ) begin
      Relu_for_y_qr_30_0_1_lpi_1_dfm <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          ActUnit_RunInst_case_11_nv_scvector_cctor_data_0_sva_1_30_0, ActUnit_RunInst_switch_lp_not_1_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_15_enex5 ) begin
      nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_16_enex5 ) begin
      nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_RunInst_case_14_nv_scvector_cctor_data_0_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( ActUnit_RunInst_switch_lp_and_815_enex5 ) begin
      ActUnit_RunInst_case_14_nv_scvector_cctor_data_0_sva_30_0 <= ActUnit_RunInst_case_11_nv_scvector_cctor_data_0_sva_1_30_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_5_for_2_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_17_enex5 ) begin
      nv_scvector_cctor_nv_scvector_5_for_2_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_18_enex5 ) begin
      nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_19_enex5 ) begin
      nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_20_enex5 ) begin
      nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_21_enex5 ) begin
      nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_22_enex5 ) begin
      nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_23_enex5 ) begin
      nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_24_enex5 ) begin
      nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_25_enex5 ) begin
      nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_26_enex5 ) begin
      nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_27_enex5 ) begin
      nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_28_enex5 ) begin
      nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_29_enex5 ) begin
      nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_6_for_3_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_enex5 ) begin
      nv_scvector_cctor_nv_scvector_6_for_3_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_6_for_12_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_15_enex5 ) begin
      nv_scvector_cctor_nv_scvector_6_for_12_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_RunInst_case_15_nv_scvector_cctor_data_0_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( ActUnit_RunInst_switch_lp_and_816_enex5 ) begin
      ActUnit_RunInst_case_15_nv_scvector_cctor_data_0_sva_30_0 <= ActUnit_RunInst_case_11_nv_scvector_cctor_data_0_sva_1_30_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_6_for_2_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_16_enex5 ) begin
      nv_scvector_cctor_nv_scvector_6_for_2_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_6_for_4_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_17_enex5 ) begin
      nv_scvector_cctor_nv_scvector_6_for_4_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_6_for_5_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_18_enex5 ) begin
      nv_scvector_cctor_nv_scvector_6_for_5_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_6_for_6_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_19_enex5 ) begin
      nv_scvector_cctor_nv_scvector_6_for_6_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_6_for_7_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_20_enex5 ) begin
      nv_scvector_cctor_nv_scvector_6_for_7_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_6_for_8_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_21_enex5 ) begin
      nv_scvector_cctor_nv_scvector_6_for_8_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_6_for_9_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_22_enex5 ) begin
      nv_scvector_cctor_nv_scvector_6_for_9_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_6_for_10_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_23_enex5 ) begin
      nv_scvector_cctor_nv_scvector_6_for_10_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_6_for_11_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_24_enex5 ) begin
      nv_scvector_cctor_nv_scvector_6_for_11_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_6_for_13_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_25_enex5 ) begin
      nv_scvector_cctor_nv_scvector_6_for_13_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_6_for_14_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_26_enex5 ) begin
      nv_scvector_cctor_nv_scvector_6_for_14_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_6_for_15_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_27_enex5 ) begin
      nv_scvector_cctor_nv_scvector_6_for_15_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_6_for_16_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= 31'b0000000000000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_28_enex5 ) begin
      nv_scvector_cctor_nv_scvector_6_for_16_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0
          <= nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_config_in_InstFetch_return_sva_7_2 <= 6'b000000;
    end
    else if ( ActUnit_RunInst_curr_inst_and_enex5 ) begin
      act_config_in_InstFetch_return_sva_7_2 <= act_config_in_InstFetch_mux_tmp[7:2];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Tanh_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
          <= 1'b0;
      Tanh_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
          <= 1'b0;
      Tanh_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
          <= 1'b0;
    end
    else if ( operator_32_8_true_AC_TRN_AC_WRAP_and_cse ) begin
      Tanh_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_3_less_tmp;
      Tanh_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_3_less_5_tmp;
      Tanh_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_3_less_6_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= 1'b0;
    end
    else if ( ActUnit_RunInst_switch_lp_and_812_cse & and_dcpl_51 & and_dcpl_47 &
        (~ operator_32_8_true_AC_TRN_AC_WRAP_2_less_15_tmp) ) begin
      Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_1_less_15_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= 1'b0;
    end
    else if ( ActUnit_RunInst_switch_lp_and_812_cse & and_dcpl_51 & and_dcpl_47 &
        (~ operator_32_8_true_AC_TRN_AC_WRAP_2_less_14_tmp) ) begin
      Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_1_less_14_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= 1'b0;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_cse & and_dcpl_51 & and_dcpl_47
        & (~ operator_32_8_true_AC_TRN_AC_WRAP_2_less_13_tmp) ) begin
      Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= $signed({1'b0, 26'b10000000000000000000000000}) < $signed(({nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
          , nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0}));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= 1'b0;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_cse & and_dcpl_51 & and_dcpl_47
        & (~ operator_32_8_true_AC_TRN_AC_WRAP_2_less_12_tmp) ) begin
      Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= $signed({1'b0, 26'b10000000000000000000000000}) < $signed(({nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
          , nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0}));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
          <= 1'b0;
      Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
          <= 1'b0;
    end
    else if ( operator_32_8_true_AC_TRN_AC_WRAP_2_and_cse ) begin
      Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_12_tmp;
      Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_13_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
          <= 1'b0;
      Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
          <= 1'b0;
    end
    else if ( operator_32_8_true_AC_TRN_AC_WRAP_2_and_17_cse ) begin
      Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_14_tmp;
      Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_15_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= 1'b0;
      Gelu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= 1'b0;
      Gelu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
          <= 1'b0;
      Gelu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
          <= 1'b0;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_7_cse ) begin
      Gelu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_15_tmp_1;
      Gelu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_14_tmp_1;
      Gelu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_3_less_14_tmp;
      Gelu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_3_less_15_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= 1'b0;
      Gelu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
          <= 1'b0;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_9_cse ) begin
      Gelu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_13_tmp_1;
      Gelu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_3_less_13_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= 1'b0;
      Gelu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
          <= 1'b0;
      Gelu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= 1'b0;
      Gelu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= 1'b0;
      Gelu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
          <= 1'b0;
      Gelu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
          <= 1'b0;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_13_cse ) begin
      Gelu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_4_tmp_1;
      Gelu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_3_less_4_tmp;
      Gelu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_10_tmp_1;
      Gelu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_9_tmp_1;
      Gelu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_3_less_9_tmp;
      Gelu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_3_less_10_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= 1'b0;
      Gelu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= 1'b0;
      Gelu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= 1'b0;
      Gelu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
          <= 1'b0;
      Gelu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
          <= 1'b0;
      Gelu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
          <= 1'b0;
      Gelu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= 1'b0;
      Gelu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= 1'b0;
      Gelu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
          <= 1'b0;
      Gelu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
          <= 1'b0;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_7_cse ) begin
      Gelu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_3_tmp_1;
      Gelu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_2_tmp_1;
      Gelu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_1_tmp_1;
      Gelu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_3_less_1_tmp;
      Gelu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_3_less_2_tmp;
      Gelu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_3_less_3_tmp;
      Gelu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_8_tmp_1;
      Gelu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_7_tmp_1;
      Gelu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_3_less_7_tmp;
      Gelu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_3_less_8_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= 1'b0;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_3_cse & and_dcpl_51 & and_dcpl_47
        & (~ operator_32_8_true_AC_TRN_AC_WRAP_2_less_11_tmp) ) begin
      Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= $signed({1'b0, 26'b10000000000000000000000000}) < $signed(({nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
          , nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0}));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= 1'b0;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_3_cse & and_dcpl_51 & and_dcpl_47
        & (~ operator_32_8_true_AC_TRN_AC_WRAP_2_less_10_tmp) ) begin
      Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= $signed({1'b0, 26'b10000000000000000000000000}) < $signed(({nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
          , nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0}));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
          <= 1'b0;
      Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
          <= 1'b0;
    end
    else if ( operator_32_8_true_AC_TRN_AC_WRAP_2_and_19_cse ) begin
      Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_10_tmp;
      Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_11_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= 1'b0;
      Gelu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= 1'b0;
      Gelu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
          <= 1'b0;
      Gelu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
          <= 1'b0;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_11_cse ) begin
      Gelu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_12_tmp_1;
      Gelu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_11_tmp_1;
      Gelu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_3_less_11_tmp;
      Gelu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_3_less_12_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= 1'b0;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_5_cse & and_dcpl_51 & and_dcpl_47
        & (~ operator_32_8_true_AC_TRN_AC_WRAP_2_less_9_tmp) ) begin
      Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= $signed({1'b0, 26'b10000000000000000000000000}) < $signed(({nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
          , nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0}));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= 1'b0;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_5_cse & and_dcpl_51 & (act_config_in_InstFetch_mux_tmp[6])
        & (~ operator_32_8_true_AC_TRN_AC_WRAP_2_less_8_tmp) & (~ (act_config_in_InstFetch_mux_tmp[4]))
        ) begin
      Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= $signed({1'b0, 26'b10000000000000000000000000}) < $signed(({nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
          , nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0}));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
          <= 1'b0;
      Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
          <= 1'b0;
    end
    else if ( operator_32_8_true_AC_TRN_AC_WRAP_2_and_21_cse ) begin
      Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_8_tmp;
      Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_9_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= 1'b0;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_7_cse & and_dcpl_51 & and_dcpl_47
        & (~ operator_32_8_true_AC_TRN_AC_WRAP_2_less_7_tmp) ) begin
      Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= $signed({1'b0, 26'b10000000000000000000000000}) < $signed(({nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
          , nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0}));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= 1'b0;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_7_cse & and_dcpl_51 & and_dcpl_47
        & (~ operator_32_8_true_AC_TRN_AC_WRAP_2_less_6_tmp) ) begin
      Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= $signed({1'b0, 26'b10000000000000000000000000}) < $signed(({nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
          , nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0}));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
          <= 1'b0;
      Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
          <= 1'b0;
    end
    else if ( operator_32_8_true_AC_TRN_AC_WRAP_2_and_23_cse ) begin
      Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_6_tmp;
      Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_7_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= 1'b0;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_9_cse & and_dcpl_51 & and_dcpl_47
        & (~ operator_32_8_true_AC_TRN_AC_WRAP_2_less_5_tmp) ) begin
      Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= $signed({1'b0, 26'b10000000000000000000000000}) < $signed(({nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
          , nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0}));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= 1'b0;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_9_cse & and_dcpl_51 & and_dcpl_47
        & (~ operator_32_8_true_AC_TRN_AC_WRAP_2_less_4_tmp) ) begin
      Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= $signed({1'b0, 26'b10000000000000000000000000}) < $signed(({nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
          , nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0}));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
          <= 1'b0;
      Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
          <= 1'b0;
    end
    else if ( operator_32_8_true_AC_TRN_AC_WRAP_2_and_25_cse ) begin
      Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_4_tmp;
      Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_5_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= 1'b0;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_11_cse & and_dcpl_51 & and_dcpl_47
        & (~ operator_32_8_true_AC_TRN_AC_WRAP_2_less_3_tmp) ) begin
      Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= $signed({1'b0, 26'b10000000000000000000000000}) < $signed(({nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
          , nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0}));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= 1'b0;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_11_cse & and_dcpl_51 & and_dcpl_47
        & (~ operator_32_8_true_AC_TRN_AC_WRAP_2_less_2_tmp) ) begin
      Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= $signed({1'b0, 26'b10000000000000000000000000}) < $signed(({nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
          , nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0}));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
          <= 1'b0;
      Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
          <= 1'b0;
    end
    else if ( operator_32_8_true_AC_TRN_AC_WRAP_2_and_27_cse ) begin
      Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_2_tmp;
      Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_3_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= 1'b0;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_13_cse & and_dcpl_51 & and_dcpl_47
        & (~ operator_32_8_true_AC_TRN_AC_WRAP_2_less_1_tmp) ) begin
      Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= $signed({1'b0, 26'b10000000000000000000000000}) < $signed(({nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
          , nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0}));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= 1'b0;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_13_cse & and_dcpl_51 & and_dcpl_47
        & (~ operator_32_8_true_AC_TRN_AC_WRAP_2_less_tmp) ) begin
      Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= $signed({1'b0, 26'b10000000000000000000000000}) < $signed(({nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31
          , nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0}));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
          <= 1'b0;
      Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
          <= 1'b0;
    end
    else if ( operator_32_8_true_AC_TRN_AC_WRAP_2_and_29_cse ) begin
      Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_tmp;
      Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_2_less_1_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_asn_262_itm <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~ or_dcpl_440) & or_71_cse ) begin
      while_asn_262_itm <= is_start_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_RunInst_switch_lp_and_16_tmp <= 1'b0;
      ActUnit_RunInst_switch_lp_and_32_tmp <= 1'b0;
    end
    else if ( ActUnit_RunInst_switch_lp_and_808_cse ) begin
      ActUnit_RunInst_switch_lp_and_16_tmp <= MUX_s_1_2_2(ActUnit_RunInst_switch_lp_equal_tmp_9,
          ActUnit_RunInst_switch_lp_and_16_tmp_mx0w1, and_dcpl_788);
      ActUnit_RunInst_switch_lp_and_32_tmp <= MUX_s_1_2_2(ActUnit_RunInst_switch_lp_equal_tmp_1_mx0w0,
          ActUnit_RunInst_switch_lp_and_32_tmp_mx0w1, and_dcpl_788);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva
          <= 1'b0;
    end
    else if ( ActUnitRun_wen & (((ActUnit_RunInst_case_2_for_i_4_0_sva_2[4]) & ((~(((is_start_sva
        | (~ (fsm_output[0]))) & (fsm_output[2])) | (fsm_output[3]) | (fsm_output[1])))
        | (fsm_output[4]))) | and_dcpl_554 | ActUnit_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva_mx0c2
        | ActUnit_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva_mx0c3
        | and_dcpl_814) ) begin
      ActUnit_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva
          <= MUX1HOT_s_1_4_2(ActUnit_RunInst_switch_lp_equal_tmp_3_mx0w0, start_PopNB_mioi_return_rsc_z_mxwt,
          ActUnit_CheckStart_if_ActUnit_CheckStart_if_and_itm_1, act_config_InstIncr_act_config_InstIncr_if_and_svs_1,
          {and_dcpl_554 , ActUnit_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva_mx0c2
          , ActUnit_RunInst_switch_lp_or_3_nl , and_dcpl_814});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_for_i_4_0_sva_3_0 <= 4'b0000;
    end
    else if ( ActUnitRun_wen & ((~ (ActUnit_RunInst_case_2_for_i_4_0_sva_2[4])) |
        ActUnit_PushOutput_if_for_i_4_0_sva_3_0_mx0c0 | (mux_213_nl & nor_734_cse))
        ) begin
      ActUnit_PushOutput_if_for_i_4_0_sva_3_0 <= MUX_v_4_2_2(4'b0000, (ActUnit_RunInst_case_2_for_i_4_0_sva_2[3:0]),
          ActUnit_PushOutput_if_for_i_not_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_0_sva_8_31 <= 1'b0;
      act_regs_data_0_0_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_64_ssc ) begin
      act_regs_data_0_0_sva_8_31 <= MUX1HOT_s_1_4_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_31,
          nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_68_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_0_0_sva_dfm_2_31, {and_dcpl_557 , and_dcpl_852 , act_regs_data_and_404_ssc
          , act_regs_data_and_405_ssc});
      act_regs_data_0_0_sva_8_30_0 <= MUX1HOT_v_31_4_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_30_0,
          nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_141_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_0_0_sva_dfm_2_30_0, {and_dcpl_557 , and_dcpl_852 , act_regs_data_and_404_ssc
          , act_regs_data_and_405_ssc});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_1_sva_8_31 <= 1'b0;
      act_regs_data_0_1_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_65_ssc ) begin
      act_regs_data_0_1_sva_8_31 <= act_regs_data_mux1h_74_nl & (~ and_dcpl_554);
      act_regs_data_0_1_sva_8_30_0 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          act_regs_data_mux1h_575_nl, not_3696_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_10_sva_8_31 <= 1'b0;
      act_regs_data_0_10_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_66_ssc ) begin
      act_regs_data_0_10_sva_8_31 <= act_regs_data_mux1h_79_nl & (~ and_dcpl_554);
      act_regs_data_0_10_sva_8_30_0 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          act_regs_data_mux1h_567_nl, not_3697_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_11_sva_8_31 <= 1'b0;
      act_regs_data_0_11_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_67_ssc ) begin
      act_regs_data_0_11_sva_8_31 <= act_regs_data_mux1h_84_nl & (~ and_dcpl_554);
      act_regs_data_0_11_sva_8_30_0 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          act_regs_data_mux1h_566_nl, not_3698_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_12_sva_8_31 <= 1'b0;
      act_regs_data_0_12_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_68_ssc ) begin
      act_regs_data_0_12_sva_8_31 <= act_regs_data_mux1h_89_nl & (~ and_dcpl_554);
      act_regs_data_0_12_sva_8_30_0 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          act_regs_data_mux1h_565_nl, not_3699_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_13_sva_8_31 <= 1'b0;
      act_regs_data_0_13_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_69_ssc ) begin
      act_regs_data_0_13_sva_8_31 <= act_regs_data_mux1h_94_nl & (~ and_dcpl_554);
      act_regs_data_0_13_sva_8_30_0 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          act_regs_data_mux1h_564_nl, not_3700_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_14_sva_8_31 <= 1'b0;
      act_regs_data_0_14_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_70_ssc ) begin
      act_regs_data_0_14_sva_8_31 <= act_regs_data_mux1h_99_nl & (~ and_dcpl_554);
      act_regs_data_0_14_sva_8_30_0 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          act_regs_data_mux1h_563_nl, not_3701_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_15_sva_8_31 <= 1'b0;
      act_regs_data_0_15_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_71_ssc ) begin
      act_regs_data_0_15_sva_8_31 <= act_regs_data_mux1h_104_nl & (~ and_dcpl_554);
      act_regs_data_0_15_sva_8_30_0 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          act_regs_data_mux1h_562_nl, not_3702_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_2_sva_8_31 <= 1'b0;
      act_regs_data_0_2_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_72_ssc ) begin
      act_regs_data_0_2_sva_8_31 <= act_regs_data_mux1h_109_nl & (~ and_dcpl_554);
      act_regs_data_0_2_sva_8_30_0 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          act_regs_data_mux1h_574_nl, not_3703_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_3_sva_8_31 <= 1'b0;
      act_regs_data_0_3_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_73_ssc ) begin
      act_regs_data_0_3_sva_8_31 <= act_regs_data_mux1h_114_nl & (~ and_dcpl_554);
      act_regs_data_0_3_sva_8_30_0 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          act_regs_data_mux1h_573_nl, not_3704_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_4_sva_8_31 <= 1'b0;
      act_regs_data_0_4_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_74_ssc ) begin
      act_regs_data_0_4_sva_8_31 <= act_regs_data_mux1h_119_nl & (~ and_dcpl_554);
      act_regs_data_0_4_sva_8_30_0 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          act_regs_data_mux1h_572_nl, not_3705_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_5_sva_8_31 <= 1'b0;
      act_regs_data_0_5_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_75_ssc ) begin
      act_regs_data_0_5_sva_8_31 <= act_regs_data_mux1h_124_nl & (~ and_dcpl_554);
      act_regs_data_0_5_sva_8_30_0 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          act_regs_data_mux1h_571_nl, not_3706_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_6_sva_8_31 <= 1'b0;
      act_regs_data_0_6_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_76_ssc ) begin
      act_regs_data_0_6_sva_8_31 <= act_regs_data_mux1h_129_nl & (~ and_dcpl_554);
      act_regs_data_0_6_sva_8_30_0 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          act_regs_data_mux1h_570_nl, not_3707_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_7_sva_8_31 <= 1'b0;
      act_regs_data_0_7_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_77_ssc ) begin
      act_regs_data_0_7_sva_8_31 <= act_regs_data_mux1h_134_nl & (~ and_dcpl_554);
      act_regs_data_0_7_sva_8_30_0 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          act_regs_data_mux1h_569_nl, not_3708_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_8_sva_8_31 <= 1'b0;
      act_regs_data_0_8_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_78_ssc ) begin
      act_regs_data_0_8_sva_8_31 <= act_regs_data_mux1h_139_nl & (~ and_dcpl_554);
      act_regs_data_0_8_sva_8_30_0 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          act_regs_data_mux1h_568_nl, not_3709_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_449 | and_dcpl_901)) | and_dcpl_557 |
        and_dcpl_900 | and_dcpl_852) ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_31 <= MUX1HOT_s_1_4_2(ActUnit_RunInst_case_2_for_ActUnit_RunInst_case_2_for_and_nl,
          Gelu_for_Gelu_for_and_11_nl, ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_2_31,
          nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_6_nl, {and_dcpl_557
          , and_dcpl_900 , and_dcpl_832 , and_dcpl_852});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1225_tmp ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_30_0 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_90_nl, nor_771_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_config_inst_counter_sva_dfm_3 <= 5'b00000;
    end
    else if ( ActUnitRun_wen & mux_217_nl ) begin
      act_config_inst_counter_sva_dfm_3 <= MUX1HOT_v_5_3_2(act_read_addrs_sva_2_mx0w0,
          ({{4{ActUnit_DecodeAxiRead_unequal_tmp_1}}, ActUnit_DecodeAxiRead_unequal_tmp_1}),
          act_config_inst_counter_sva, {nor_340_nl , and_1140_nl , or_996_tmp});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_read_req_valid_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( ActUnitRun_wen & (and_dcpl_909 | and_dcpl_829) ) begin
      act_read_req_valid_lpi_1_dfm_6 <= MUX_s_1_2_2(ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_2_tmp,
          ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_5_nl, and_dcpl_829);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_read_for_mux_15_itm <= 32'b00000000000000000000000000000000;
      act_mem_banks_read_for_mux_14_itm <= 32'b00000000000000000000000000000000;
      act_mem_banks_read_for_mux_13_itm <= 32'b00000000000000000000000000000000;
      act_mem_banks_read_for_mux_12_itm <= 32'b00000000000000000000000000000000;
      act_mem_banks_read_for_mux_11_itm <= 32'b00000000000000000000000000000000;
      act_mem_banks_read_for_mux_10_itm <= 32'b00000000000000000000000000000000;
      act_mem_banks_read_for_mux_9_itm <= 32'b00000000000000000000000000000000;
      act_mem_banks_read_for_mux_8_itm <= 32'b00000000000000000000000000000000;
      act_mem_banks_read_for_mux_7_itm <= 32'b00000000000000000000000000000000;
      act_mem_banks_read_for_mux_6_itm <= 32'b00000000000000000000000000000000;
      act_mem_banks_read_for_mux_5_itm <= 32'b00000000000000000000000000000000;
      act_mem_banks_read_for_mux_4_itm <= 32'b00000000000000000000000000000000;
      act_mem_banks_read_for_mux_3_itm <= 32'b00000000000000000000000000000000;
      act_mem_banks_read_for_mux_2_itm <= 32'b00000000000000000000000000000000;
      act_mem_banks_read_for_mux_1_itm <= 32'b00000000000000000000000000000000;
      act_mem_banks_read_for_mux_itm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_read_for_and_cse ) begin
      act_mem_banks_read_for_mux_15_itm <= MUX_v_32_32_2(act_mem_banks_bank_a_0_31_0_sva_dfm,
          act_mem_banks_bank_a_1_31_0_sva_dfm, act_mem_banks_bank_a_2_31_0_sva_dfm,
          act_mem_banks_bank_a_3_31_0_sva_dfm, act_mem_banks_bank_a_4_31_0_sva_dfm,
          act_mem_banks_bank_a_5_31_0_sva_dfm, act_mem_banks_bank_a_6_31_0_sva_dfm,
          act_mem_banks_bank_a_7_31_0_sva_dfm, act_mem_banks_bank_a_8_31_0_sva_dfm,
          act_mem_banks_bank_a_9_31_0_sva_dfm, act_mem_banks_bank_a_10_31_0_sva_dfm,
          act_mem_banks_bank_a_11_31_0_sva_dfm, act_mem_banks_bank_a_12_31_0_sva_dfm,
          act_mem_banks_bank_a_13_31_0_sva_dfm, act_mem_banks_bank_a_14_31_0_sva_dfm,
          act_mem_banks_bank_a_15_31_0_sva_dfm, act_mem_banks_bank_a_16_31_0_sva_dfm,
          act_mem_banks_bank_a_17_31_0_sva_dfm, act_mem_banks_bank_a_18_31_0_sva_dfm,
          act_mem_banks_bank_a_19_31_0_sva_dfm, act_mem_banks_bank_a_20_31_0_sva_dfm,
          act_mem_banks_bank_a_21_31_0_sva_dfm, act_mem_banks_bank_a_22_31_0_sva_dfm,
          act_mem_banks_bank_a_23_31_0_sva_dfm, act_mem_banks_bank_a_24_31_0_sva_dfm,
          act_mem_banks_bank_a_25_31_0_sva_dfm, act_mem_banks_bank_a_26_31_0_sva_dfm,
          act_mem_banks_bank_a_27_31_0_sva_dfm, act_mem_banks_bank_a_28_31_0_sva_dfm,
          act_mem_banks_bank_a_29_31_0_sva_dfm, act_mem_banks_bank_a_30_31_0_sva_dfm,
          act_mem_banks_bank_a_31_31_0_sva_dfm, while_mux_53_ssc_mx0);
      act_mem_banks_read_for_mux_14_itm <= MUX_v_32_32_2(act_mem_banks_bank_a_0_63_32_sva_dfm,
          act_mem_banks_bank_a_1_63_32_sva_dfm, act_mem_banks_bank_a_2_63_32_sva_dfm,
          act_mem_banks_bank_a_3_63_32_sva_dfm, act_mem_banks_bank_a_4_63_32_sva_dfm,
          act_mem_banks_bank_a_5_63_32_sva_dfm, act_mem_banks_bank_a_6_63_32_sva_dfm,
          act_mem_banks_bank_a_7_63_32_sva_dfm, act_mem_banks_bank_a_8_63_32_sva_dfm,
          act_mem_banks_bank_a_9_63_32_sva_dfm, act_mem_banks_bank_a_10_63_32_sva_dfm,
          act_mem_banks_bank_a_11_63_32_sva_dfm, act_mem_banks_bank_a_12_63_32_sva_dfm,
          act_mem_banks_bank_a_13_63_32_sva_dfm, act_mem_banks_bank_a_14_63_32_sva_dfm,
          act_mem_banks_bank_a_15_63_32_sva_dfm, act_mem_banks_bank_a_16_63_32_sva_dfm,
          act_mem_banks_bank_a_17_63_32_sva_dfm, act_mem_banks_bank_a_18_63_32_sva_dfm,
          act_mem_banks_bank_a_19_63_32_sva_dfm, act_mem_banks_bank_a_20_63_32_sva_dfm,
          act_mem_banks_bank_a_21_63_32_sva_dfm, act_mem_banks_bank_a_22_63_32_sva_dfm,
          act_mem_banks_bank_a_23_63_32_sva_dfm, act_mem_banks_bank_a_24_63_32_sva_dfm,
          act_mem_banks_bank_a_25_63_32_sva_dfm, act_mem_banks_bank_a_26_63_32_sva_dfm,
          act_mem_banks_bank_a_27_63_32_sva_dfm, act_mem_banks_bank_a_28_63_32_sva_dfm,
          act_mem_banks_bank_a_29_63_32_sva_dfm, act_mem_banks_bank_a_30_63_32_sva_dfm,
          act_mem_banks_bank_a_31_63_32_sva_dfm, while_mux_53_ssc_mx0);
      act_mem_banks_read_for_mux_13_itm <= MUX_v_32_32_2(act_mem_banks_bank_a_0_95_64_sva_dfm,
          act_mem_banks_bank_a_1_95_64_sva_dfm, act_mem_banks_bank_a_2_95_64_sva_dfm,
          act_mem_banks_bank_a_3_95_64_sva_dfm, act_mem_banks_bank_a_4_95_64_sva_dfm,
          act_mem_banks_bank_a_5_95_64_sva_dfm, act_mem_banks_bank_a_6_95_64_sva_dfm,
          act_mem_banks_bank_a_7_95_64_sva_dfm, act_mem_banks_bank_a_8_95_64_sva_dfm,
          act_mem_banks_bank_a_9_95_64_sva_dfm, act_mem_banks_bank_a_10_95_64_sva_dfm,
          act_mem_banks_bank_a_11_95_64_sva_dfm, act_mem_banks_bank_a_12_95_64_sva_dfm,
          act_mem_banks_bank_a_13_95_64_sva_dfm, act_mem_banks_bank_a_14_95_64_sva_dfm,
          act_mem_banks_bank_a_15_95_64_sva_dfm, act_mem_banks_bank_a_16_95_64_sva_dfm,
          act_mem_banks_bank_a_17_95_64_sva_dfm, act_mem_banks_bank_a_18_95_64_sva_dfm,
          act_mem_banks_bank_a_19_95_64_sva_dfm, act_mem_banks_bank_a_20_95_64_sva_dfm,
          act_mem_banks_bank_a_21_95_64_sva_dfm, act_mem_banks_bank_a_22_95_64_sva_dfm,
          act_mem_banks_bank_a_23_95_64_sva_dfm, act_mem_banks_bank_a_24_95_64_sva_dfm,
          act_mem_banks_bank_a_25_95_64_sva_dfm, act_mem_banks_bank_a_26_95_64_sva_dfm,
          act_mem_banks_bank_a_27_95_64_sva_dfm, act_mem_banks_bank_a_28_95_64_sva_dfm,
          act_mem_banks_bank_a_29_95_64_sva_dfm, act_mem_banks_bank_a_30_95_64_sva_dfm,
          act_mem_banks_bank_a_31_95_64_sva_dfm, while_mux_53_ssc_mx0);
      act_mem_banks_read_for_mux_12_itm <= MUX_v_32_32_2(act_mem_banks_bank_a_0_127_96_sva_dfm,
          act_mem_banks_bank_a_1_127_96_sva_dfm, act_mem_banks_bank_a_2_127_96_sva_dfm,
          act_mem_banks_bank_a_3_127_96_sva_dfm, act_mem_banks_bank_a_4_127_96_sva_dfm,
          act_mem_banks_bank_a_5_127_96_sva_dfm, act_mem_banks_bank_a_6_127_96_sva_dfm,
          act_mem_banks_bank_a_7_127_96_sva_dfm, act_mem_banks_bank_a_8_127_96_sva_dfm,
          act_mem_banks_bank_a_9_127_96_sva_dfm, act_mem_banks_bank_a_10_127_96_sva_dfm,
          act_mem_banks_bank_a_11_127_96_sva_dfm, act_mem_banks_bank_a_12_127_96_sva_dfm,
          act_mem_banks_bank_a_13_127_96_sva_dfm, act_mem_banks_bank_a_14_127_96_sva_dfm,
          act_mem_banks_bank_a_15_127_96_sva_dfm, act_mem_banks_bank_a_16_127_96_sva_dfm,
          act_mem_banks_bank_a_17_127_96_sva_dfm, act_mem_banks_bank_a_18_127_96_sva_dfm,
          act_mem_banks_bank_a_19_127_96_sva_dfm, act_mem_banks_bank_a_20_127_96_sva_dfm,
          act_mem_banks_bank_a_21_127_96_sva_dfm, act_mem_banks_bank_a_22_127_96_sva_dfm,
          act_mem_banks_bank_a_23_127_96_sva_dfm, act_mem_banks_bank_a_24_127_96_sva_dfm,
          act_mem_banks_bank_a_25_127_96_sva_dfm, act_mem_banks_bank_a_26_127_96_sva_dfm,
          act_mem_banks_bank_a_27_127_96_sva_dfm, act_mem_banks_bank_a_28_127_96_sva_dfm,
          act_mem_banks_bank_a_29_127_96_sva_dfm, act_mem_banks_bank_a_30_127_96_sva_dfm,
          act_mem_banks_bank_a_31_127_96_sva_dfm, while_mux_53_ssc_mx0);
      act_mem_banks_read_for_mux_11_itm <= MUX_v_32_32_2(act_mem_banks_bank_a_0_159_128_sva_dfm,
          act_mem_banks_bank_a_1_159_128_sva_dfm, act_mem_banks_bank_a_2_159_128_sva_dfm,
          act_mem_banks_bank_a_3_159_128_sva_dfm, act_mem_banks_bank_a_4_159_128_sva_dfm,
          act_mem_banks_bank_a_5_159_128_sva_dfm, act_mem_banks_bank_a_6_159_128_sva_dfm,
          act_mem_banks_bank_a_7_159_128_sva_dfm, act_mem_banks_bank_a_8_159_128_sva_dfm,
          act_mem_banks_bank_a_9_159_128_sva_dfm, act_mem_banks_bank_a_10_159_128_sva_dfm,
          act_mem_banks_bank_a_11_159_128_sva_dfm, act_mem_banks_bank_a_12_159_128_sva_dfm,
          act_mem_banks_bank_a_13_159_128_sva_dfm, act_mem_banks_bank_a_14_159_128_sva_dfm,
          act_mem_banks_bank_a_15_159_128_sva_dfm, act_mem_banks_bank_a_16_159_128_sva_dfm,
          act_mem_banks_bank_a_17_159_128_sva_dfm, act_mem_banks_bank_a_18_159_128_sva_dfm,
          act_mem_banks_bank_a_19_159_128_sva_dfm, act_mem_banks_bank_a_20_159_128_sva_dfm,
          act_mem_banks_bank_a_21_159_128_sva_dfm, act_mem_banks_bank_a_22_159_128_sva_dfm,
          act_mem_banks_bank_a_23_159_128_sva_dfm, act_mem_banks_bank_a_24_159_128_sva_dfm,
          act_mem_banks_bank_a_25_159_128_sva_dfm, act_mem_banks_bank_a_26_159_128_sva_dfm,
          act_mem_banks_bank_a_27_159_128_sva_dfm, act_mem_banks_bank_a_28_159_128_sva_dfm,
          act_mem_banks_bank_a_29_159_128_sva_dfm, act_mem_banks_bank_a_30_159_128_sva_dfm,
          act_mem_banks_bank_a_31_159_128_sva_dfm, while_mux_53_ssc_mx0);
      act_mem_banks_read_for_mux_10_itm <= MUX_v_32_32_2(act_mem_banks_bank_a_0_191_160_sva_dfm,
          act_mem_banks_bank_a_1_191_160_sva_dfm, act_mem_banks_bank_a_2_191_160_sva_dfm,
          act_mem_banks_bank_a_3_191_160_sva_dfm, act_mem_banks_bank_a_4_191_160_sva_dfm,
          act_mem_banks_bank_a_5_191_160_sva_dfm, act_mem_banks_bank_a_6_191_160_sva_dfm,
          act_mem_banks_bank_a_7_191_160_sva_dfm, act_mem_banks_bank_a_8_191_160_sva_dfm,
          act_mem_banks_bank_a_9_191_160_sva_dfm, act_mem_banks_bank_a_10_191_160_sva_dfm,
          act_mem_banks_bank_a_11_191_160_sva_dfm, act_mem_banks_bank_a_12_191_160_sva_dfm,
          act_mem_banks_bank_a_13_191_160_sva_dfm, act_mem_banks_bank_a_14_191_160_sva_dfm,
          act_mem_banks_bank_a_15_191_160_sva_dfm, act_mem_banks_bank_a_16_191_160_sva_dfm,
          act_mem_banks_bank_a_17_191_160_sva_dfm, act_mem_banks_bank_a_18_191_160_sva_dfm,
          act_mem_banks_bank_a_19_191_160_sva_dfm, act_mem_banks_bank_a_20_191_160_sva_dfm,
          act_mem_banks_bank_a_21_191_160_sva_dfm, act_mem_banks_bank_a_22_191_160_sva_dfm,
          act_mem_banks_bank_a_23_191_160_sva_dfm, act_mem_banks_bank_a_24_191_160_sva_dfm,
          act_mem_banks_bank_a_25_191_160_sva_dfm, act_mem_banks_bank_a_26_191_160_sva_dfm,
          act_mem_banks_bank_a_27_191_160_sva_dfm, act_mem_banks_bank_a_28_191_160_sva_dfm,
          act_mem_banks_bank_a_29_191_160_sva_dfm, act_mem_banks_bank_a_30_191_160_sva_dfm,
          act_mem_banks_bank_a_31_191_160_sva_dfm, while_mux_53_ssc_mx0);
      act_mem_banks_read_for_mux_9_itm <= MUX_v_32_32_2(act_mem_banks_bank_a_0_223_192_sva_dfm,
          act_mem_banks_bank_a_1_223_192_sva_dfm, act_mem_banks_bank_a_2_223_192_sva_dfm,
          act_mem_banks_bank_a_3_223_192_sva_dfm, act_mem_banks_bank_a_4_223_192_sva_dfm,
          act_mem_banks_bank_a_5_223_192_sva_dfm, act_mem_banks_bank_a_6_223_192_sva_dfm,
          act_mem_banks_bank_a_7_223_192_sva_dfm, act_mem_banks_bank_a_8_223_192_sva_dfm,
          act_mem_banks_bank_a_9_223_192_sva_dfm, act_mem_banks_bank_a_10_223_192_sva_dfm,
          act_mem_banks_bank_a_11_223_192_sva_dfm, act_mem_banks_bank_a_12_223_192_sva_dfm,
          act_mem_banks_bank_a_13_223_192_sva_dfm, act_mem_banks_bank_a_14_223_192_sva_dfm,
          act_mem_banks_bank_a_15_223_192_sva_dfm, act_mem_banks_bank_a_16_223_192_sva_dfm,
          act_mem_banks_bank_a_17_223_192_sva_dfm, act_mem_banks_bank_a_18_223_192_sva_dfm,
          act_mem_banks_bank_a_19_223_192_sva_dfm, act_mem_banks_bank_a_20_223_192_sva_dfm,
          act_mem_banks_bank_a_21_223_192_sva_dfm, act_mem_banks_bank_a_22_223_192_sva_dfm,
          act_mem_banks_bank_a_23_223_192_sva_dfm, act_mem_banks_bank_a_24_223_192_sva_dfm,
          act_mem_banks_bank_a_25_223_192_sva_dfm, act_mem_banks_bank_a_26_223_192_sva_dfm,
          act_mem_banks_bank_a_27_223_192_sva_dfm, act_mem_banks_bank_a_28_223_192_sva_dfm,
          act_mem_banks_bank_a_29_223_192_sva_dfm, act_mem_banks_bank_a_30_223_192_sva_dfm,
          act_mem_banks_bank_a_31_223_192_sva_dfm, while_mux_53_ssc_mx0);
      act_mem_banks_read_for_mux_8_itm <= MUX_v_32_32_2(act_mem_banks_bank_a_0_255_224_sva_dfm,
          act_mem_banks_bank_a_1_255_224_sva_dfm, act_mem_banks_bank_a_2_255_224_sva_dfm,
          act_mem_banks_bank_a_3_255_224_sva_dfm, act_mem_banks_bank_a_4_255_224_sva_dfm,
          act_mem_banks_bank_a_5_255_224_sva_dfm, act_mem_banks_bank_a_6_255_224_sva_dfm,
          act_mem_banks_bank_a_7_255_224_sva_dfm, act_mem_banks_bank_a_8_255_224_sva_dfm,
          act_mem_banks_bank_a_9_255_224_sva_dfm, act_mem_banks_bank_a_10_255_224_sva_dfm,
          act_mem_banks_bank_a_11_255_224_sva_dfm, act_mem_banks_bank_a_12_255_224_sva_dfm,
          act_mem_banks_bank_a_13_255_224_sva_dfm, act_mem_banks_bank_a_14_255_224_sva_dfm,
          act_mem_banks_bank_a_15_255_224_sva_dfm, act_mem_banks_bank_a_16_255_224_sva_dfm,
          act_mem_banks_bank_a_17_255_224_sva_dfm, act_mem_banks_bank_a_18_255_224_sva_dfm,
          act_mem_banks_bank_a_19_255_224_sva_dfm, act_mem_banks_bank_a_20_255_224_sva_dfm,
          act_mem_banks_bank_a_21_255_224_sva_dfm, act_mem_banks_bank_a_22_255_224_sva_dfm,
          act_mem_banks_bank_a_23_255_224_sva_dfm, act_mem_banks_bank_a_24_255_224_sva_dfm,
          act_mem_banks_bank_a_25_255_224_sva_dfm, act_mem_banks_bank_a_26_255_224_sva_dfm,
          act_mem_banks_bank_a_27_255_224_sva_dfm, act_mem_banks_bank_a_28_255_224_sva_dfm,
          act_mem_banks_bank_a_29_255_224_sva_dfm, act_mem_banks_bank_a_30_255_224_sva_dfm,
          act_mem_banks_bank_a_31_255_224_sva_dfm, while_mux_53_ssc_mx0);
      act_mem_banks_read_for_mux_7_itm <= MUX_v_32_32_2(act_mem_banks_bank_a_0_287_256_sva_dfm,
          act_mem_banks_bank_a_1_287_256_sva_dfm, act_mem_banks_bank_a_2_287_256_sva_dfm,
          act_mem_banks_bank_a_3_287_256_sva_dfm, act_mem_banks_bank_a_4_287_256_sva_dfm,
          act_mem_banks_bank_a_5_287_256_sva_dfm, act_mem_banks_bank_a_6_287_256_sva_dfm,
          act_mem_banks_bank_a_7_287_256_sva_dfm, act_mem_banks_bank_a_8_287_256_sva_dfm,
          act_mem_banks_bank_a_9_287_256_sva_dfm, act_mem_banks_bank_a_10_287_256_sva_dfm,
          act_mem_banks_bank_a_11_287_256_sva_dfm, act_mem_banks_bank_a_12_287_256_sva_dfm,
          act_mem_banks_bank_a_13_287_256_sva_dfm, act_mem_banks_bank_a_14_287_256_sva_dfm,
          act_mem_banks_bank_a_15_287_256_sva_dfm, act_mem_banks_bank_a_16_287_256_sva_dfm,
          act_mem_banks_bank_a_17_287_256_sva_dfm, act_mem_banks_bank_a_18_287_256_sva_dfm,
          act_mem_banks_bank_a_19_287_256_sva_dfm, act_mem_banks_bank_a_20_287_256_sva_dfm,
          act_mem_banks_bank_a_21_287_256_sva_dfm, act_mem_banks_bank_a_22_287_256_sva_dfm,
          act_mem_banks_bank_a_23_287_256_sva_dfm, act_mem_banks_bank_a_24_287_256_sva_dfm,
          act_mem_banks_bank_a_25_287_256_sva_dfm, act_mem_banks_bank_a_26_287_256_sva_dfm,
          act_mem_banks_bank_a_27_287_256_sva_dfm, act_mem_banks_bank_a_28_287_256_sva_dfm,
          act_mem_banks_bank_a_29_287_256_sva_dfm, act_mem_banks_bank_a_30_287_256_sva_dfm,
          act_mem_banks_bank_a_31_287_256_sva_dfm, while_mux_53_ssc_mx0);
      act_mem_banks_read_for_mux_6_itm <= MUX_v_32_32_2(act_mem_banks_bank_a_0_319_288_sva_dfm,
          act_mem_banks_bank_a_1_319_288_sva_dfm, act_mem_banks_bank_a_2_319_288_sva_dfm,
          act_mem_banks_bank_a_3_319_288_sva_dfm, act_mem_banks_bank_a_4_319_288_sva_dfm,
          act_mem_banks_bank_a_5_319_288_sva_dfm, act_mem_banks_bank_a_6_319_288_sva_dfm,
          act_mem_banks_bank_a_7_319_288_sva_dfm, act_mem_banks_bank_a_8_319_288_sva_dfm,
          act_mem_banks_bank_a_9_319_288_sva_dfm, act_mem_banks_bank_a_10_319_288_sva_dfm,
          act_mem_banks_bank_a_11_319_288_sva_dfm, act_mem_banks_bank_a_12_319_288_sva_dfm,
          act_mem_banks_bank_a_13_319_288_sva_dfm, act_mem_banks_bank_a_14_319_288_sva_dfm,
          act_mem_banks_bank_a_15_319_288_sva_dfm, act_mem_banks_bank_a_16_319_288_sva_dfm,
          act_mem_banks_bank_a_17_319_288_sva_dfm, act_mem_banks_bank_a_18_319_288_sva_dfm,
          act_mem_banks_bank_a_19_319_288_sva_dfm, act_mem_banks_bank_a_20_319_288_sva_dfm,
          act_mem_banks_bank_a_21_319_288_sva_dfm, act_mem_banks_bank_a_22_319_288_sva_dfm,
          act_mem_banks_bank_a_23_319_288_sva_dfm, act_mem_banks_bank_a_24_319_288_sva_dfm,
          act_mem_banks_bank_a_25_319_288_sva_dfm, act_mem_banks_bank_a_26_319_288_sva_dfm,
          act_mem_banks_bank_a_27_319_288_sva_dfm, act_mem_banks_bank_a_28_319_288_sva_dfm,
          act_mem_banks_bank_a_29_319_288_sva_dfm, act_mem_banks_bank_a_30_319_288_sva_dfm,
          act_mem_banks_bank_a_31_319_288_sva_dfm, while_mux_53_ssc_mx0);
      act_mem_banks_read_for_mux_5_itm <= MUX_v_32_32_2(act_mem_banks_bank_a_0_351_320_sva_dfm,
          act_mem_banks_bank_a_1_351_320_sva_dfm, act_mem_banks_bank_a_2_351_320_sva_dfm,
          act_mem_banks_bank_a_3_351_320_sva_dfm, act_mem_banks_bank_a_4_351_320_sva_dfm,
          act_mem_banks_bank_a_5_351_320_sva_dfm, act_mem_banks_bank_a_6_351_320_sva_dfm,
          act_mem_banks_bank_a_7_351_320_sva_dfm, act_mem_banks_bank_a_8_351_320_sva_dfm,
          act_mem_banks_bank_a_9_351_320_sva_dfm, act_mem_banks_bank_a_10_351_320_sva_dfm,
          act_mem_banks_bank_a_11_351_320_sva_dfm, act_mem_banks_bank_a_12_351_320_sva_dfm,
          act_mem_banks_bank_a_13_351_320_sva_dfm, act_mem_banks_bank_a_14_351_320_sva_dfm,
          act_mem_banks_bank_a_15_351_320_sva_dfm, act_mem_banks_bank_a_16_351_320_sva_dfm,
          act_mem_banks_bank_a_17_351_320_sva_dfm, act_mem_banks_bank_a_18_351_320_sva_dfm,
          act_mem_banks_bank_a_19_351_320_sva_dfm, act_mem_banks_bank_a_20_351_320_sva_dfm,
          act_mem_banks_bank_a_21_351_320_sva_dfm, act_mem_banks_bank_a_22_351_320_sva_dfm,
          act_mem_banks_bank_a_23_351_320_sva_dfm, act_mem_banks_bank_a_24_351_320_sva_dfm,
          act_mem_banks_bank_a_25_351_320_sva_dfm, act_mem_banks_bank_a_26_351_320_sva_dfm,
          act_mem_banks_bank_a_27_351_320_sva_dfm, act_mem_banks_bank_a_28_351_320_sva_dfm,
          act_mem_banks_bank_a_29_351_320_sva_dfm, act_mem_banks_bank_a_30_351_320_sva_dfm,
          act_mem_banks_bank_a_31_351_320_sva_dfm, while_mux_53_ssc_mx0);
      act_mem_banks_read_for_mux_4_itm <= MUX_v_32_32_2(act_mem_banks_bank_a_0_383_352_sva_dfm,
          act_mem_banks_bank_a_1_383_352_sva_dfm, act_mem_banks_bank_a_2_383_352_sva_dfm,
          act_mem_banks_bank_a_3_383_352_sva_dfm, act_mem_banks_bank_a_4_383_352_sva_dfm,
          act_mem_banks_bank_a_5_383_352_sva_dfm, act_mem_banks_bank_a_6_383_352_sva_dfm,
          act_mem_banks_bank_a_7_383_352_sva_dfm, act_mem_banks_bank_a_8_383_352_sva_dfm,
          act_mem_banks_bank_a_9_383_352_sva_dfm, act_mem_banks_bank_a_10_383_352_sva_dfm,
          act_mem_banks_bank_a_11_383_352_sva_dfm, act_mem_banks_bank_a_12_383_352_sva_dfm,
          act_mem_banks_bank_a_13_383_352_sva_dfm, act_mem_banks_bank_a_14_383_352_sva_dfm,
          act_mem_banks_bank_a_15_383_352_sva_dfm, act_mem_banks_bank_a_16_383_352_sva_dfm,
          act_mem_banks_bank_a_17_383_352_sva_dfm, act_mem_banks_bank_a_18_383_352_sva_dfm,
          act_mem_banks_bank_a_19_383_352_sva_dfm, act_mem_banks_bank_a_20_383_352_sva_dfm,
          act_mem_banks_bank_a_21_383_352_sva_dfm, act_mem_banks_bank_a_22_383_352_sva_dfm,
          act_mem_banks_bank_a_23_383_352_sva_dfm, act_mem_banks_bank_a_24_383_352_sva_dfm,
          act_mem_banks_bank_a_25_383_352_sva_dfm, act_mem_banks_bank_a_26_383_352_sva_dfm,
          act_mem_banks_bank_a_27_383_352_sva_dfm, act_mem_banks_bank_a_28_383_352_sva_dfm,
          act_mem_banks_bank_a_29_383_352_sva_dfm, act_mem_banks_bank_a_30_383_352_sva_dfm,
          act_mem_banks_bank_a_31_383_352_sva_dfm, while_mux_53_ssc_mx0);
      act_mem_banks_read_for_mux_3_itm <= MUX_v_32_32_2(act_mem_banks_bank_a_0_415_384_sva_dfm,
          act_mem_banks_bank_a_1_415_384_sva_dfm, act_mem_banks_bank_a_2_415_384_sva_dfm,
          act_mem_banks_bank_a_3_415_384_sva_dfm, act_mem_banks_bank_a_4_415_384_sva_dfm,
          act_mem_banks_bank_a_5_415_384_sva_dfm, act_mem_banks_bank_a_6_415_384_sva_dfm,
          act_mem_banks_bank_a_7_415_384_sva_dfm, act_mem_banks_bank_a_8_415_384_sva_dfm,
          act_mem_banks_bank_a_9_415_384_sva_dfm, act_mem_banks_bank_a_10_415_384_sva_dfm,
          act_mem_banks_bank_a_11_415_384_sva_dfm, act_mem_banks_bank_a_12_415_384_sva_dfm,
          act_mem_banks_bank_a_13_415_384_sva_dfm, act_mem_banks_bank_a_14_415_384_sva_dfm,
          act_mem_banks_bank_a_15_415_384_sva_dfm, act_mem_banks_bank_a_16_415_384_sva_dfm,
          act_mem_banks_bank_a_17_415_384_sva_dfm, act_mem_banks_bank_a_18_415_384_sva_dfm,
          act_mem_banks_bank_a_19_415_384_sva_dfm, act_mem_banks_bank_a_20_415_384_sva_dfm,
          act_mem_banks_bank_a_21_415_384_sva_dfm, act_mem_banks_bank_a_22_415_384_sva_dfm,
          act_mem_banks_bank_a_23_415_384_sva_dfm, act_mem_banks_bank_a_24_415_384_sva_dfm,
          act_mem_banks_bank_a_25_415_384_sva_dfm, act_mem_banks_bank_a_26_415_384_sva_dfm,
          act_mem_banks_bank_a_27_415_384_sva_dfm, act_mem_banks_bank_a_28_415_384_sva_dfm,
          act_mem_banks_bank_a_29_415_384_sva_dfm, act_mem_banks_bank_a_30_415_384_sva_dfm,
          act_mem_banks_bank_a_31_415_384_sva_dfm, while_mux_53_ssc_mx0);
      act_mem_banks_read_for_mux_2_itm <= MUX_v_32_32_2(act_mem_banks_bank_a_0_447_416_sva_dfm,
          act_mem_banks_bank_a_1_447_416_sva_dfm, act_mem_banks_bank_a_2_447_416_sva_dfm,
          act_mem_banks_bank_a_3_447_416_sva_dfm, act_mem_banks_bank_a_4_447_416_sva_dfm,
          act_mem_banks_bank_a_5_447_416_sva_dfm, act_mem_banks_bank_a_6_447_416_sva_dfm,
          act_mem_banks_bank_a_7_447_416_sva_dfm, act_mem_banks_bank_a_8_447_416_sva_dfm,
          act_mem_banks_bank_a_9_447_416_sva_dfm, act_mem_banks_bank_a_10_447_416_sva_dfm,
          act_mem_banks_bank_a_11_447_416_sva_dfm, act_mem_banks_bank_a_12_447_416_sva_dfm,
          act_mem_banks_bank_a_13_447_416_sva_dfm, act_mem_banks_bank_a_14_447_416_sva_dfm,
          act_mem_banks_bank_a_15_447_416_sva_dfm, act_mem_banks_bank_a_16_447_416_sva_dfm,
          act_mem_banks_bank_a_17_447_416_sva_dfm, act_mem_banks_bank_a_18_447_416_sva_dfm,
          act_mem_banks_bank_a_19_447_416_sva_dfm, act_mem_banks_bank_a_20_447_416_sva_dfm,
          act_mem_banks_bank_a_21_447_416_sva_dfm, act_mem_banks_bank_a_22_447_416_sva_dfm,
          act_mem_banks_bank_a_23_447_416_sva_dfm, act_mem_banks_bank_a_24_447_416_sva_dfm,
          act_mem_banks_bank_a_25_447_416_sva_dfm, act_mem_banks_bank_a_26_447_416_sva_dfm,
          act_mem_banks_bank_a_27_447_416_sva_dfm, act_mem_banks_bank_a_28_447_416_sva_dfm,
          act_mem_banks_bank_a_29_447_416_sva_dfm, act_mem_banks_bank_a_30_447_416_sva_dfm,
          act_mem_banks_bank_a_31_447_416_sva_dfm, while_mux_53_ssc_mx0);
      act_mem_banks_read_for_mux_1_itm <= MUX_v_32_32_2(act_mem_banks_bank_a_0_479_448_sva_dfm,
          act_mem_banks_bank_a_1_479_448_sva_dfm, act_mem_banks_bank_a_2_479_448_sva_dfm,
          act_mem_banks_bank_a_3_479_448_sva_dfm, act_mem_banks_bank_a_4_479_448_sva_dfm,
          act_mem_banks_bank_a_5_479_448_sva_dfm, act_mem_banks_bank_a_6_479_448_sva_dfm,
          act_mem_banks_bank_a_7_479_448_sva_dfm, act_mem_banks_bank_a_8_479_448_sva_dfm,
          act_mem_banks_bank_a_9_479_448_sva_dfm, act_mem_banks_bank_a_10_479_448_sva_dfm,
          act_mem_banks_bank_a_11_479_448_sva_dfm, act_mem_banks_bank_a_12_479_448_sva_dfm,
          act_mem_banks_bank_a_13_479_448_sva_dfm, act_mem_banks_bank_a_14_479_448_sva_dfm,
          act_mem_banks_bank_a_15_479_448_sva_dfm, act_mem_banks_bank_a_16_479_448_sva_dfm,
          act_mem_banks_bank_a_17_479_448_sva_dfm, act_mem_banks_bank_a_18_479_448_sva_dfm,
          act_mem_banks_bank_a_19_479_448_sva_dfm, act_mem_banks_bank_a_20_479_448_sva_dfm,
          act_mem_banks_bank_a_21_479_448_sva_dfm, act_mem_banks_bank_a_22_479_448_sva_dfm,
          act_mem_banks_bank_a_23_479_448_sva_dfm, act_mem_banks_bank_a_24_479_448_sva_dfm,
          act_mem_banks_bank_a_25_479_448_sva_dfm, act_mem_banks_bank_a_26_479_448_sva_dfm,
          act_mem_banks_bank_a_27_479_448_sva_dfm, act_mem_banks_bank_a_28_479_448_sva_dfm,
          act_mem_banks_bank_a_29_479_448_sva_dfm, act_mem_banks_bank_a_30_479_448_sva_dfm,
          act_mem_banks_bank_a_31_479_448_sva_dfm, while_mux_53_ssc_mx0);
      act_mem_banks_read_for_mux_itm <= MUX_v_32_32_2(act_mem_banks_bank_a_0_511_480_sva_dfm,
          act_mem_banks_bank_a_1_511_480_sva_dfm, act_mem_banks_bank_a_2_511_480_sva_dfm,
          act_mem_banks_bank_a_3_511_480_sva_dfm, act_mem_banks_bank_a_4_511_480_sva_dfm,
          act_mem_banks_bank_a_5_511_480_sva_dfm, act_mem_banks_bank_a_6_511_480_sva_dfm,
          act_mem_banks_bank_a_7_511_480_sva_dfm, act_mem_banks_bank_a_8_511_480_sva_dfm,
          act_mem_banks_bank_a_9_511_480_sva_dfm, act_mem_banks_bank_a_10_511_480_sva_dfm,
          act_mem_banks_bank_a_11_511_480_sva_dfm, act_mem_banks_bank_a_12_511_480_sva_dfm,
          act_mem_banks_bank_a_13_511_480_sva_dfm, act_mem_banks_bank_a_14_511_480_sva_dfm,
          act_mem_banks_bank_a_15_511_480_sva_dfm, act_mem_banks_bank_a_16_511_480_sva_dfm,
          act_mem_banks_bank_a_17_511_480_sva_dfm, act_mem_banks_bank_a_18_511_480_sva_dfm,
          act_mem_banks_bank_a_19_511_480_sva_dfm, act_mem_banks_bank_a_20_511_480_sva_dfm,
          act_mem_banks_bank_a_21_511_480_sva_dfm, act_mem_banks_bank_a_22_511_480_sva_dfm,
          act_mem_banks_bank_a_23_511_480_sva_dfm, act_mem_banks_bank_a_24_511_480_sva_dfm,
          act_mem_banks_bank_a_25_511_480_sva_dfm, act_mem_banks_bank_a_26_511_480_sva_dfm,
          act_mem_banks_bank_a_27_511_480_sva_dfm, act_mem_banks_bank_a_28_511_480_sva_dfm,
          act_mem_banks_bank_a_29_511_480_sva_dfm, act_mem_banks_bank_a_30_511_480_sva_dfm,
          act_mem_banks_bank_a_31_511_480_sva_dfm, while_mux_53_ssc_mx0);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_0_sva_dfm_3 <= 1'b0;
      rva_out_reg_data_8_sva_dfm_3 <= 1'b0;
      rva_out_reg_data_29_24_sva_dfm_3 <= 6'b000000;
      rva_out_reg_data_39_32_sva_dfm_3 <= 8'b00000000;
      rva_out_reg_data_52_48_sva_dfm_3 <= 5'b00000;
      rva_out_reg_data_71_64_sva_dfm_3 <= 8'b00000000;
    end
    else if ( rva_out_reg_data_and_62_cse ) begin
      rva_out_reg_data_0_sva_dfm_3 <= MUX_s_1_2_2(ActUnit_DecodeAxi_mux_93_nl, ActUnit_PushOutput_if_for_and_stg_2_7_sva,
          is_start_sva);
      rva_out_reg_data_8_sva_dfm_3 <= MUX_s_1_2_2(ActUnit_DecodeAxi_mux_94_nl, Gelu_for_and_2_cse_sva,
          is_start_sva);
      rva_out_reg_data_29_24_sva_dfm_3 <= MUX1HOT_v_6_4_2(rva_out_reg_data_29_24_sva_dfm_6,
          act_config_num_inst_sva, act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_20_nl,
          (act_config_inst_regs_3_sva_dfm_5[5:0]), {while_asn_1331 , while_asn_1333
          , while_and_203_cse , while_and_204_cse});
      rva_out_reg_data_39_32_sva_dfm_3 <= MUX1HOT_v_8_4_2(rva_out_reg_data_39_32_sva_dfm_6,
          act_config_num_output_sva, act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_21_nl,
          act_config_inst_regs_4_sva_dfm_5, {while_asn_1331 , while_asn_1333 , while_and_203_cse
          , while_and_204_cse});
      rva_out_reg_data_52_48_sva_dfm_3 <= MUX1HOT_v_5_4_2(rva_out_reg_data_52_48_sva_dfm_6,
          act_config_buffer_addr_base_sva, act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_22_nl,
          (act_config_inst_regs_6_sva_dfm_5[4:0]), {while_asn_1331 , while_asn_1333
          , while_and_203_cse , while_and_204_cse});
      rva_out_reg_data_71_64_sva_dfm_3 <= MUX1HOT_v_8_4_2(rva_out_reg_data_71_64_sva_dfm_6,
          act_config_output_addr_base_sva, act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_23_nl,
          act_config_inst_regs_8_sva_dfm_5, {while_asn_1331 , while_asn_1333 , while_and_203_cse
          , while_and_204_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      w_axi_rsp_lpi_1_dfm_1 <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_423 | or_dcpl_322)) ) begin
      w_axi_rsp_lpi_1_dfm_1 <= ~(ActUnit_DecodeAxi_rva_in_reg_rw_sva_mx1 | (~ ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_mx1)
          | is_start_sva);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_RunInst_case_3_act_port_reg_data_sva <= 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ActUnit_RunInst_case_3_act_port_reg_data_and_cse & act_port_PopNB_mioi_return_rsc_z_mxwt
        & is_start_sva & ActUnit_RunInst_switch_lp_equal_tmp_2 ) begin
      ActUnit_RunInst_case_3_act_port_reg_data_sva <= act_port_PopNB_mioi_data_data_rsc_z_mxwt;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_config_output_counter_sva_dfm_3 <= 8'b00000000;
      is_incr_lpi_1_dfm_1 <= 1'b0;
      act_config_is_zero_first_sva_dfm_4 <= 1'b0;
    end
    else if ( act_config_output_counter_and_1_cse ) begin
      act_config_output_counter_sva_dfm_3 <= MUX_v_8_2_2(({{7{ActUnit_DecodeAxiRead_unequal_tmp_1}},
          ActUnit_DecodeAxiRead_unequal_tmp_1}), act_config_output_counter_sva, or_997_nl);
      is_incr_lpi_1_dfm_1 <= act_port_PopNB_mioi_return_rsc_z_mxwt | (~ ActUnit_RunInst_switch_lp_equal_tmp_2)
          | (~ is_start_sva);
      act_config_is_zero_first_sva_dfm_4 <= MUX_s_1_2_2(ActUnit_DecodeAxiWrite_mux_4_nl,
          act_config_is_zero_first_sva, and_dcpl_908);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_nor_cse <= 1'b0;
      reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_2_cse <= 1'b0;
      reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_1_cse <= 1'b0;
      reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_cse <= 1'b0;
      ActUnit_RunInst_switch_lp_and_48_tmp <= 1'b0;
      ActUnit_RunInst_switch_lp_and_tmp <= 1'b0;
      while_nor_48_itm <= 1'b0;
      while_nor_32_itm <= 1'b0;
      while_nor_16_itm <= 1'b0;
      while_nor_itm <= 1'b0;
    end
    else if ( ActUnit_RunInst_case_3_act_port_reg_data_and_cse ) begin
      reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_nor_cse <= Tanh_for_nor_cse_sva_mx0w0;
      reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_2_cse <= Tanh_for_and_2_cse_sva_mx0w0;
      reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_1_cse <= Tanh_for_and_1_cse_sva_mx0w0;
      reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_cse <= Tanh_for_and_cse_sva_mx0w0;
      ActUnit_RunInst_switch_lp_and_48_tmp <= ActUnit_RunInst_switch_lp_and_48_tmp_mx0w0;
      ActUnit_RunInst_switch_lp_and_tmp <= ActUnit_RunInst_switch_lp_and_tmp_mx0w0;
      while_nor_48_itm <= ~(ActUnit_RunInst_switch_lp_and_16_tmp | ActUnit_RunInst_switch_lp_and_32_tmp
          | ActUnit_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva
          | ActUnit_RunInst_switch_lp_nor_tmp | ((~ Tanh_for_and_2_cse_sva_mx0w0)
          & ActUnit_RunInst_switch_lp_equal_tmp_4) | ((~ Tanh_for_and_2_cse_sva_mx0w0)
          & ActUnit_RunInst_switch_lp_equal_tmp_5) | ((~ Tanh_for_and_2_cse_sva_mx0w0)
          & ActUnit_RunInst_switch_lp_equal_tmp_6) | ((~ Tanh_for_and_2_cse_sva_mx0w0)
          & ActUnit_RunInst_switch_lp_equal_tmp_7) | ((~ Tanh_for_and_2_cse_sva_mx0w0)
          & ActUnit_RunInst_switch_lp_equal_tmp_8) | ((~ ActUnit_RunInst_switch_lp_and_48_tmp_mx0w0)
          & ActUnit_RunInst_switch_lp_equal_tmp_2));
      while_nor_32_itm <= ~(ActUnit_RunInst_switch_lp_and_16_tmp | ActUnit_RunInst_switch_lp_and_32_tmp
          | ActUnit_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva
          | ActUnit_RunInst_switch_lp_nor_tmp | ((~ Tanh_for_and_cse_sva_mx0w0) &
          ActUnit_RunInst_switch_lp_equal_tmp_4) | ((~ Tanh_for_and_cse_sva_mx0w0)
          & ActUnit_RunInst_switch_lp_equal_tmp_5) | ((~ Tanh_for_and_cse_sva_mx0w0)
          & ActUnit_RunInst_switch_lp_equal_tmp_6) | ((~ Tanh_for_and_cse_sva_mx0w0)
          & ActUnit_RunInst_switch_lp_equal_tmp_7) | ((~ Tanh_for_and_cse_sva_mx0w0)
          & ActUnit_RunInst_switch_lp_equal_tmp_8) | ((~ ActUnit_RunInst_switch_lp_and_32_tmp_mx0w1)
          & ActUnit_RunInst_switch_lp_equal_tmp_2));
      while_nor_16_itm <= ~(ActUnit_RunInst_switch_lp_and_16_tmp | ActUnit_RunInst_switch_lp_and_32_tmp
          | ActUnit_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva
          | ActUnit_RunInst_switch_lp_nor_tmp | ((~ Tanh_for_and_1_cse_sva_mx0w0)
          & ActUnit_RunInst_switch_lp_equal_tmp_4) | ((~ Tanh_for_and_1_cse_sva_mx0w0)
          & ActUnit_RunInst_switch_lp_equal_tmp_5) | ((~ Tanh_for_and_1_cse_sva_mx0w0)
          & ActUnit_RunInst_switch_lp_equal_tmp_6) | ((~ Tanh_for_and_1_cse_sva_mx0w0)
          & ActUnit_RunInst_switch_lp_equal_tmp_7) | ((~ Tanh_for_and_1_cse_sva_mx0w0)
          & ActUnit_RunInst_switch_lp_equal_tmp_8) | ((~ ActUnit_RunInst_switch_lp_and_16_tmp_mx0w1)
          & ActUnit_RunInst_switch_lp_equal_tmp_2));
      while_nor_itm <= ~(ActUnit_RunInst_switch_lp_and_16_tmp | ActUnit_RunInst_switch_lp_and_32_tmp
          | ActUnit_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva
          | ActUnit_RunInst_switch_lp_nor_tmp | ((~ Tanh_for_nor_cse_sva_mx0w0) &
          ActUnit_RunInst_switch_lp_equal_tmp_4) | ((~ Tanh_for_nor_cse_sva_mx0w0)
          & ActUnit_RunInst_switch_lp_equal_tmp_5) | ((~ Tanh_for_nor_cse_sva_mx0w0)
          & ActUnit_RunInst_switch_lp_equal_tmp_6) | ((~ Tanh_for_nor_cse_sva_mx0w0)
          & ActUnit_RunInst_switch_lp_equal_tmp_7) | ((~ Tanh_for_nor_cse_sva_mx0w0)
          & ActUnit_RunInst_switch_lp_equal_tmp_8) | ((~ ActUnit_RunInst_switch_lp_and_tmp_mx0w0)
          & ActUnit_RunInst_switch_lp_equal_tmp_2));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_get_slc_2U_NVUINT8_return_2_sva <= 2'b00;
    end
    else if ( ActUnitRun_wen & (mux_tmp_214 | (fsm_output[4])) & and_dcpl_377 ) begin
      nvhls_get_slc_2U_NVUINT8_return_2_sva <= MUX_v_2_32_2((act_config_inst_regs_0_sva_dfm_5[3:2]),
          (act_config_inst_regs_1_sva_dfm_5[3:2]), (act_config_inst_regs_2_sva_dfm_5[3:2]),
          (act_config_inst_regs_3_sva_dfm_5[3:2]), (act_config_inst_regs_4_sva_dfm_5[3:2]),
          (act_config_inst_regs_5_sva_dfm_5[3:2]), (act_config_inst_regs_6_sva_dfm_5[3:2]),
          (act_config_inst_regs_7_sva_dfm_5[3:2]), (act_config_inst_regs_8_sva_dfm_5[3:2]),
          (act_config_inst_regs_9_sva_dfm_5[3:2]), (act_config_inst_regs_10_sva_dfm_5[3:2]),
          (act_config_inst_regs_11_sva_dfm_5[3:2]), (act_config_inst_regs_12_sva_dfm_5[3:2]),
          (act_config_inst_regs_13_sva_dfm_5[3:2]), (act_config_inst_regs_14_sva_dfm_5[3:2]),
          (act_config_inst_regs_15_sva_dfm_5[3:2]), ActUnit_DecodeAxiWrite_if_mux_5_nl,
          ActUnit_DecodeAxiWrite_if_mux_7_nl, ActUnit_DecodeAxiWrite_if_mux_9_nl,
          ActUnit_DecodeAxiWrite_if_mux_11_nl, ActUnit_DecodeAxiWrite_if_mux_13_nl,
          ActUnit_DecodeAxiWrite_if_mux_15_nl, ActUnit_DecodeAxiWrite_if_mux_17_nl,
          ActUnit_DecodeAxiWrite_if_mux_19_nl, ActUnit_DecodeAxiWrite_if_mux_21_nl,
          ActUnit_DecodeAxiWrite_if_mux_23_nl, ActUnit_DecodeAxiWrite_if_mux_25_nl,
          ActUnit_DecodeAxiWrite_if_mux_27_nl, ActUnit_DecodeAxiWrite_if_mux_29_nl,
          ActUnit_DecodeAxiWrite_if_mux_31_nl, ActUnit_DecodeAxiWrite_if_mux_33_nl,
          ActUnit_DecodeAxiWrite_if_mux_35_nl, act_config_inst_counter_sva);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_15_sva_8_31 <= 1'b0;
      act_regs_data_3_15_sva_8_30_0 <= 31'b0000000000000000000000000000000;
      act_regs_data_3_14_sva_8_31 <= 1'b0;
      act_regs_data_3_14_sva_8_30_0 <= 31'b0000000000000000000000000000000;
      act_regs_data_3_13_sva_8_31 <= 1'b0;
      act_regs_data_3_13_sva_8_30_0 <= 31'b0000000000000000000000000000000;
      act_regs_data_3_12_sva_8_31 <= 1'b0;
      act_regs_data_3_12_sva_8_30_0 <= 31'b0000000000000000000000000000000;
      act_regs_data_3_11_sva_8_31 <= 1'b0;
      act_regs_data_3_11_sva_8_30_0 <= 31'b0000000000000000000000000000000;
      act_regs_data_3_10_sva_8_31 <= 1'b0;
      act_regs_data_3_10_sva_8_30_0 <= 31'b0000000000000000000000000000000;
      act_regs_data_3_9_sva_8_31 <= 1'b0;
      act_regs_data_3_9_sva_8_30_0 <= 31'b0000000000000000000000000000000;
      act_regs_data_3_8_sva_8_31 <= 1'b0;
      act_regs_data_3_8_sva_8_30_0 <= 31'b0000000000000000000000000000000;
      act_regs_data_3_7_sva_8_31 <= 1'b0;
      act_regs_data_3_7_sva_8_30_0 <= 31'b0000000000000000000000000000000;
      act_regs_data_3_6_sva_8_31 <= 1'b0;
      act_regs_data_3_6_sva_8_30_0 <= 31'b0000000000000000000000000000000;
      act_regs_data_3_5_sva_8_31 <= 1'b0;
      act_regs_data_3_5_sva_8_30_0 <= 31'b0000000000000000000000000000000;
      act_regs_data_3_4_sva_8_31 <= 1'b0;
      act_regs_data_3_4_sva_8_30_0 <= 31'b0000000000000000000000000000000;
      act_regs_data_3_3_sva_8_31 <= 1'b0;
      act_regs_data_3_3_sva_8_30_0 <= 31'b0000000000000000000000000000000;
      act_regs_data_3_2_sva_8_31 <= 1'b0;
      act_regs_data_3_2_sva_8_30_0 <= 31'b0000000000000000000000000000000;
      act_regs_data_3_1_sva_8_31 <= 1'b0;
      act_regs_data_3_1_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_284_cse ) begin
      act_regs_data_3_15_sva_8_31 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_3_15_sva_dfm_2_31, or_832_ssc);
      act_regs_data_3_15_sva_8_30_0 <= MUX_v_31_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_3_15_sva_dfm_2_30_0, or_832_ssc);
      act_regs_data_3_14_sva_8_31 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_3_14_sva_dfm_2_31, or_833_ssc);
      act_regs_data_3_14_sva_8_30_0 <= MUX_v_31_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_3_14_sva_dfm_2_30_0, or_833_ssc);
      act_regs_data_3_13_sva_8_31 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_3_13_sva_dfm_2_31, or_836_ssc);
      act_regs_data_3_13_sva_8_30_0 <= MUX_v_31_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_3_13_sva_dfm_2_30_0, or_836_ssc);
      act_regs_data_3_12_sva_8_31 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_3_12_sva_dfm_2_31, or_837_ssc);
      act_regs_data_3_12_sva_8_30_0 <= MUX_v_31_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_3_12_sva_dfm_2_30_0, or_837_ssc);
      act_regs_data_3_11_sva_8_31 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_3_11_sva_dfm_2_31, or_838_ssc);
      act_regs_data_3_11_sva_8_30_0 <= MUX_v_31_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_3_11_sva_dfm_2_30_0, or_838_ssc);
      act_regs_data_3_10_sva_8_31 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_3_10_sva_dfm_2_31, or_839_ssc);
      act_regs_data_3_10_sva_8_30_0 <= MUX_v_31_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_3_10_sva_dfm_2_30_0, or_839_ssc);
      act_regs_data_3_9_sva_8_31 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_3_9_sva_dfm_2_31, or_840_ssc);
      act_regs_data_3_9_sva_8_30_0 <= MUX_v_31_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_3_9_sva_dfm_2_30_0, or_840_ssc);
      act_regs_data_3_8_sva_8_31 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_3_8_sva_dfm_2_31, or_841_ssc);
      act_regs_data_3_8_sva_8_30_0 <= MUX_v_31_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_3_8_sva_dfm_2_30_0, or_841_ssc);
      act_regs_data_3_7_sva_8_31 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_3_7_sva_dfm_2_31, or_842_ssc);
      act_regs_data_3_7_sva_8_30_0 <= MUX_v_31_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_3_7_sva_dfm_2_30_0, or_842_ssc);
      act_regs_data_3_6_sva_8_31 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_3_6_sva_dfm_2_31, or_843_ssc);
      act_regs_data_3_6_sva_8_30_0 <= MUX_v_31_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_3_6_sva_dfm_2_30_0, or_843_ssc);
      act_regs_data_3_5_sva_8_31 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_3_5_sva_dfm_2_31, or_844_ssc);
      act_regs_data_3_5_sva_8_30_0 <= MUX_v_31_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_3_5_sva_dfm_2_30_0, or_844_ssc);
      act_regs_data_3_4_sva_8_31 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_3_4_sva_dfm_2_31, or_845_ssc);
      act_regs_data_3_4_sva_8_30_0 <= MUX_v_31_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_3_4_sva_dfm_2_30_0, or_845_ssc);
      act_regs_data_3_3_sva_8_31 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_3_3_sva_dfm_2_31, or_846_ssc);
      act_regs_data_3_3_sva_8_30_0 <= MUX_v_31_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_3_3_sva_dfm_2_30_0, or_846_ssc);
      act_regs_data_3_2_sva_8_31 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_3_2_sva_dfm_2_31, or_847_ssc);
      act_regs_data_3_2_sva_8_30_0 <= MUX_v_31_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_3_2_sva_dfm_2_30_0, or_847_ssc);
      act_regs_data_3_1_sva_8_31 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_3_1_sva_dfm_2_31, or_848_ssc);
      act_regs_data_3_1_sva_8_30_0 <= MUX_v_31_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_3_1_sva_dfm_2_30_0, or_848_ssc);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_0_sva_8_31 <= 1'b0;
      act_regs_data_3_0_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_94_ssc ) begin
      act_regs_data_3_0_sva_8_31 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_69_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_3_0_sva_dfm_2_31, {(~ and_dcpl_849) , act_regs_data_and_434_ssc
          , act_regs_data_and_435_ssc});
      act_regs_data_3_0_sva_8_30_0 <= MUX1HOT_v_31_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_174_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_3_0_sva_dfm_2_30_0, {(~ and_dcpl_849) , act_regs_data_and_434_ssc
          , act_regs_data_and_435_ssc});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_15_sva_8_31 <= 1'b0;
      act_regs_data_2_15_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_95_ssc ) begin
      act_regs_data_2_15_sva_8_31 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_104_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_2_15_sva_dfm_2_31, {(~ and_dcpl_849) , act_regs_data_and_436_ssc
          , act_regs_data_and_437_ssc});
      act_regs_data_2_15_sva_8_30_0 <= MUX1HOT_v_31_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_173_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_2_15_sva_dfm_2_30_0, {(~ and_dcpl_849) , act_regs_data_and_436_ssc
          , act_regs_data_and_437_ssc});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_14_sva_8_31 <= 1'b0;
      act_regs_data_2_14_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_96_ssc ) begin
      act_regs_data_2_14_sva_8_31 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_97_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_2_14_sva_dfm_2_31, {(~ and_dcpl_849) , act_regs_data_and_438_ssc
          , act_regs_data_and_439_ssc});
      act_regs_data_2_14_sva_8_30_0 <= MUX1HOT_v_31_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_171_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_2_14_sva_dfm_2_30_0, {(~ and_dcpl_849) , act_regs_data_and_438_ssc
          , act_regs_data_and_439_ssc});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_13_sva_8_31 <= 1'b0;
      act_regs_data_2_13_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_97_ssc ) begin
      act_regs_data_2_13_sva_8_31 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_90_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_2_13_sva_dfm_2_31, {(~ and_dcpl_849) , act_regs_data_and_440_ssc
          , act_regs_data_and_441_ssc});
      act_regs_data_2_13_sva_8_30_0 <= MUX1HOT_v_31_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_169_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_2_13_sva_dfm_2_30_0, {(~ and_dcpl_849) , act_regs_data_and_440_ssc
          , act_regs_data_and_441_ssc});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_12_sva_8_31 <= 1'b0;
      act_regs_data_2_12_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_98_ssc ) begin
      act_regs_data_2_12_sva_8_31 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_83_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_2_12_sva_dfm_2_31, {(~ and_dcpl_849) , act_regs_data_and_442_ssc
          , act_regs_data_and_443_ssc});
      act_regs_data_2_12_sva_8_30_0 <= MUX1HOT_v_31_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_167_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_2_12_sva_dfm_2_30_0, {(~ and_dcpl_849) , act_regs_data_and_442_ssc
          , act_regs_data_and_443_ssc});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_11_sva_8_31 <= 1'b0;
      act_regs_data_2_11_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_99_ssc ) begin
      act_regs_data_2_11_sva_8_31 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_76_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_2_11_sva_dfm_2_31, {(~ and_dcpl_849) , act_regs_data_and_444_ssc
          , act_regs_data_and_445_ssc});
      act_regs_data_2_11_sva_8_30_0 <= MUX1HOT_v_31_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_165_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_2_11_sva_dfm_2_30_0, {(~ and_dcpl_849) , act_regs_data_and_444_ssc
          , act_regs_data_and_445_ssc});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_10_sva_8_31 <= 1'b0;
      act_regs_data_2_10_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_100_ssc ) begin
      act_regs_data_2_10_sva_8_31 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_12_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_2_10_sva_dfm_2_31, {(~ and_dcpl_849) , act_regs_data_and_446_ssc
          , act_regs_data_and_447_ssc});
      act_regs_data_2_10_sva_8_30_0 <= MUX1HOT_v_31_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_163_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_2_10_sva_dfm_2_30_0, {(~ and_dcpl_849) , act_regs_data_and_446_ssc
          , act_regs_data_and_447_ssc});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_9_sva_8_31 <= 1'b0;
      act_regs_data_2_9_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_101_ssc ) begin
      act_regs_data_2_9_sva_8_31 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_62_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_2_9_sva_dfm_2_31, {(~ and_dcpl_849) , act_regs_data_and_448_ssc
          , act_regs_data_and_449_ssc});
      act_regs_data_2_9_sva_8_30_0 <= MUX1HOT_v_31_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_161_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_2_9_sva_dfm_2_30_0, {(~ and_dcpl_849) , act_regs_data_and_448_ssc
          , act_regs_data_and_449_ssc});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_8_sva_8_31 <= 1'b0;
      act_regs_data_2_8_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_102_ssc ) begin
      act_regs_data_2_8_sva_8_31 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_54_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_2_8_sva_dfm_2_31, {(~ and_dcpl_849) , act_regs_data_and_450_ssc
          , act_regs_data_and_451_ssc});
      act_regs_data_2_8_sva_8_30_0 <= MUX1HOT_v_31_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_159_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_2_8_sva_dfm_2_30_0, {(~ and_dcpl_849) , act_regs_data_and_450_ssc
          , act_regs_data_and_451_ssc});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_7_sva_8_31 <= 1'b0;
      act_regs_data_2_7_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_103_ssc ) begin
      act_regs_data_2_7_sva_8_31 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_47_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_2_7_sva_dfm_2_31, {(~ and_dcpl_849) , act_regs_data_and_452_ssc
          , act_regs_data_and_453_ssc});
      act_regs_data_2_7_sva_8_30_0 <= MUX1HOT_v_31_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_157_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_2_7_sva_dfm_2_30_0, {(~ and_dcpl_849) , act_regs_data_and_452_ssc
          , act_regs_data_and_453_ssc});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_6_sva_8_31 <= 1'b0;
      act_regs_data_2_6_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_104_ssc ) begin
      act_regs_data_2_6_sva_8_31 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_40_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_2_6_sva_dfm_2_31, {(~ and_dcpl_849) , act_regs_data_and_454_ssc
          , act_regs_data_and_455_ssc});
      act_regs_data_2_6_sva_8_30_0 <= MUX1HOT_v_31_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_155_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_2_6_sva_dfm_2_30_0, {(~ and_dcpl_849) , act_regs_data_and_454_ssc
          , act_regs_data_and_455_ssc});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_5_sva_8_31 <= 1'b0;
      act_regs_data_2_5_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_105_ssc ) begin
      act_regs_data_2_5_sva_8_31 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_33_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_2_5_sva_dfm_2_31, {(~ and_dcpl_849) , act_regs_data_and_456_ssc
          , act_regs_data_and_457_ssc});
      act_regs_data_2_5_sva_8_30_0 <= MUX1HOT_v_31_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_153_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_2_5_sva_dfm_2_30_0, {(~ and_dcpl_849) , act_regs_data_and_456_ssc
          , act_regs_data_and_457_ssc});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_4_sva_8_31 <= 1'b0;
      act_regs_data_2_4_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_106_ssc ) begin
      act_regs_data_2_4_sva_8_31 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_26_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_2_4_sva_dfm_2_31, {(~ and_dcpl_849) , act_regs_data_and_458_ssc
          , act_regs_data_and_459_ssc});
      act_regs_data_2_4_sva_8_30_0 <= MUX1HOT_v_31_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_151_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_2_4_sva_dfm_2_30_0, {(~ and_dcpl_849) , act_regs_data_and_458_ssc
          , act_regs_data_and_459_ssc});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_3_sva_8_31 <= 1'b0;
      act_regs_data_2_3_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_107_ssc ) begin
      act_regs_data_2_3_sva_8_31 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_19_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_2_3_sva_dfm_2_31, {(~ and_dcpl_849) , act_regs_data_and_460_ssc
          , act_regs_data_and_461_ssc});
      act_regs_data_2_3_sva_8_30_0 <= MUX1HOT_v_31_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_149_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_2_3_sva_dfm_2_30_0, {(~ and_dcpl_849) , act_regs_data_and_460_ssc
          , act_regs_data_and_461_ssc});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_2_sva_8_31 <= 1'b0;
      act_regs_data_2_2_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_108_ssc ) begin
      act_regs_data_2_2_sva_8_31 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_111_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_2_2_sva_dfm_2_31, {(~ and_dcpl_849) , act_regs_data_and_462_ssc
          , act_regs_data_and_463_ssc});
      act_regs_data_2_2_sva_8_30_0 <= MUX1HOT_v_31_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_147_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_2_2_sva_dfm_2_30_0, {(~ and_dcpl_849) , act_regs_data_and_462_ssc
          , act_regs_data_and_463_ssc});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_1_sva_8_31 <= 1'b0;
      act_regs_data_2_1_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_109_ssc ) begin
      act_regs_data_2_1_sva_8_31 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_5_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_2_1_sva_dfm_2_31, {(~ and_dcpl_849) , act_regs_data_and_464_ssc
          , act_regs_data_and_465_ssc});
      act_regs_data_2_1_sva_8_30_0 <= MUX1HOT_v_31_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_145_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_2_1_sva_dfm_2_30_0, {(~ and_dcpl_849) , act_regs_data_and_464_ssc
          , act_regs_data_and_465_ssc});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_0_sva_8_31 <= 1'b0;
      act_regs_data_2_0_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_110_ssc ) begin
      act_regs_data_2_0_sva_8_31 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_67_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_2_0_sva_dfm_2_31, {(~ and_dcpl_849) , act_regs_data_and_466_ssc
          , act_regs_data_and_467_ssc});
      act_regs_data_2_0_sva_8_30_0 <= MUX1HOT_v_31_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_143_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_2_0_sva_dfm_2_30_0, {(~ and_dcpl_849) , act_regs_data_and_466_ssc
          , act_regs_data_and_467_ssc});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_15_sva_8_31 <= 1'b0;
      act_regs_data_1_15_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_111_ssc ) begin
      act_regs_data_1_15_sva_8_31 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_102_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_1_15_sva_dfm_2_31, {(~ and_dcpl_849) , act_regs_data_and_468_ssc
          , act_regs_data_and_469_ssc});
      act_regs_data_1_15_sva_8_30_0 <= MUX1HOT_v_31_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_142_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_1_15_sva_dfm_2_30_0, {(~ and_dcpl_849) , act_regs_data_and_468_ssc
          , act_regs_data_and_469_ssc});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_14_sva_8_31 <= 1'b0;
      act_regs_data_1_14_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_112_ssc ) begin
      act_regs_data_1_14_sva_8_31 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_95_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_1_14_sva_dfm_2_31, {(~ and_dcpl_849) , act_regs_data_and_470_ssc
          , act_regs_data_and_471_ssc});
      act_regs_data_1_14_sva_8_30_0 <= MUX1HOT_v_31_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_144_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_1_14_sva_dfm_2_30_0, {(~ and_dcpl_849) , act_regs_data_and_470_ssc
          , act_regs_data_and_471_ssc});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_13_sva_8_31 <= 1'b0;
      act_regs_data_1_13_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_113_ssc ) begin
      act_regs_data_1_13_sva_8_31 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_88_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_1_13_sva_dfm_2_31, {(~ and_dcpl_849) , act_regs_data_and_472_ssc
          , act_regs_data_and_473_ssc});
      act_regs_data_1_13_sva_8_30_0 <= MUX1HOT_v_31_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_146_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_1_13_sva_dfm_2_30_0, {(~ and_dcpl_849) , act_regs_data_and_472_ssc
          , act_regs_data_and_473_ssc});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_12_sva_8_31 <= 1'b0;
      act_regs_data_1_12_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_114_ssc ) begin
      act_regs_data_1_12_sva_8_31 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_81_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_1_12_sva_dfm_2_31, {(~ and_dcpl_849) , act_regs_data_and_474_ssc
          , act_regs_data_and_475_ssc});
      act_regs_data_1_12_sva_8_30_0 <= MUX1HOT_v_31_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_148_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_1_12_sva_dfm_2_30_0, {(~ and_dcpl_849) , act_regs_data_and_474_ssc
          , act_regs_data_and_475_ssc});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_11_sva_8_31 <= 1'b0;
      act_regs_data_1_11_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_115_ssc ) begin
      act_regs_data_1_11_sva_8_31 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_74_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_1_11_sva_dfm_2_31, {(~ and_dcpl_849) , act_regs_data_and_476_ssc
          , act_regs_data_and_477_ssc});
      act_regs_data_1_11_sva_8_30_0 <= MUX1HOT_v_31_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_150_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_1_11_sva_dfm_2_30_0, {(~ and_dcpl_849) , act_regs_data_and_476_ssc
          , act_regs_data_and_477_ssc});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_10_sva_8_31 <= 1'b0;
      act_regs_data_1_10_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_116_ssc ) begin
      act_regs_data_1_10_sva_8_31 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_10_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_1_10_sva_dfm_2_31, {(~ and_dcpl_849) , act_regs_data_and_478_ssc
          , act_regs_data_and_479_ssc});
      act_regs_data_1_10_sva_8_30_0 <= MUX1HOT_v_31_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_152_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_1_10_sva_dfm_2_30_0, {(~ and_dcpl_849) , act_regs_data_and_478_ssc
          , act_regs_data_and_479_ssc});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_9_sva_8_31 <= 1'b0;
      act_regs_data_1_9_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_117_ssc ) begin
      act_regs_data_1_9_sva_8_31 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_60_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_1_9_sva_dfm_2_31, {(~ and_dcpl_849) , act_regs_data_and_480_ssc
          , act_regs_data_and_481_ssc});
      act_regs_data_1_9_sva_8_30_0 <= MUX1HOT_v_31_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_154_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_1_9_sva_dfm_2_30_0, {(~ and_dcpl_849) , act_regs_data_and_480_ssc
          , act_regs_data_and_481_ssc});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_8_sva_8_31 <= 1'b0;
      act_regs_data_1_8_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_118_ssc ) begin
      act_regs_data_1_8_sva_8_31 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_52_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_1_8_sva_dfm_2_31, {(~ and_dcpl_849) , act_regs_data_and_482_ssc
          , act_regs_data_and_483_ssc});
      act_regs_data_1_8_sva_8_30_0 <= MUX1HOT_v_31_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_156_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_1_8_sva_dfm_2_30_0, {(~ and_dcpl_849) , act_regs_data_and_482_ssc
          , act_regs_data_and_483_ssc});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_7_sva_8_31 <= 1'b0;
      act_regs_data_1_7_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_119_ssc ) begin
      act_regs_data_1_7_sva_8_31 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_45_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_1_7_sva_dfm_2_31, {(~ and_dcpl_849) , act_regs_data_and_484_ssc
          , act_regs_data_and_485_ssc});
      act_regs_data_1_7_sva_8_30_0 <= MUX1HOT_v_31_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_158_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_1_7_sva_dfm_2_30_0, {(~ and_dcpl_849) , act_regs_data_and_484_ssc
          , act_regs_data_and_485_ssc});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_6_sva_8_31 <= 1'b0;
      act_regs_data_1_6_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_120_ssc ) begin
      act_regs_data_1_6_sva_8_31 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_38_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_1_6_sva_dfm_2_31, {(~ and_dcpl_849) , act_regs_data_and_486_ssc
          , act_regs_data_and_487_ssc});
      act_regs_data_1_6_sva_8_30_0 <= MUX1HOT_v_31_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_160_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_1_6_sva_dfm_2_30_0, {(~ and_dcpl_849) , act_regs_data_and_486_ssc
          , act_regs_data_and_487_ssc});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_5_sva_8_31 <= 1'b0;
      act_regs_data_1_5_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_121_ssc ) begin
      act_regs_data_1_5_sva_8_31 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_31_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_1_5_sva_dfm_2_31, {(~ and_dcpl_849) , act_regs_data_and_488_ssc
          , act_regs_data_and_489_ssc});
      act_regs_data_1_5_sva_8_30_0 <= MUX1HOT_v_31_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_162_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_1_5_sva_dfm_2_30_0, {(~ and_dcpl_849) , act_regs_data_and_488_ssc
          , act_regs_data_and_489_ssc});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_4_sva_8_31 <= 1'b0;
      act_regs_data_1_4_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_122_ssc ) begin
      act_regs_data_1_4_sva_8_31 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_24_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_1_4_sva_dfm_2_31, {(~ and_dcpl_849) , act_regs_data_and_490_ssc
          , act_regs_data_and_491_ssc});
      act_regs_data_1_4_sva_8_30_0 <= MUX1HOT_v_31_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_164_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_1_4_sva_dfm_2_30_0, {(~ and_dcpl_849) , act_regs_data_and_490_ssc
          , act_regs_data_and_491_ssc});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_3_sva_8_31 <= 1'b0;
      act_regs_data_1_3_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_123_ssc ) begin
      act_regs_data_1_3_sva_8_31 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_17_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_1_3_sva_dfm_2_31, {(~ and_dcpl_849) , act_regs_data_and_492_ssc
          , act_regs_data_and_493_ssc});
      act_regs_data_1_3_sva_8_30_0 <= MUX1HOT_v_31_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_166_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_1_3_sva_dfm_2_30_0, {(~ and_dcpl_849) , act_regs_data_and_492_ssc
          , act_regs_data_and_493_ssc});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_2_sva_8_31 <= 1'b0;
      act_regs_data_1_2_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_124_ssc ) begin
      act_regs_data_1_2_sva_8_31 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_109_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_1_2_sva_dfm_2_31, {(~ and_dcpl_849) , act_regs_data_and_494_ssc
          , act_regs_data_and_495_ssc});
      act_regs_data_1_2_sva_8_30_0 <= MUX1HOT_v_31_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_168_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_1_2_sva_dfm_2_30_0, {(~ and_dcpl_849) , act_regs_data_and_494_ssc
          , act_regs_data_and_495_ssc});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_1_sva_8_31 <= 1'b0;
      act_regs_data_1_1_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_125_ssc ) begin
      act_regs_data_1_1_sva_8_31 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_3_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_1_1_sva_dfm_2_31, {(~ and_dcpl_849) , act_regs_data_and_496_ssc
          , act_regs_data_and_497_ssc});
      act_regs_data_1_1_sva_8_30_0 <= MUX1HOT_v_31_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_170_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_1_1_sva_dfm_2_30_0, {(~ and_dcpl_849) , act_regs_data_and_496_ssc
          , act_regs_data_and_497_ssc});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_0_sva_8_31 <= 1'b0;
      act_regs_data_1_0_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_126_ssc ) begin
      act_regs_data_1_0_sva_8_31 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_66_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_1_0_sva_dfm_2_31, {(~ and_dcpl_849) , act_regs_data_and_498_ssc
          , act_regs_data_and_499_ssc});
      act_regs_data_1_0_sva_8_30_0 <= MUX1HOT_v_31_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_172_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_1_0_sva_dfm_2_30_0, {(~ and_dcpl_849) , act_regs_data_and_498_ssc
          , act_regs_data_and_499_ssc});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_9_sva_8_31 <= 1'b0;
      act_regs_data_0_9_sva_8_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( act_regs_data_and_127_ssc ) begin
      act_regs_data_0_9_sva_8_31 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_59_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_0_9_sva_dfm_2_31, {(~ and_dcpl_849) , act_regs_data_and_500_ssc
          , act_regs_data_and_501_ssc});
      act_regs_data_0_9_sva_8_30_0 <= MUX1HOT_v_31_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_175_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          act_regs_data_0_9_sva_dfm_2_30_0, {(~ and_dcpl_849) , act_regs_data_and_500_ssc
          , act_regs_data_and_501_ssc});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_CheckStart_start_reg_sva <= 1'b0;
    end
    else if ( ActUnit_CheckStart_start_reg_and_tmp ) begin
      ActUnit_CheckStart_start_reg_sva <= MUX1HOT_s_1_4_2(ActUnit_RunInst_switch_lp_and_32_tmp,
          ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_23_nl, start_PopNB_mioi_data_rsc_z_mxwt,
          while_and_64_nl, {and_dcpl_909 , and_dcpl_829 , and_dcpl_613 , and_dcpl_814});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_y_2_lpi_1_dfm_1_31 <= 1'b0;
      Silu_for_y_2_lpi_1_dfm_1_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( Silu_for_y_and_ssc ) begin
      Silu_for_y_2_lpi_1_dfm_1_31 <= (z_out_3_29_1[28]) & (~ Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
          & (~ Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs);
      Silu_for_y_2_lpi_1_dfm_1_30_0 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          Silu_for_else_mux_1_nl, operator_32_8_true_AC_TRN_AC_WRAP_2_not_34_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & (((~ or_dcpl_495) & mux_223_nl) | and_dcpl_592 | and_dcpl_997
        | and_dcpl_852) ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_31 <= ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_10_nl
          & (~ and_dcpl_997);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1228_tmp ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_30_0 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_83_nl, nor_772_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_y_4_lpi_1_dfm_1_31 <= 1'b0;
      Silu_for_y_4_lpi_1_dfm_1_30_0 <= 31'b0000000000000000000000000000000;
      Silu_for_y_3_lpi_1_dfm_1_31 <= 1'b0;
      Silu_for_y_3_lpi_1_dfm_1_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( Silu_for_y_and_13_ssc ) begin
      Silu_for_y_4_lpi_1_dfm_1_31 <= (z_out_4_29_1[28]) & (~ Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
          & (~ Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs);
      Silu_for_y_4_lpi_1_dfm_1_30_0 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          Silu_for_else_mux_3_nl, operator_32_8_true_AC_TRN_AC_WRAP_2_not_36_nl);
      Silu_for_y_3_lpi_1_dfm_1_31 <= (z_out_3_29_1[28]) & (~ Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
          & (~ Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs);
      Silu_for_y_3_lpi_1_dfm_1_30_0 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          Silu_for_else_mux_2_nl, operator_32_8_true_AC_TRN_AC_WRAP_2_not_35_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_else_else_slc_Tanh_for_1_else_else_mul_1_cmp_z_46_0_itm <= 47'b00000000000000000000000000000000000000000000000;
    end
    else if ( ActUnitRun_wen & (~ and_dcpl_614) & and_dcpl_162 & (act_config_in_InstFetch_return_sva_7_2[2])
        & (~ Gelu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs)
        & (~ Gelu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
        ) begin
      Gelu_for_else_else_slc_Tanh_for_1_else_else_mul_1_cmp_z_46_0_itm <= Tanh_for_1_else_else_mul_1_cmp_z[46:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_y_6_lpi_1_dfm_1_31 <= 1'b0;
      Silu_for_y_6_lpi_1_dfm_1_30_0 <= 31'b0000000000000000000000000000000;
      Silu_for_y_5_lpi_1_dfm_1_31 <= 1'b0;
      Silu_for_y_5_lpi_1_dfm_1_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( Silu_for_y_and_15_ssc ) begin
      Silu_for_y_6_lpi_1_dfm_1_31 <= (z_out_4_29_1[28]) & (~ Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
          & (~ Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs);
      Silu_for_y_6_lpi_1_dfm_1_30_0 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          Silu_for_else_mux_5_nl, operator_32_8_true_AC_TRN_AC_WRAP_2_not_38_nl);
      Silu_for_y_5_lpi_1_dfm_1_31 <= (z_out_3_29_1[28]) & (~ Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
          & (~ Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs);
      Silu_for_y_5_lpi_1_dfm_1_30_0 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          Silu_for_else_mux_4_nl, operator_32_8_true_AC_TRN_AC_WRAP_2_not_37_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_else_else_slc_Tanh_for_1_else_else_mul_cmp_15_z_46_0_itm <= 47'b00000000000000000000000000000000000000000000000;
    end
    else if ( Gelu_for_else_else_and_1_cse & and_dcpl_162 & (act_config_in_InstFetch_return_sva_7_2[2])
        & (~ Gelu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
        & (~ Gelu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs)
        ) begin
      Gelu_for_else_else_slc_Tanh_for_1_else_else_mul_cmp_15_z_46_0_itm <= Tanh_for_1_else_else_mul_cmp_15_z[46:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_else_else_slc_Tanh_for_1_else_else_mul_cmp_z_46_0_itm <= 47'b00000000000000000000000000000000000000000000000;
    end
    else if ( Gelu_for_else_else_and_1_cse & and_dcpl_162 & (act_config_in_InstFetch_return_sva_7_2[2])
        & (~ Gelu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs)
        & (~ Gelu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
        ) begin
      Gelu_for_else_else_slc_Tanh_for_1_else_else_mul_cmp_z_46_0_itm <= Tanh_for_1_else_else_mul_cmp_z[46:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_else_else_slc_Tanh_for_1_else_else_mul_cmp_12_z_46_0_itm <= 47'b00000000000000000000000000000000000000000000000;
    end
    else if ( Gelu_for_else_else_and_1_cse & and_dcpl_162 & (act_config_in_InstFetch_return_sva_7_2[2])
        & (~ Gelu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs)
        & (~ Gelu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
        ) begin
      Gelu_for_else_else_slc_Tanh_for_1_else_else_mul_cmp_12_z_46_0_itm <= Tanh_for_1_else_else_mul_cmp_12_z[46:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_else_else_slc_Tanh_for_1_else_else_mul_cmp_13_z_46_0_itm <= 47'b00000000000000000000000000000000000000000000000;
    end
    else if ( ActUnitRun_wen & (mux_227_nl | (fsm_output[4])) & and_dcpl_162 & (act_config_in_InstFetch_return_sva_7_2[2])
        & (~ Tanh_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs)
        & (~ Tanh_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)
        ) begin
      Gelu_for_else_else_slc_Tanh_for_1_else_else_mul_cmp_13_z_46_0_itm <= Tanh_for_1_else_else_mul_cmp_13_z[46:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_y_8_lpi_1_dfm_1_31 <= 1'b0;
      Silu_for_y_8_lpi_1_dfm_1_30_0 <= 31'b0000000000000000000000000000000;
      Silu_for_y_7_lpi_1_dfm_1_31 <= 1'b0;
      Silu_for_y_7_lpi_1_dfm_1_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( Silu_for_y_and_17_ssc ) begin
      Silu_for_y_8_lpi_1_dfm_1_31 <= (z_out_3_29_1[28]) & (~ Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
          & (~ Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs);
      Silu_for_y_8_lpi_1_dfm_1_30_0 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          Silu_for_else_mux_7_nl, operator_32_8_true_AC_TRN_AC_WRAP_2_not_40_nl);
      Silu_for_y_7_lpi_1_dfm_1_31 <= (z_out_4_29_1[28]) & (~ Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
          & (~ Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs);
      Silu_for_y_7_lpi_1_dfm_1_30_0 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          Silu_for_else_mux_6_nl, operator_32_8_true_AC_TRN_AC_WRAP_2_not_39_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_y_9_lpi_1_dfm_1_31 <= 1'b0;
      Silu_for_y_9_lpi_1_dfm_1_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( Silu_for_y_and_19_ssc ) begin
      Silu_for_y_9_lpi_1_dfm_1_31 <= (z_out_4_29_1[28]) & (~ Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
          & (~ Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs);
      Silu_for_y_9_lpi_1_dfm_1_30_0 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          Silu_for_else_mux_8_nl, operator_32_8_true_AC_TRN_AC_WRAP_2_not_41_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_474 | (~ mux_229_itm))) | and_dcpl_576
        | and_dcpl_997 | and_dcpl_852) ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_31 <= ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_15_nl
          & (~ and_dcpl_997);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1231_tmp ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_30_0 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_78_nl, nor_773_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_497 | (~ mux_229_itm))) | and_dcpl_576
        | and_dcpl_997 | and_dcpl_852) ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_31 <= ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_20_nl
          & (~ and_dcpl_997);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1234_tmp ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_30_0 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_82_nl, nor_774_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_31 <= 1'b0;
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( Silu_for_y_and_7_cse ) begin
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_31 <= MUX_s_1_2_2(Gelu_for_Gelu_for_and_nl,
          ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_2_31, and_dcpl_832);
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_30_0 <= MUX_v_31_2_2(Gelu_for_Gelu_for_and_19_nl,
          ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_2_30_0, and_dcpl_832);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_y_12_lpi_1_dfm_1_31 <= 1'b0;
      Silu_for_y_12_lpi_1_dfm_1_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( Silu_for_y_and_8_ssc ) begin
      Silu_for_y_12_lpi_1_dfm_1_31 <= (z_out_3_29_1[28]) & (~ Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
          & (~ Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs);
      Silu_for_y_12_lpi_1_dfm_1_30_0 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          Silu_for_else_mux_11_nl, operator_32_8_true_AC_TRN_AC_WRAP_2_not_42_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_477 | (~ mux_231_itm))) | and_dcpl_578
        | and_dcpl_997 | and_dcpl_852) ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_31 <= ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_25_nl
          & (~ and_dcpl_997);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1237_tmp ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_30_0 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_77_nl, nor_775_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_499 | (~ mux_231_itm))) | and_dcpl_578
        | and_dcpl_997 | and_dcpl_852) ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_31 <= ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_30_nl
          & (~ and_dcpl_997);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1240_tmp ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_30_0 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_81_nl, nor_776_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_y_14_lpi_1_dfm_1_31 <= 1'b0;
      Silu_for_y_14_lpi_1_dfm_1_30_0 <= 31'b0000000000000000000000000000000;
      Silu_for_y_13_lpi_1_dfm_1_31 <= 1'b0;
      Silu_for_y_13_lpi_1_dfm_1_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( Silu_for_y_and_20_ssc ) begin
      Silu_for_y_14_lpi_1_dfm_1_31 <= (z_out_3_29_1[28]) & (~ Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
          & (~ Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs);
      Silu_for_y_14_lpi_1_dfm_1_30_0 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          Silu_for_else_mux_13_nl, operator_32_8_true_AC_TRN_AC_WRAP_2_not_44_nl);
      Silu_for_y_13_lpi_1_dfm_1_31 <= (z_out_4_29_1[28]) & (~ Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
          & (~ Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs);
      Silu_for_y_13_lpi_1_dfm_1_30_0 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          Silu_for_else_mux_12_nl, operator_32_8_true_AC_TRN_AC_WRAP_2_not_43_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_480 | (~ mux_234_itm))) | and_dcpl_1006
        | and_dcpl_997 | and_dcpl_852) ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_31 <= ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_35_nl
          & (~ and_dcpl_997);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1243_tmp ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_30_0 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_76_nl, nor_777_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_482 | (~ mux_234_itm))) | and_dcpl_1006
        | and_dcpl_997 | and_dcpl_852) ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_31 <= ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_40_nl
          & (~ and_dcpl_997);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1246_tmp ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_30_0 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_88_nl, nor_778_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_y_lpi_1_dfm_1_31 <= 1'b0;
      Silu_for_y_lpi_1_dfm_1_30_0 <= 31'b0000000000000000000000000000000;
      Silu_for_y_15_lpi_1_dfm_1_31 <= 1'b0;
      Silu_for_y_15_lpi_1_dfm_1_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( Silu_for_y_and_22_ssc ) begin
      Silu_for_y_lpi_1_dfm_1_31 <= (z_out_3_29_1[28]) & (~ Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
          & (~ Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs);
      Silu_for_y_lpi_1_dfm_1_30_0 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          Silu_for_else_mux_15_nl, operator_32_8_true_AC_TRN_AC_WRAP_2_not_46_nl);
      Silu_for_y_15_lpi_1_dfm_1_31 <= (z_out_4_29_1[28]) & (~ Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
          & (~ Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs);
      Silu_for_y_15_lpi_1_dfm_1_30_0 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          Silu_for_else_mux_14_nl, operator_32_8_true_AC_TRN_AC_WRAP_2_not_45_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_484 | and_dcpl_901)) | and_dcpl_900 |
        and_dcpl_997 | and_dcpl_852) ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_31 <= ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_45_nl
          & (~ and_dcpl_997);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1250_tmp ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_30_0 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_87_nl, nor_779_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_487 | and_dcpl_901)) | and_dcpl_900 |
        and_dcpl_997 | and_dcpl_852) ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_31 <= ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_50_nl
          & (~ and_dcpl_997);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1254_tmp ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_30_0 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_86_nl, nor_780_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_1_sva_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_456 | and_dcpl_799)) | and_dcpl_1007 |
        and_dcpl_997 | and_dcpl_852) ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_1_sva_31 <= ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_55_nl
          & (~ and_dcpl_997);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_1_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1261_tmp ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_1_sva_30_0 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_89_nl, nor_781_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_462 | and_dcpl_799)) | and_dcpl_1007 |
        and_dcpl_997 | and_dcpl_852) ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_31 <= ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_60_nl
          & (~ and_dcpl_997);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1268_tmp ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_30_0 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_80_nl, nor_782_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_469 | and_dcpl_799)) | and_dcpl_1007 |
        and_dcpl_997 | and_dcpl_852) ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_31 <= ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_65_nl
          & (~ and_dcpl_997);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1275_tmp ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_30_0 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_79_nl, nor_783_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_489 | and_dcpl_799)) | and_dcpl_1007 |
        and_dcpl_997 | and_dcpl_852) ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_31 <= ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_70_nl
          & (~ and_dcpl_997);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1282_tmp ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_30_0 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_85_nl, nor_784_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_492 | and_dcpl_799)) | and_dcpl_1007 |
        and_dcpl_997 | and_dcpl_852) ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_31 <= ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_75_nl
          & (~ and_dcpl_997);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1289_tmp ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_30_0 <= MUX_v_31_2_2(31'b0000000000000000000000000000000,
          ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_84_nl, nor_785_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_0_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_563 | or_dcpl_451 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_0_0_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_273_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_0_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1291_tmp ) begin
      act_regs_data_0_0_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_0_0_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[30:0]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_1_exs_5_30_0, Relu_for_y_qr_30_0_1_lpi_1_dfm, ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_30_0,
          ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_299_cse , act_regs_data_and_300_cse , act_regs_data_and_301_cse
          , act_regs_data_and_302_cse , act_regs_data_and_303_cse , act_regs_data_and_304_cse
          , act_regs_data_and_305_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_1_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_563 | or_dcpl_458 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_0_1_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_272_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_1_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1293_tmp ) begin
      act_regs_data_0_1_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_0_1_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[62:32]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_2_exs_5_30_0, Relu_for_y_qr_30_0_2_lpi_1_dfm, Silu_for_y_2_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_299_cse , act_regs_data_and_300_cse , act_regs_data_and_301_cse
          , act_regs_data_and_302_cse , act_regs_data_and_303_cse , act_regs_data_and_304_cse
          , act_regs_data_and_305_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_2_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_567 | or_dcpl_451 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_0_2_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_271_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_2_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1295_tmp ) begin
      act_regs_data_0_2_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_0_2_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[94:64]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_3_exs_5_30_0, Relu_for_y_qr_30_0_3_lpi_1_dfm, Silu_for_y_3_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_299_cse , act_regs_data_and_300_cse , act_regs_data_and_301_cse
          , act_regs_data_and_302_cse , act_regs_data_and_303_cse , act_regs_data_and_304_cse
          , act_regs_data_and_305_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_3_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_567 | or_dcpl_458 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_0_3_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_270_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_3_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1297_tmp ) begin
      act_regs_data_0_3_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_0_3_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[126:96]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_4_exs_5_30_0, Relu_for_y_qr_30_0_4_lpi_1_dfm, Silu_for_y_4_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_299_cse , act_regs_data_and_300_cse , act_regs_data_and_301_cse
          , act_regs_data_and_302_cse , act_regs_data_and_303_cse , act_regs_data_and_304_cse
          , act_regs_data_and_305_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_4_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_563 | or_dcpl_490 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_0_4_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_269_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_4_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1299_tmp ) begin
      act_regs_data_0_4_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_0_4_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[158:128]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_5_exs_5_30_0, Relu_for_y_qr_30_0_5_lpi_1_dfm, Silu_for_y_5_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_299_cse , act_regs_data_and_300_cse , act_regs_data_and_301_cse
          , act_regs_data_and_302_cse , act_regs_data_and_303_cse , act_regs_data_and_304_cse
          , act_regs_data_and_305_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_5_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_563 | or_dcpl_493 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_0_5_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_268_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_5_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1301_tmp ) begin
      act_regs_data_0_5_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_0_5_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[190:160]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_6_exs_5_30_0, Relu_for_y_qr_30_0_6_lpi_1_dfm, Silu_for_y_6_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_299_cse , act_regs_data_and_300_cse , act_regs_data_and_301_cse
          , act_regs_data_and_302_cse , act_regs_data_and_303_cse , act_regs_data_and_304_cse
          , act_regs_data_and_305_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_6_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_567 | or_dcpl_490 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_0_6_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_267_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_6_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1303_tmp ) begin
      act_regs_data_0_6_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_0_6_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[222:192]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_7_exs_5_30_0, Relu_for_y_qr_30_0_7_lpi_1_dfm, Silu_for_y_7_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_299_cse , act_regs_data_and_300_cse , act_regs_data_and_301_cse
          , act_regs_data_and_302_cse , act_regs_data_and_303_cse , act_regs_data_and_304_cse
          , act_regs_data_and_305_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_7_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_567 | or_dcpl_493 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_0_7_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_266_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_7_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1305_tmp ) begin
      act_regs_data_0_7_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_0_7_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[254:224]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_8_exs_5_30_0, Relu_for_y_qr_30_0_8_lpi_1_dfm, Silu_for_y_8_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_299_cse , act_regs_data_and_300_cse , act_regs_data_and_301_cse
          , act_regs_data_and_302_cse , act_regs_data_and_303_cse , act_regs_data_and_304_cse
          , act_regs_data_and_305_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_8_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_563 | or_dcpl_464 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_0_8_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_265_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_8_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1307_tmp ) begin
      act_regs_data_0_8_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_0_8_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[286:256]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_9_exs_5_30_0, Relu_for_y_qr_30_0_9_lpi_1_dfm, Silu_for_y_9_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_299_cse , act_regs_data_and_300_cse , act_regs_data_and_301_cse
          , act_regs_data_and_302_cse , act_regs_data_and_303_cse , act_regs_data_and_304_cse
          , act_regs_data_and_305_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_9_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_563 | or_dcpl_471 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_0_9_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_264_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_9_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1309_tmp ) begin
      act_regs_data_0_9_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_0_9_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[318:288]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_10_exs_5_30_0, Relu_for_y_qr_30_0_10_lpi_1_dfm, ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_30_0,
          Gelu_for_y_10_lpi_1_dfm_2_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_299_cse , act_regs_data_and_300_cse , act_regs_data_and_301_cse
          , act_regs_data_and_302_cse , act_regs_data_and_303_cse , act_regs_data_and_304_cse
          , act_regs_data_and_305_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_10_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_567 | or_dcpl_464 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_0_10_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_263_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_10_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1311_tmp ) begin
      act_regs_data_0_10_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_0_10_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[350:320]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_11_exs_5_30_0, Relu_for_y_qr_30_0_11_lpi_1_dfm, ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_30_0,
          Gelu_for_y_11_lpi_1_dfm_2_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_299_cse , act_regs_data_and_300_cse , act_regs_data_and_301_cse
          , act_regs_data_and_302_cse , act_regs_data_and_303_cse , act_regs_data_and_304_cse
          , act_regs_data_and_305_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_11_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_567 | or_dcpl_471 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_0_11_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_262_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_11_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1313_tmp ) begin
      act_regs_data_0_11_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_0_11_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[382:352]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_12_exs_5_30_0, Relu_for_y_qr_30_0_12_lpi_1_dfm, Silu_for_y_12_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_299_cse , act_regs_data_and_300_cse , act_regs_data_and_301_cse
          , act_regs_data_and_302_cse , act_regs_data_and_303_cse , act_regs_data_and_304_cse
          , act_regs_data_and_305_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_12_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_563 | or_dcpl_475 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_0_12_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_261_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_12_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1315_tmp ) begin
      act_regs_data_0_12_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_0_12_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[414:384]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_13_exs_5_30_0, Relu_for_y_qr_30_0_13_lpi_1_dfm, Silu_for_y_13_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_1_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_299_cse , act_regs_data_and_300_cse , act_regs_data_and_301_cse
          , act_regs_data_and_302_cse , act_regs_data_and_303_cse , act_regs_data_and_304_cse
          , act_regs_data_and_305_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_13_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_563 | or_dcpl_478 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_0_13_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_260_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_13_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1317_tmp ) begin
      act_regs_data_0_13_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_0_13_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[446:416]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_14_exs_5_30_0, Relu_for_y_qr_30_0_14_lpi_1_dfm, Silu_for_y_14_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_299_cse , act_regs_data_and_300_cse , act_regs_data_and_301_cse
          , act_regs_data_and_302_cse , act_regs_data_and_303_cse , act_regs_data_and_304_cse
          , act_regs_data_and_305_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_14_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_567 | or_dcpl_475 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_0_14_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_259_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_14_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1319_tmp ) begin
      act_regs_data_0_14_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_0_14_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[478:448]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_15_exs_5_30_0, Relu_for_y_qr_30_0_15_lpi_1_dfm, Silu_for_y_15_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_299_cse , act_regs_data_and_300_cse , act_regs_data_and_301_cse
          , act_regs_data_and_302_cse , act_regs_data_and_303_cse , act_regs_data_and_304_cse
          , act_regs_data_and_305_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_15_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_567 | or_dcpl_478 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_0_15_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_258_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_15_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1321_tmp ) begin
      act_regs_data_0_15_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_0_15_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[510:480]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_16_exs_5_30_0, Relu_for_y_qr_30_0_lpi_1_dfm, Silu_for_y_lpi_1_dfm_1_30_0,
          Gelu_for_y_lpi_1_dfm_2_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_299_cse , act_regs_data_and_300_cse , act_regs_data_and_301_cse
          , act_regs_data_and_302_cse , act_regs_data_and_303_cse , act_regs_data_and_304_cse
          , act_regs_data_and_305_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_0_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_583 | or_dcpl_451 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_1_0_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_257_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_0_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1323_tmp ) begin
      act_regs_data_1_0_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_1_0_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[30:0]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_1_exs_5_30_0, Relu_for_y_qr_30_0_1_lpi_1_dfm, ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_30_0,
          ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_523_cse , act_regs_data_and_524_cse , act_regs_data_and_525_cse
          , act_regs_data_and_526_cse , act_regs_data_and_527_cse , act_regs_data_and_528_cse
          , act_regs_data_and_529_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_1_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_583 | or_dcpl_458 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_1_1_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_256_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_1_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1325_tmp ) begin
      act_regs_data_1_1_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_1_1_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[62:32]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_2_exs_5_30_0, Relu_for_y_qr_30_0_2_lpi_1_dfm, Silu_for_y_2_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_523_cse , act_regs_data_and_524_cse , act_regs_data_and_525_cse
          , act_regs_data_and_526_cse , act_regs_data_and_527_cse , act_regs_data_and_528_cse
          , act_regs_data_and_529_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_2_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_586 | or_dcpl_451 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_1_2_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_255_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_2_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1327_tmp ) begin
      act_regs_data_1_2_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_1_2_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[94:64]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_3_exs_5_30_0, Relu_for_y_qr_30_0_3_lpi_1_dfm, Silu_for_y_3_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_523_cse , act_regs_data_and_524_cse , act_regs_data_and_525_cse
          , act_regs_data_and_526_cse , act_regs_data_and_527_cse , act_regs_data_and_528_cse
          , act_regs_data_and_529_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_3_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_586 | or_dcpl_458 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_1_3_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_254_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_3_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1329_tmp ) begin
      act_regs_data_1_3_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_1_3_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[126:96]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_4_exs_5_30_0, Relu_for_y_qr_30_0_4_lpi_1_dfm, Silu_for_y_4_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_523_cse , act_regs_data_and_524_cse , act_regs_data_and_525_cse
          , act_regs_data_and_526_cse , act_regs_data_and_527_cse , act_regs_data_and_528_cse
          , act_regs_data_and_529_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_4_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_583 | or_dcpl_490 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_1_4_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_253_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_4_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1331_tmp ) begin
      act_regs_data_1_4_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_1_4_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[158:128]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_5_exs_5_30_0, Relu_for_y_qr_30_0_5_lpi_1_dfm, Silu_for_y_5_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_523_cse , act_regs_data_and_524_cse , act_regs_data_and_525_cse
          , act_regs_data_and_526_cse , act_regs_data_and_527_cse , act_regs_data_and_528_cse
          , act_regs_data_and_529_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_5_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_583 | or_dcpl_493 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_1_5_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_252_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_5_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1333_tmp ) begin
      act_regs_data_1_5_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_1_5_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[190:160]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_6_exs_5_30_0, Relu_for_y_qr_30_0_6_lpi_1_dfm, Silu_for_y_6_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_523_cse , act_regs_data_and_524_cse , act_regs_data_and_525_cse
          , act_regs_data_and_526_cse , act_regs_data_and_527_cse , act_regs_data_and_528_cse
          , act_regs_data_and_529_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_6_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_586 | or_dcpl_490 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_1_6_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_251_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_6_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1335_tmp ) begin
      act_regs_data_1_6_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_1_6_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[222:192]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_7_exs_5_30_0, Relu_for_y_qr_30_0_7_lpi_1_dfm, Silu_for_y_7_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_523_cse , act_regs_data_and_524_cse , act_regs_data_and_525_cse
          , act_regs_data_and_526_cse , act_regs_data_and_527_cse , act_regs_data_and_528_cse
          , act_regs_data_and_529_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_7_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_586 | or_dcpl_493 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_1_7_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_250_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_7_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1337_tmp ) begin
      act_regs_data_1_7_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_1_7_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[254:224]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_8_exs_5_30_0, Relu_for_y_qr_30_0_8_lpi_1_dfm, Silu_for_y_8_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_523_cse , act_regs_data_and_524_cse , act_regs_data_and_525_cse
          , act_regs_data_and_526_cse , act_regs_data_and_527_cse , act_regs_data_and_528_cse
          , act_regs_data_and_529_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_8_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_583 | or_dcpl_464 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_1_8_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_249_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_8_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1339_tmp ) begin
      act_regs_data_1_8_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_1_8_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[286:256]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_9_exs_5_30_0, Relu_for_y_qr_30_0_9_lpi_1_dfm, Silu_for_y_9_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_523_cse , act_regs_data_and_524_cse , act_regs_data_and_525_cse
          , act_regs_data_and_526_cse , act_regs_data_and_527_cse , act_regs_data_and_528_cse
          , act_regs_data_and_529_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_9_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_583 | or_dcpl_471 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_1_9_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_248_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_9_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1341_tmp ) begin
      act_regs_data_1_9_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_1_9_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[318:288]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_10_exs_5_30_0, Relu_for_y_qr_30_0_10_lpi_1_dfm, ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_30_0,
          Gelu_for_y_10_lpi_1_dfm_2_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_523_cse , act_regs_data_and_524_cse , act_regs_data_and_525_cse
          , act_regs_data_and_526_cse , act_regs_data_and_527_cse , act_regs_data_and_528_cse
          , act_regs_data_and_529_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_10_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_586 | or_dcpl_464 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_1_10_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_247_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_10_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1343_tmp ) begin
      act_regs_data_1_10_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_1_10_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[350:320]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_11_exs_5_30_0, Relu_for_y_qr_30_0_11_lpi_1_dfm, ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_30_0,
          Gelu_for_y_11_lpi_1_dfm_2_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_523_cse , act_regs_data_and_524_cse , act_regs_data_and_525_cse
          , act_regs_data_and_526_cse , act_regs_data_and_527_cse , act_regs_data_and_528_cse
          , act_regs_data_and_529_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_11_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_586 | or_dcpl_471 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_1_11_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_246_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_11_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1345_tmp ) begin
      act_regs_data_1_11_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_1_11_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[382:352]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_12_exs_5_30_0, Relu_for_y_qr_30_0_12_lpi_1_dfm, Silu_for_y_12_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_523_cse , act_regs_data_and_524_cse , act_regs_data_and_525_cse
          , act_regs_data_and_526_cse , act_regs_data_and_527_cse , act_regs_data_and_528_cse
          , act_regs_data_and_529_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_12_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_583 | or_dcpl_475 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_1_12_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_245_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_12_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1347_tmp ) begin
      act_regs_data_1_12_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_1_12_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[414:384]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_13_exs_5_30_0, Relu_for_y_qr_30_0_13_lpi_1_dfm, Silu_for_y_13_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_1_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_523_cse , act_regs_data_and_524_cse , act_regs_data_and_525_cse
          , act_regs_data_and_526_cse , act_regs_data_and_527_cse , act_regs_data_and_528_cse
          , act_regs_data_and_529_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_13_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_583 | or_dcpl_478 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_1_13_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_244_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_13_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1349_tmp ) begin
      act_regs_data_1_13_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_1_13_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[446:416]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_14_exs_5_30_0, Relu_for_y_qr_30_0_14_lpi_1_dfm, Silu_for_y_14_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_523_cse , act_regs_data_and_524_cse , act_regs_data_and_525_cse
          , act_regs_data_and_526_cse , act_regs_data_and_527_cse , act_regs_data_and_528_cse
          , act_regs_data_and_529_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_14_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_586 | or_dcpl_475 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_1_14_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_243_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_14_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1351_tmp ) begin
      act_regs_data_1_14_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_1_14_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[478:448]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_15_exs_5_30_0, Relu_for_y_qr_30_0_15_lpi_1_dfm, Silu_for_y_15_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_523_cse , act_regs_data_and_524_cse , act_regs_data_and_525_cse
          , act_regs_data_and_526_cse , act_regs_data_and_527_cse , act_regs_data_and_528_cse
          , act_regs_data_and_529_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_15_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_586 | or_dcpl_478 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_1_15_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_242_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_15_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1353_tmp ) begin
      act_regs_data_1_15_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_1_15_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[510:480]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_16_exs_5_30_0, Relu_for_y_qr_30_0_lpi_1_dfm, Silu_for_y_lpi_1_dfm_1_30_0,
          Gelu_for_y_lpi_1_dfm_2_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_523_cse , act_regs_data_and_524_cse , act_regs_data_and_525_cse
          , act_regs_data_and_526_cse , act_regs_data_and_527_cse , act_regs_data_and_528_cse
          , act_regs_data_and_529_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_0_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_602 | or_dcpl_451 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_2_0_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_241_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_0_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1355_tmp ) begin
      act_regs_data_2_0_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_2_0_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[30:0]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_1_exs_5_30_0, Relu_for_y_qr_30_0_1_lpi_1_dfm, ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_30_0,
          ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_635_cse , act_regs_data_and_636_cse , act_regs_data_and_637_cse
          , act_regs_data_and_638_cse , act_regs_data_and_639_cse , act_regs_data_and_640_cse
          , act_regs_data_and_641_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_1_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_602 | or_dcpl_458 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_2_1_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_240_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_1_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1357_tmp ) begin
      act_regs_data_2_1_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_2_1_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[62:32]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_2_exs_5_30_0, Relu_for_y_qr_30_0_2_lpi_1_dfm, Silu_for_y_2_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_635_cse , act_regs_data_and_636_cse , act_regs_data_and_637_cse
          , act_regs_data_and_638_cse , act_regs_data_and_639_cse , act_regs_data_and_640_cse
          , act_regs_data_and_641_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_2_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_605 | or_dcpl_451 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_2_2_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_239_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_2_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1359_tmp ) begin
      act_regs_data_2_2_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_2_2_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[94:64]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_3_exs_5_30_0, Relu_for_y_qr_30_0_3_lpi_1_dfm, Silu_for_y_3_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_635_cse , act_regs_data_and_636_cse , act_regs_data_and_637_cse
          , act_regs_data_and_638_cse , act_regs_data_and_639_cse , act_regs_data_and_640_cse
          , act_regs_data_and_641_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_3_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_605 | or_dcpl_458 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_2_3_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_238_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_3_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1361_tmp ) begin
      act_regs_data_2_3_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_2_3_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[126:96]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_4_exs_5_30_0, Relu_for_y_qr_30_0_4_lpi_1_dfm, Silu_for_y_4_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_635_cse , act_regs_data_and_636_cse , act_regs_data_and_637_cse
          , act_regs_data_and_638_cse , act_regs_data_and_639_cse , act_regs_data_and_640_cse
          , act_regs_data_and_641_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_4_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_602 | or_dcpl_490 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_2_4_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_237_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_4_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1363_tmp ) begin
      act_regs_data_2_4_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_2_4_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[158:128]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_5_exs_5_30_0, Relu_for_y_qr_30_0_5_lpi_1_dfm, Silu_for_y_5_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_635_cse , act_regs_data_and_636_cse , act_regs_data_and_637_cse
          , act_regs_data_and_638_cse , act_regs_data_and_639_cse , act_regs_data_and_640_cse
          , act_regs_data_and_641_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_5_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_602 | or_dcpl_493 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_2_5_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_236_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_5_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1365_tmp ) begin
      act_regs_data_2_5_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_2_5_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[190:160]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_6_exs_5_30_0, Relu_for_y_qr_30_0_6_lpi_1_dfm, Silu_for_y_6_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_635_cse , act_regs_data_and_636_cse , act_regs_data_and_637_cse
          , act_regs_data_and_638_cse , act_regs_data_and_639_cse , act_regs_data_and_640_cse
          , act_regs_data_and_641_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_6_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_605 | or_dcpl_490 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_2_6_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_235_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_6_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1367_tmp ) begin
      act_regs_data_2_6_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_2_6_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[222:192]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_7_exs_5_30_0, Relu_for_y_qr_30_0_7_lpi_1_dfm, Silu_for_y_7_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_635_cse , act_regs_data_and_636_cse , act_regs_data_and_637_cse
          , act_regs_data_and_638_cse , act_regs_data_and_639_cse , act_regs_data_and_640_cse
          , act_regs_data_and_641_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_7_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_605 | or_dcpl_493 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_2_7_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_234_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_7_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1369_tmp ) begin
      act_regs_data_2_7_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_2_7_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[254:224]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_8_exs_5_30_0, Relu_for_y_qr_30_0_8_lpi_1_dfm, Silu_for_y_8_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_635_cse , act_regs_data_and_636_cse , act_regs_data_and_637_cse
          , act_regs_data_and_638_cse , act_regs_data_and_639_cse , act_regs_data_and_640_cse
          , act_regs_data_and_641_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_8_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_602 | or_dcpl_464 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_2_8_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_233_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_8_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1371_tmp ) begin
      act_regs_data_2_8_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_2_8_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[286:256]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_9_exs_5_30_0, Relu_for_y_qr_30_0_9_lpi_1_dfm, Silu_for_y_9_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_635_cse , act_regs_data_and_636_cse , act_regs_data_and_637_cse
          , act_regs_data_and_638_cse , act_regs_data_and_639_cse , act_regs_data_and_640_cse
          , act_regs_data_and_641_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_9_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_602 | or_dcpl_471 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_2_9_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_232_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_9_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1373_tmp ) begin
      act_regs_data_2_9_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_2_9_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[318:288]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_10_exs_5_30_0, Relu_for_y_qr_30_0_10_lpi_1_dfm, ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_30_0,
          Gelu_for_y_10_lpi_1_dfm_2_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_635_cse , act_regs_data_and_636_cse , act_regs_data_and_637_cse
          , act_regs_data_and_638_cse , act_regs_data_and_639_cse , act_regs_data_and_640_cse
          , act_regs_data_and_641_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_10_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_605 | or_dcpl_464 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_2_10_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_231_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_10_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1375_tmp ) begin
      act_regs_data_2_10_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_2_10_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[350:320]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_11_exs_5_30_0, Relu_for_y_qr_30_0_11_lpi_1_dfm, ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_30_0,
          Gelu_for_y_11_lpi_1_dfm_2_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_635_cse , act_regs_data_and_636_cse , act_regs_data_and_637_cse
          , act_regs_data_and_638_cse , act_regs_data_and_639_cse , act_regs_data_and_640_cse
          , act_regs_data_and_641_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_11_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_605 | or_dcpl_471 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_2_11_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_230_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_11_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1377_tmp ) begin
      act_regs_data_2_11_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_2_11_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[382:352]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_12_exs_5_30_0, Relu_for_y_qr_30_0_12_lpi_1_dfm, Silu_for_y_12_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_635_cse , act_regs_data_and_636_cse , act_regs_data_and_637_cse
          , act_regs_data_and_638_cse , act_regs_data_and_639_cse , act_regs_data_and_640_cse
          , act_regs_data_and_641_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_12_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_602 | or_dcpl_475 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_2_12_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_229_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_12_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1379_tmp ) begin
      act_regs_data_2_12_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_2_12_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[414:384]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_13_exs_5_30_0, Relu_for_y_qr_30_0_13_lpi_1_dfm, Silu_for_y_13_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_1_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_635_cse , act_regs_data_and_636_cse , act_regs_data_and_637_cse
          , act_regs_data_and_638_cse , act_regs_data_and_639_cse , act_regs_data_and_640_cse
          , act_regs_data_and_641_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_13_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_602 | or_dcpl_478 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_2_13_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_228_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_13_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1381_tmp ) begin
      act_regs_data_2_13_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_2_13_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[446:416]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_14_exs_5_30_0, Relu_for_y_qr_30_0_14_lpi_1_dfm, Silu_for_y_14_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_635_cse , act_regs_data_and_636_cse , act_regs_data_and_637_cse
          , act_regs_data_and_638_cse , act_regs_data_and_639_cse , act_regs_data_and_640_cse
          , act_regs_data_and_641_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_14_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_605 | or_dcpl_475 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_2_14_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_227_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_14_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1383_tmp ) begin
      act_regs_data_2_14_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_2_14_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[478:448]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_15_exs_5_30_0, Relu_for_y_qr_30_0_15_lpi_1_dfm, Silu_for_y_15_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_635_cse , act_regs_data_and_636_cse , act_regs_data_and_637_cse
          , act_regs_data_and_638_cse , act_regs_data_and_639_cse , act_regs_data_and_640_cse
          , act_regs_data_and_641_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_15_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_605 | or_dcpl_478 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_2_15_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_226_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_15_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1385_tmp ) begin
      act_regs_data_2_15_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_2_15_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[510:480]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_16_exs_5_30_0, Relu_for_y_qr_30_0_lpi_1_dfm, Silu_for_y_lpi_1_dfm_1_30_0,
          Gelu_for_y_lpi_1_dfm_2_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_635_cse , act_regs_data_and_636_cse , act_regs_data_and_637_cse
          , act_regs_data_and_638_cse , act_regs_data_and_639_cse , act_regs_data_and_640_cse
          , act_regs_data_and_641_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_0_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_621 | or_dcpl_451 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_3_0_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_225_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_0_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1387_tmp ) begin
      act_regs_data_3_0_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_3_0_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[30:0]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_1_exs_5_30_0, Relu_for_y_qr_30_0_1_lpi_1_dfm, ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_30_0,
          ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_747_cse , act_regs_data_and_748_cse , act_regs_data_and_749_cse
          , act_regs_data_and_750_cse , act_regs_data_and_751_cse , act_regs_data_and_752_cse
          , act_regs_data_and_753_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_1_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_621 | or_dcpl_458 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_3_1_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_224_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_1_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1389_tmp ) begin
      act_regs_data_3_1_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_3_1_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[62:32]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_2_exs_5_30_0, Relu_for_y_qr_30_0_2_lpi_1_dfm, Silu_for_y_2_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_747_cse , act_regs_data_and_748_cse , act_regs_data_and_749_cse
          , act_regs_data_and_750_cse , act_regs_data_and_751_cse , act_regs_data_and_752_cse
          , act_regs_data_and_753_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_2_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_624 | or_dcpl_451 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_3_2_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_223_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_2_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1391_tmp ) begin
      act_regs_data_3_2_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_3_2_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[94:64]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_3_exs_5_30_0, Relu_for_y_qr_30_0_3_lpi_1_dfm, Silu_for_y_3_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_747_cse , act_regs_data_and_748_cse , act_regs_data_and_749_cse
          , act_regs_data_and_750_cse , act_regs_data_and_751_cse , act_regs_data_and_752_cse
          , act_regs_data_and_753_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_3_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_624 | or_dcpl_458 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_3_3_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_222_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_3_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1393_tmp ) begin
      act_regs_data_3_3_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_3_3_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[126:96]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_4_exs_5_30_0, Relu_for_y_qr_30_0_4_lpi_1_dfm, Silu_for_y_4_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_747_cse , act_regs_data_and_748_cse , act_regs_data_and_749_cse
          , act_regs_data_and_750_cse , act_regs_data_and_751_cse , act_regs_data_and_752_cse
          , act_regs_data_and_753_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_4_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_621 | or_dcpl_490 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_3_4_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_221_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_4_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1395_tmp ) begin
      act_regs_data_3_4_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_3_4_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[158:128]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_5_exs_5_30_0, Relu_for_y_qr_30_0_5_lpi_1_dfm, Silu_for_y_5_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_747_cse , act_regs_data_and_748_cse , act_regs_data_and_749_cse
          , act_regs_data_and_750_cse , act_regs_data_and_751_cse , act_regs_data_and_752_cse
          , act_regs_data_and_753_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_5_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_621 | or_dcpl_493 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_3_5_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_220_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_5_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1397_tmp ) begin
      act_regs_data_3_5_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_3_5_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[190:160]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_6_exs_5_30_0, Relu_for_y_qr_30_0_6_lpi_1_dfm, Silu_for_y_6_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_747_cse , act_regs_data_and_748_cse , act_regs_data_and_749_cse
          , act_regs_data_and_750_cse , act_regs_data_and_751_cse , act_regs_data_and_752_cse
          , act_regs_data_and_753_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_6_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_624 | or_dcpl_490 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_3_6_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_219_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_6_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1399_tmp ) begin
      act_regs_data_3_6_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_3_6_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[222:192]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_7_exs_5_30_0, Relu_for_y_qr_30_0_7_lpi_1_dfm, Silu_for_y_7_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_747_cse , act_regs_data_and_748_cse , act_regs_data_and_749_cse
          , act_regs_data_and_750_cse , act_regs_data_and_751_cse , act_regs_data_and_752_cse
          , act_regs_data_and_753_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_7_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_624 | or_dcpl_493 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_3_7_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_218_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_7_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1401_tmp ) begin
      act_regs_data_3_7_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_3_7_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[254:224]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_8_exs_5_30_0, Relu_for_y_qr_30_0_8_lpi_1_dfm, Silu_for_y_8_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_747_cse , act_regs_data_and_748_cse , act_regs_data_and_749_cse
          , act_regs_data_and_750_cse , act_regs_data_and_751_cse , act_regs_data_and_752_cse
          , act_regs_data_and_753_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_8_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_621 | or_dcpl_464 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_3_8_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_217_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_8_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1403_tmp ) begin
      act_regs_data_3_8_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_3_8_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[286:256]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_9_exs_5_30_0, Relu_for_y_qr_30_0_9_lpi_1_dfm, Silu_for_y_9_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_747_cse , act_regs_data_and_748_cse , act_regs_data_and_749_cse
          , act_regs_data_and_750_cse , act_regs_data_and_751_cse , act_regs_data_and_752_cse
          , act_regs_data_and_753_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_9_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_621 | or_dcpl_471 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_3_9_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_216_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_9_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1405_tmp ) begin
      act_regs_data_3_9_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_3_9_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[318:288]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_10_exs_5_30_0, Relu_for_y_qr_30_0_10_lpi_1_dfm, ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_30_0,
          Gelu_for_y_10_lpi_1_dfm_2_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_747_cse , act_regs_data_and_748_cse , act_regs_data_and_749_cse
          , act_regs_data_and_750_cse , act_regs_data_and_751_cse , act_regs_data_and_752_cse
          , act_regs_data_and_753_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_10_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_624 | or_dcpl_464 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_3_10_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_215_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_10_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1407_tmp ) begin
      act_regs_data_3_10_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_3_10_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[350:320]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_11_exs_5_30_0, Relu_for_y_qr_30_0_11_lpi_1_dfm, ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_30_0,
          Gelu_for_y_11_lpi_1_dfm_2_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_747_cse , act_regs_data_and_748_cse , act_regs_data_and_749_cse
          , act_regs_data_and_750_cse , act_regs_data_and_751_cse , act_regs_data_and_752_cse
          , act_regs_data_and_753_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_11_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_624 | or_dcpl_471 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_3_11_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_214_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_11_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1409_tmp ) begin
      act_regs_data_3_11_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_3_11_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[382:352]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_12_exs_5_30_0, Relu_for_y_qr_30_0_12_lpi_1_dfm, Silu_for_y_12_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_747_cse , act_regs_data_and_748_cse , act_regs_data_and_749_cse
          , act_regs_data_and_750_cse , act_regs_data_and_751_cse , act_regs_data_and_752_cse
          , act_regs_data_and_753_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_12_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_621 | or_dcpl_475 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_3_12_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_213_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_12_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1411_tmp ) begin
      act_regs_data_3_12_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_3_12_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[414:384]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_13_exs_5_30_0, Relu_for_y_qr_30_0_13_lpi_1_dfm, Silu_for_y_13_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_1_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_747_cse , act_regs_data_and_748_cse , act_regs_data_and_749_cse
          , act_regs_data_and_750_cse , act_regs_data_and_751_cse , act_regs_data_and_752_cse
          , act_regs_data_and_753_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_13_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_621 | or_dcpl_478 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_3_13_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_212_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_13_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1413_tmp ) begin
      act_regs_data_3_13_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_3_13_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[446:416]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_14_exs_5_30_0, Relu_for_y_qr_30_0_14_lpi_1_dfm, Silu_for_y_14_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_747_cse , act_regs_data_and_748_cse , act_regs_data_and_749_cse
          , act_regs_data_and_750_cse , act_regs_data_and_751_cse , act_regs_data_and_752_cse
          , act_regs_data_and_753_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_14_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_624 | or_dcpl_475 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_3_14_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_211_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_14_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1415_tmp ) begin
      act_regs_data_3_14_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_3_14_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[478:448]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_15_exs_5_30_0, Relu_for_y_qr_30_0_15_lpi_1_dfm, Silu_for_y_15_lpi_1_dfm_1_30_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_747_cse , act_regs_data_and_748_cse , act_regs_data_and_749_cse
          , act_regs_data_and_750_cse , act_regs_data_and_751_cse , act_regs_data_and_752_cse
          , act_regs_data_and_753_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_15_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_624 | or_dcpl_478 | (~ mux_235_itm)))
        | and_dcpl_997) ) begin
      act_regs_data_3_15_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_849);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_15_sva_dfm_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_1417_tmp ) begin
      act_regs_data_3_15_sva_dfm_2_30_0 <= MUX1HOT_v_31_8_2(act_regs_data_3_15_sva_30_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[510:480]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_0,
          Tanh_for_16_exs_5_30_0, Relu_for_y_qr_30_0_lpi_1_dfm, Silu_for_y_lpi_1_dfm_1_30_0,
          Gelu_for_y_lpi_1_dfm_2_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
          {act_regs_data_and_747_cse , act_regs_data_and_748_cse , act_regs_data_and_749_cse
          , act_regs_data_and_750_cse , act_regs_data_and_751_cse , act_regs_data_and_752_cse
          , act_regs_data_and_753_cse , and_dcpl_849});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_get_slc_2U_NVUINT8_return_3_sva <= 2'b00;
    end
    else if ( ActUnitRun_wen & (~ and_dcpl_799) & and_dcpl_370 & (~(act_config_is_zero_first_sva_dfm_4
        | act_config_is_zero_first_sva)) ) begin
      nvhls_get_slc_2U_NVUINT8_return_3_sva <= nvhls_get_slc_2U_NVUINT8_return_3_sva_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_config_InstIncr_if_act_config_InstIncr_if_if_nor_mdf_sva <= 1'b0;
    end
    else if ( ActUnitRun_wen & mux_82_nl & while_asn_262_itm & is_incr_lpi_1_dfm_1
        ) begin
      act_config_InstIncr_if_act_config_InstIncr_if_if_nor_mdf_sva <= act_config_InstIncr_if_act_config_InstIncr_if_if_nor_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_else_1_mux_1_itm <= 1'b0;
    end
    else if ( ActUnitRun_wen & while_asn_262_itm ) begin
      while_else_1_mux_1_itm <= MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4, act_config_InstIncr_mux_2_nl,
          is_incr_lpi_1_dfm_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_23_4_ftd_12
          <= 8'b00000000;
    end
    else if ( mux_578_nl & (~((fsm_output[4]) | is_start_sva)) & ActUnitRun_wen &
        (fsm_output[1]) & nor_734_cse & (fsm_output[0]) ) begin
      reg_ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_23_4_ftd_12
          <= ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_23_4_mx1_tmp_7_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_RunInst_case_11_nv_scvector_cctor_data_0_ftd_6 <= 26'b00000000000000000000000000;
    end
    else if ( ActUnit_RunInst_switch_lp_and_817_enex5 ) begin
      reg_ActUnit_RunInst_case_11_nv_scvector_cctor_data_0_ftd_6 <= ActUnit_RunInst_case_11_nv_scvector_cctor_data_0_sva_1_30_0[25:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6
          <= 26'b00000000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_3_for_and_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6
          <= nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[25:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6
          <= 26'b00000000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_3_for_and_15_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6
          <= nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[25:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6
          <= 26'b00000000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_3_for_and_16_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6
          <= nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[25:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6
          <= 26'b00000000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_3_for_and_17_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6
          <= nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[25:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6
          <= 26'b00000000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_3_for_and_18_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6
          <= nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[25:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6
          <= 26'b00000000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_3_for_and_19_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6
          <= nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[25:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6
          <= 26'b00000000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_3_for_and_20_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6
          <= nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[25:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6
          <= 26'b00000000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_3_for_and_21_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6
          <= nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[25:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6
          <= 26'b00000000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_3_for_and_22_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6
          <= nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[25:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6
          <= 26'b00000000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_3_for_and_23_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6
          <= nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[25:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6
          <= 26'b00000000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_3_for_and_24_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6
          <= nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[25:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6
          <= 26'b00000000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_3_for_and_25_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_ftd_6
          <= nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_30_0[25:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_15_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_284_cse | act_regs_data_and_859_enex5 ) begin
      reg_act_regs_data_3_15_3_enexo <= act_regs_data_and_284_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_2_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_108_ssc | act_regs_data_and_859_enex5 ) begin
      reg_act_regs_data_2_2_3_enexo <= act_regs_data_and_108_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_859_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_859_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_859_enex5 ) begin
      reg_is_start_enexo <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_15_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1417_tmp | act_regs_data_and_859_enex5 ) begin
      reg_act_regs_data_3_15_sva_dfm_2_1_enexo <= and_1417_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_15_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_95_ssc | act_regs_data_and_860_enex5 ) begin
      reg_act_regs_data_2_15_3_enexo <= act_regs_data_and_95_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_14_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_284_cse | act_regs_data_and_860_enex5 ) begin
      reg_act_regs_data_3_14_3_enexo <= act_regs_data_and_284_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_1 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_860_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_1 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_1 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_860_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_1 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_1 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_860_enex5 ) begin
      reg_is_start_enexo_1 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_14_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1415_tmp | act_regs_data_and_860_enex5 ) begin
      reg_act_regs_data_3_14_sva_dfm_2_1_enexo <= and_1415_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_14_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_96_ssc | act_regs_data_and_861_enex5 ) begin
      reg_act_regs_data_2_14_3_enexo <= act_regs_data_and_96_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_13_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_284_cse | act_regs_data_and_861_enex5 ) begin
      reg_act_regs_data_3_13_3_enexo <= act_regs_data_and_284_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_2 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_861_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_2 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_2 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_861_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_2 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_2 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_861_enex5 ) begin
      reg_is_start_enexo_2 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_13_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1413_tmp | act_regs_data_and_861_enex5 ) begin
      reg_act_regs_data_3_13_sva_dfm_2_1_enexo <= and_1413_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_12_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_284_cse | act_regs_data_and_862_enex5 ) begin
      reg_act_regs_data_3_12_3_enexo <= act_regs_data_and_284_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_3 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_862_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_3 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_13_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_97_ssc | act_regs_data_and_862_enex5 ) begin
      reg_act_regs_data_2_13_3_enexo <= act_regs_data_and_97_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_3 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_862_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_3 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_3 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_862_enex5 ) begin
      reg_is_start_enexo_3 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_12_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1411_tmp | act_regs_data_and_862_enex5 ) begin
      reg_act_regs_data_3_12_sva_dfm_2_1_enexo <= and_1411_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_11_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_284_cse | act_regs_data_and_863_enex5 ) begin
      reg_act_regs_data_3_11_3_enexo <= act_regs_data_and_284_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_4 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_863_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_4 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_12_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_98_ssc | act_regs_data_and_863_enex5 ) begin
      reg_act_regs_data_2_12_3_enexo <= act_regs_data_and_98_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_4 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_863_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_4 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_4 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_863_enex5 ) begin
      reg_is_start_enexo_4 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_11_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1409_tmp | act_regs_data_and_863_enex5 ) begin
      reg_act_regs_data_3_11_sva_dfm_2_1_enexo <= and_1409_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_10_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_284_cse | act_regs_data_and_864_enex5 ) begin
      reg_act_regs_data_3_10_3_enexo <= act_regs_data_and_284_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_5 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_864_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_5 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_11_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_99_ssc | act_regs_data_and_864_enex5 ) begin
      reg_act_regs_data_2_11_3_enexo <= act_regs_data_and_99_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_5 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_864_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_5 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_5 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_864_enex5 ) begin
      reg_is_start_enexo_5 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_10_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1407_tmp | act_regs_data_and_864_enex5 ) begin
      reg_act_regs_data_3_10_sva_dfm_2_1_enexo <= and_1407_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_0_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_94_ssc | act_regs_data_and_865_enex5 ) begin
      reg_act_regs_data_3_0_3_enexo <= act_regs_data_and_94_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_9_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_284_cse | act_regs_data_and_865_enex5 ) begin
      reg_act_regs_data_3_9_3_enexo <= act_regs_data_and_284_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_6 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_865_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_6 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_6 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_865_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_6 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_6 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_865_enex5 ) begin
      reg_is_start_enexo_6 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_9_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1405_tmp | act_regs_data_and_865_enex5 ) begin
      reg_act_regs_data_3_9_sva_dfm_2_1_enexo <= and_1405_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_8_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_284_cse | act_regs_data_and_866_enex5 ) begin
      reg_act_regs_data_3_8_3_enexo <= act_regs_data_and_284_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_7 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_866_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_7 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_9_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_101_ssc | act_regs_data_and_866_enex5 ) begin
      reg_act_regs_data_2_9_3_enexo <= act_regs_data_and_101_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_7 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_866_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_7 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_7 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_866_enex5 ) begin
      reg_is_start_enexo_7 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_8_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1403_tmp | act_regs_data_and_866_enex5 ) begin
      reg_act_regs_data_3_8_sva_dfm_2_1_enexo <= and_1403_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_7_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_284_cse | act_regs_data_and_867_enex5 ) begin
      reg_act_regs_data_3_7_3_enexo <= act_regs_data_and_284_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_8 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_867_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_8 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_8_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_102_ssc | act_regs_data_and_867_enex5 ) begin
      reg_act_regs_data_2_8_3_enexo <= act_regs_data_and_102_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_8 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_867_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_8 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_8 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_867_enex5 ) begin
      reg_is_start_enexo_8 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_7_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1401_tmp | act_regs_data_and_867_enex5 ) begin
      reg_act_regs_data_3_7_sva_dfm_2_1_enexo <= and_1401_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_6_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_284_cse | act_regs_data_and_868_enex5 ) begin
      reg_act_regs_data_3_6_3_enexo <= act_regs_data_and_284_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_9 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_868_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_9 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_7_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_103_ssc | act_regs_data_and_868_enex5 ) begin
      reg_act_regs_data_2_7_3_enexo <= act_regs_data_and_103_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_9 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_868_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_9 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_9 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_868_enex5 ) begin
      reg_is_start_enexo_9 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_6_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1399_tmp | act_regs_data_and_868_enex5 ) begin
      reg_act_regs_data_3_6_sva_dfm_2_1_enexo <= and_1399_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_5_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_284_cse | act_regs_data_and_869_enex5 ) begin
      reg_act_regs_data_3_5_3_enexo <= act_regs_data_and_284_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_10 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_869_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_10 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_6_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_104_ssc | act_regs_data_and_869_enex5 ) begin
      reg_act_regs_data_2_6_3_enexo <= act_regs_data_and_104_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_10 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_869_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_10 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_10 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_869_enex5 ) begin
      reg_is_start_enexo_10 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_5_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1397_tmp | act_regs_data_and_869_enex5 ) begin
      reg_act_regs_data_3_5_sva_dfm_2_1_enexo <= and_1397_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_4_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_284_cse | act_regs_data_and_870_enex5 ) begin
      reg_act_regs_data_3_4_3_enexo <= act_regs_data_and_284_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_11 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_870_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_11 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_5_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_105_ssc | act_regs_data_and_870_enex5 ) begin
      reg_act_regs_data_2_5_3_enexo <= act_regs_data_and_105_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_11 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_870_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_11 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_11 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_870_enex5 ) begin
      reg_is_start_enexo_11 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_4_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1395_tmp | act_regs_data_and_870_enex5 ) begin
      reg_act_regs_data_3_4_sva_dfm_2_1_enexo <= and_1395_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_3_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_284_cse | act_regs_data_and_871_enex5 ) begin
      reg_act_regs_data_3_3_3_enexo <= act_regs_data_and_284_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_12 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_871_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_12 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_4_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_106_ssc | act_regs_data_and_871_enex5 ) begin
      reg_act_regs_data_2_4_3_enexo <= act_regs_data_and_106_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_12 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_871_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_12 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_12 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_871_enex5 ) begin
      reg_is_start_enexo_12 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_3_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1393_tmp | act_regs_data_and_871_enex5 ) begin
      reg_act_regs_data_3_3_sva_dfm_2_1_enexo <= and_1393_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_2_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_284_cse | act_regs_data_and_872_enex5 ) begin
      reg_act_regs_data_3_2_3_enexo <= act_regs_data_and_284_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_3_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_107_ssc | act_regs_data_and_872_enex5 ) begin
      reg_act_regs_data_2_3_3_enexo <= act_regs_data_and_107_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_13 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_872_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_13 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_13 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_872_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_13 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_13 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_872_enex5 ) begin
      reg_is_start_enexo_13 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_2_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1391_tmp | act_regs_data_and_872_enex5 ) begin
      reg_act_regs_data_3_2_sva_dfm_2_1_enexo <= and_1391_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_1_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_284_cse | act_regs_data_and_873_enex5 ) begin
      reg_act_regs_data_3_1_3_enexo <= act_regs_data_and_284_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_14 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_873_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_14 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_10_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_100_ssc | act_regs_data_and_873_enex5 ) begin
      reg_act_regs_data_2_10_3_enexo <= act_regs_data_and_100_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_14 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_873_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_14 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_14 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_873_enex5 ) begin
      reg_is_start_enexo_14 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_1_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1389_tmp | act_regs_data_and_873_enex5 ) begin
      reg_act_regs_data_3_1_sva_dfm_2_1_enexo <= and_1389_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_0_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_94_ssc | act_regs_data_and_874_enex5 ) begin
      reg_act_regs_data_3_0_3_enexo_1 <= act_regs_data_and_94_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_1_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_109_ssc | act_regs_data_and_874_enex5 ) begin
      reg_act_regs_data_2_1_3_enexo <= act_regs_data_and_109_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_15 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_874_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_15 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_15 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_874_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_15 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_15 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_874_enex5 ) begin
      reg_is_start_enexo_15 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_0_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1387_tmp | act_regs_data_and_874_enex5 ) begin
      reg_act_regs_data_3_0_sva_dfm_2_1_enexo <= and_1387_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_15_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_95_ssc | act_regs_data_and_875_enex5 ) begin
      reg_act_regs_data_2_15_3_enexo_1 <= act_regs_data_and_95_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_16 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_875_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_16 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_16 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_875_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_16 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_2_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_124_ssc | act_regs_data_and_875_enex5 ) begin
      reg_act_regs_data_1_2_3_enexo <= act_regs_data_and_124_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_16 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_875_enex5 ) begin
      reg_is_start_enexo_16 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_15_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1385_tmp | act_regs_data_and_875_enex5 ) begin
      reg_act_regs_data_2_15_sva_dfm_2_1_enexo <= and_1385_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_14_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_96_ssc | act_regs_data_and_876_enex5 ) begin
      reg_act_regs_data_2_14_3_enexo_1 <= act_regs_data_and_96_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_15_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_111_ssc | act_regs_data_and_876_enex5 ) begin
      reg_act_regs_data_1_15_3_enexo <= act_regs_data_and_111_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_17 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_876_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_17 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_17 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_876_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_17 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_17 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_876_enex5 ) begin
      reg_is_start_enexo_17 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_14_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1383_tmp | act_regs_data_and_876_enex5 ) begin
      reg_act_regs_data_2_14_sva_dfm_2_1_enexo <= and_1383_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_14_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_112_ssc | act_regs_data_and_877_enex5 ) begin
      reg_act_regs_data_1_14_3_enexo <= act_regs_data_and_112_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_18 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_877_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_18 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_13_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_97_ssc | act_regs_data_and_877_enex5 ) begin
      reg_act_regs_data_2_13_3_enexo_1 <= act_regs_data_and_97_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_18 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_877_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_18 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_18 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_877_enex5 ) begin
      reg_is_start_enexo_18 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_13_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1381_tmp | act_regs_data_and_877_enex5 ) begin
      reg_act_regs_data_2_13_sva_dfm_2_1_enexo <= and_1381_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_13_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_113_ssc | act_regs_data_and_878_enex5 ) begin
      reg_act_regs_data_1_13_3_enexo <= act_regs_data_and_113_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_19 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_878_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_19 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_12_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_98_ssc | act_regs_data_and_878_enex5 ) begin
      reg_act_regs_data_2_12_3_enexo_1 <= act_regs_data_and_98_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_19 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_878_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_19 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_19 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_878_enex5 ) begin
      reg_is_start_enexo_19 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_12_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1379_tmp | act_regs_data_and_878_enex5 ) begin
      reg_act_regs_data_2_12_sva_dfm_2_1_enexo <= and_1379_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_12_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_114_ssc | act_regs_data_and_879_enex5 ) begin
      reg_act_regs_data_1_12_3_enexo <= act_regs_data_and_114_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_20 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_879_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_20 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_11_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_99_ssc | act_regs_data_and_879_enex5 ) begin
      reg_act_regs_data_2_11_3_enexo_1 <= act_regs_data_and_99_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_20 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_879_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_20 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_20 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_879_enex5 ) begin
      reg_is_start_enexo_20 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_11_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1377_tmp | act_regs_data_and_879_enex5 ) begin
      reg_act_regs_data_2_11_sva_dfm_2_1_enexo <= and_1377_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_11_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_115_ssc | act_regs_data_and_880_enex5 ) begin
      reg_act_regs_data_1_11_3_enexo <= act_regs_data_and_115_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_21 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_880_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_21 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_10_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_100_ssc | act_regs_data_and_880_enex5 ) begin
      reg_act_regs_data_2_10_3_enexo_1 <= act_regs_data_and_100_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_21 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_880_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_21 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_21 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_880_enex5 ) begin
      reg_is_start_enexo_21 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_10_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1375_tmp | act_regs_data_and_880_enex5 ) begin
      reg_act_regs_data_2_10_sva_dfm_2_1_enexo <= and_1375_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_0_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_110_ssc | act_regs_data_and_881_enex5 ) begin
      reg_act_regs_data_2_0_3_enexo <= act_regs_data_and_110_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_22 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_881_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_22 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_9_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_101_ssc | act_regs_data_and_881_enex5 ) begin
      reg_act_regs_data_2_9_3_enexo_1 <= act_regs_data_and_101_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_22 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_881_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_22 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_22 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_881_enex5 ) begin
      reg_is_start_enexo_22 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_9_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1373_tmp | act_regs_data_and_881_enex5 ) begin
      reg_act_regs_data_2_9_sva_dfm_2_1_enexo <= and_1373_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_23 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_882_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_23 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_8_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_102_ssc | act_regs_data_and_882_enex5 ) begin
      reg_act_regs_data_2_8_3_enexo_1 <= act_regs_data_and_102_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_23 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_882_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_23 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_9_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_117_ssc | act_regs_data_and_882_enex5 ) begin
      reg_act_regs_data_1_9_3_enexo <= act_regs_data_and_117_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_23 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_882_enex5 ) begin
      reg_is_start_enexo_23 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_8_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1371_tmp | act_regs_data_and_882_enex5 ) begin
      reg_act_regs_data_2_8_sva_dfm_2_1_enexo <= and_1371_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_24 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_883_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_24 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_7_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_103_ssc | act_regs_data_and_883_enex5 ) begin
      reg_act_regs_data_2_7_3_enexo_1 <= act_regs_data_and_103_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_24 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_883_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_24 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_8_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_118_ssc | act_regs_data_and_883_enex5 ) begin
      reg_act_regs_data_1_8_3_enexo <= act_regs_data_and_118_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_24 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_883_enex5 ) begin
      reg_is_start_enexo_24 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_7_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1369_tmp | act_regs_data_and_883_enex5 ) begin
      reg_act_regs_data_2_7_sva_dfm_2_1_enexo <= and_1369_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_25 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_884_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_25 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_6_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_104_ssc | act_regs_data_and_884_enex5 ) begin
      reg_act_regs_data_2_6_3_enexo_1 <= act_regs_data_and_104_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_25 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_884_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_25 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_7_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_119_ssc | act_regs_data_and_884_enex5 ) begin
      reg_act_regs_data_1_7_3_enexo <= act_regs_data_and_119_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_25 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_884_enex5 ) begin
      reg_is_start_enexo_25 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_6_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1367_tmp | act_regs_data_and_884_enex5 ) begin
      reg_act_regs_data_2_6_sva_dfm_2_1_enexo <= and_1367_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_26 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_885_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_26 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_5_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_105_ssc | act_regs_data_and_885_enex5 ) begin
      reg_act_regs_data_2_5_3_enexo_1 <= act_regs_data_and_105_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_26 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_885_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_26 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_6_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_120_ssc | act_regs_data_and_885_enex5 ) begin
      reg_act_regs_data_1_6_3_enexo <= act_regs_data_and_120_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_26 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_885_enex5 ) begin
      reg_is_start_enexo_26 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_5_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1365_tmp | act_regs_data_and_885_enex5 ) begin
      reg_act_regs_data_2_5_sva_dfm_2_1_enexo <= and_1365_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_27 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_886_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_27 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_4_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_106_ssc | act_regs_data_and_886_enex5 ) begin
      reg_act_regs_data_2_4_3_enexo_1 <= act_regs_data_and_106_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_27 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_886_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_27 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_5_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_121_ssc | act_regs_data_and_886_enex5 ) begin
      reg_act_regs_data_1_5_3_enexo <= act_regs_data_and_121_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_27 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_886_enex5 ) begin
      reg_is_start_enexo_27 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_4_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1363_tmp | act_regs_data_and_886_enex5 ) begin
      reg_act_regs_data_2_4_sva_dfm_2_1_enexo <= and_1363_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_3_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_107_ssc | act_regs_data_and_887_enex5 ) begin
      reg_act_regs_data_2_3_3_enexo_1 <= act_regs_data_and_107_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_28 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_887_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_28 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_28 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_887_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_28 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_4_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_122_ssc | act_regs_data_and_887_enex5 ) begin
      reg_act_regs_data_1_4_3_enexo <= act_regs_data_and_122_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_28 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_887_enex5 ) begin
      reg_is_start_enexo_28 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_3_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1361_tmp | act_regs_data_and_887_enex5 ) begin
      reg_act_regs_data_2_3_sva_dfm_2_1_enexo <= and_1361_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_2_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_108_ssc | act_regs_data_and_888_enex5 ) begin
      reg_act_regs_data_2_2_3_enexo_1 <= act_regs_data_and_108_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_29 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_888_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_29 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_29 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_888_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_29 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_3_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_123_ssc | act_regs_data_and_888_enex5 ) begin
      reg_act_regs_data_1_3_3_enexo <= act_regs_data_and_123_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_29 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_888_enex5 ) begin
      reg_is_start_enexo_29 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_2_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1359_tmp | act_regs_data_and_888_enex5 ) begin
      reg_act_regs_data_2_2_sva_dfm_2_1_enexo <= and_1359_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_1_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_109_ssc | act_regs_data_and_889_enex5 ) begin
      reg_act_regs_data_2_1_3_enexo_1 <= act_regs_data_and_109_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_10_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_116_ssc | act_regs_data_and_889_enex5 ) begin
      reg_act_regs_data_1_10_3_enexo <= act_regs_data_and_116_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_30 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_889_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_30 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_30 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_889_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_30 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_30 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_889_enex5 ) begin
      reg_is_start_enexo_30 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_1_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1357_tmp | act_regs_data_and_889_enex5 ) begin
      reg_act_regs_data_2_1_sva_dfm_2_1_enexo <= and_1357_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_0_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_110_ssc | act_regs_data_and_890_enex5 ) begin
      reg_act_regs_data_2_0_3_enexo_1 <= act_regs_data_and_110_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_31 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_890_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_31 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_31 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_890_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_31 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_1_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_125_ssc | act_regs_data_and_890_enex5 ) begin
      reg_act_regs_data_1_1_3_enexo <= act_regs_data_and_125_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_31 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_890_enex5 ) begin
      reg_is_start_enexo_31 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_0_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1355_tmp | act_regs_data_and_890_enex5 ) begin
      reg_act_regs_data_2_0_sva_dfm_2_1_enexo <= and_1355_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_15_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_111_ssc | act_regs_data_and_891_enex5 ) begin
      reg_act_regs_data_1_15_3_enexo_1 <= act_regs_data_and_111_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_32 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_891_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_32 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_32 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_891_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_32 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_2_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_72_ssc | act_regs_data_and_891_enex5 ) begin
      reg_act_regs_data_0_2_3_enexo <= act_regs_data_and_72_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_32 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_891_enex5 ) begin
      reg_is_start_enexo_32 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_15_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1353_tmp | act_regs_data_and_891_enex5 ) begin
      reg_act_regs_data_1_15_sva_dfm_2_1_enexo <= and_1353_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_14_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_112_ssc | act_regs_data_and_892_enex5 ) begin
      reg_act_regs_data_1_14_3_enexo_1 <= act_regs_data_and_112_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_33 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_892_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_33 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_33 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_892_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_33 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_33 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_892_enex5 ) begin
      reg_is_start_enexo_33 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_14_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1351_tmp | act_regs_data_and_892_enex5 ) begin
      reg_act_regs_data_1_14_sva_dfm_2_1_enexo <= and_1351_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_15_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_71_ssc | act_regs_data_and_892_enex5 ) begin
      reg_act_regs_data_0_15_3_enexo <= act_regs_data_and_71_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_13_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_113_ssc | act_regs_data_and_893_enex5 ) begin
      reg_act_regs_data_1_13_3_enexo_1 <= act_regs_data_and_113_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_34 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_893_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_34 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_34 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_893_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_34 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_34 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_893_enex5 ) begin
      reg_is_start_enexo_34 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_13_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1349_tmp | act_regs_data_and_893_enex5 ) begin
      reg_act_regs_data_1_13_sva_dfm_2_1_enexo <= and_1349_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_14_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_70_ssc | act_regs_data_and_893_enex5 ) begin
      reg_act_regs_data_0_14_3_enexo <= act_regs_data_and_70_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_12_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_114_ssc | act_regs_data_and_894_enex5 ) begin
      reg_act_regs_data_1_12_3_enexo_1 <= act_regs_data_and_114_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_35 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_894_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_35 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_35 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_894_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_35 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_35 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_894_enex5 ) begin
      reg_is_start_enexo_35 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_13_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_69_ssc | act_regs_data_and_894_enex5 ) begin
      reg_act_regs_data_0_13_3_enexo <= act_regs_data_and_69_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_12_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1347_tmp | act_regs_data_and_894_enex5 ) begin
      reg_act_regs_data_1_12_sva_dfm_2_1_enexo <= and_1347_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_11_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_115_ssc | act_regs_data_and_895_enex5 ) begin
      reg_act_regs_data_1_11_3_enexo_1 <= act_regs_data_and_115_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_36 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_895_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_36 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_36 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_895_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_36 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_36 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_895_enex5 ) begin
      reg_is_start_enexo_36 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_12_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_68_ssc | act_regs_data_and_895_enex5 ) begin
      reg_act_regs_data_0_12_3_enexo <= act_regs_data_and_68_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_11_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1345_tmp | act_regs_data_and_895_enex5 ) begin
      reg_act_regs_data_1_11_sva_dfm_2_1_enexo <= and_1345_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_10_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_116_ssc | act_regs_data_and_896_enex5 ) begin
      reg_act_regs_data_1_10_3_enexo_1 <= act_regs_data_and_116_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_37 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_896_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_37 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_37 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_896_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_37 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_37 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_896_enex5 ) begin
      reg_is_start_enexo_37 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_11_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_67_ssc | act_regs_data_and_896_enex5 ) begin
      reg_act_regs_data_0_11_3_enexo <= act_regs_data_and_67_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_10_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1343_tmp | act_regs_data_and_896_enex5 ) begin
      reg_act_regs_data_1_10_sva_dfm_2_1_enexo <= and_1343_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_0_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_126_ssc | act_regs_data_and_897_enex5 ) begin
      reg_act_regs_data_1_0_3_enexo <= act_regs_data_and_126_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_38 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_897_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_38 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_38 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_897_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_38 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_9_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_117_ssc | act_regs_data_and_897_enex5 ) begin
      reg_act_regs_data_1_9_3_enexo_1 <= act_regs_data_and_117_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_38 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_897_enex5 ) begin
      reg_is_start_enexo_38 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_9_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1341_tmp | act_regs_data_and_897_enex5 ) begin
      reg_act_regs_data_1_9_sva_dfm_2_1_enexo <= and_1341_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_9_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_127_ssc | act_regs_data_and_898_enex5 ) begin
      reg_act_regs_data_0_9_3_enexo <= act_regs_data_and_127_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_39 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_898_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_39 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_39 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_898_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_39 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_8_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_118_ssc | act_regs_data_and_898_enex5 ) begin
      reg_act_regs_data_1_8_3_enexo_1 <= act_regs_data_and_118_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_39 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_898_enex5 ) begin
      reg_is_start_enexo_39 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_8_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1339_tmp | act_regs_data_and_898_enex5 ) begin
      reg_act_regs_data_1_8_sva_dfm_2_1_enexo <= and_1339_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_40 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_899_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_40 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_8_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_78_ssc | act_regs_data_and_899_enex5 ) begin
      reg_act_regs_data_0_8_3_enexo <= act_regs_data_and_78_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_40 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_899_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_40 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_7_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_119_ssc | act_regs_data_and_899_enex5 ) begin
      reg_act_regs_data_1_7_3_enexo_1 <= act_regs_data_and_119_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_40 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_899_enex5 ) begin
      reg_is_start_enexo_40 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_7_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1337_tmp | act_regs_data_and_899_enex5 ) begin
      reg_act_regs_data_1_7_sva_dfm_2_1_enexo <= and_1337_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_41 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_900_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_41 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_7_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_77_ssc | act_regs_data_and_900_enex5 ) begin
      reg_act_regs_data_0_7_3_enexo <= act_regs_data_and_77_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_41 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_900_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_41 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_6_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_120_ssc | act_regs_data_and_900_enex5 ) begin
      reg_act_regs_data_1_6_3_enexo_1 <= act_regs_data_and_120_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_41 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_900_enex5 ) begin
      reg_is_start_enexo_41 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_6_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1335_tmp | act_regs_data_and_900_enex5 ) begin
      reg_act_regs_data_1_6_sva_dfm_2_1_enexo <= and_1335_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_6_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_76_ssc | act_regs_data_and_901_enex5 ) begin
      reg_act_regs_data_0_6_3_enexo <= act_regs_data_and_76_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_42 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_901_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_42 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_42 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_901_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_42 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_5_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_121_ssc | act_regs_data_and_901_enex5 ) begin
      reg_act_regs_data_1_5_3_enexo_1 <= act_regs_data_and_121_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_42 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_901_enex5 ) begin
      reg_is_start_enexo_42 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_5_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1333_tmp | act_regs_data_and_901_enex5 ) begin
      reg_act_regs_data_1_5_sva_dfm_2_1_enexo <= and_1333_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_5_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_75_ssc | act_regs_data_and_902_enex5 ) begin
      reg_act_regs_data_0_5_3_enexo <= act_regs_data_and_75_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_43 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_902_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_43 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_43 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_902_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_43 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_4_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_122_ssc | act_regs_data_and_902_enex5 ) begin
      reg_act_regs_data_1_4_3_enexo_1 <= act_regs_data_and_122_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_43 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_902_enex5 ) begin
      reg_is_start_enexo_43 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_4_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1331_tmp | act_regs_data_and_902_enex5 ) begin
      reg_act_regs_data_1_4_sva_dfm_2_1_enexo <= and_1331_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_44 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_903_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_44 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_44 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_903_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_44 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_4_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_74_ssc | act_regs_data_and_903_enex5 ) begin
      reg_act_regs_data_0_4_3_enexo <= act_regs_data_and_74_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_3_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_123_ssc | act_regs_data_and_903_enex5 ) begin
      reg_act_regs_data_1_3_3_enexo_1 <= act_regs_data_and_123_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_44 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_903_enex5 ) begin
      reg_is_start_enexo_44 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_3_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1329_tmp | act_regs_data_and_903_enex5 ) begin
      reg_act_regs_data_1_3_sva_dfm_2_1_enexo <= and_1329_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_45 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_904_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_45 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_45 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_904_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_45 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_3_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_73_ssc | act_regs_data_and_904_enex5 ) begin
      reg_act_regs_data_0_3_3_enexo <= act_regs_data_and_73_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_2_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_124_ssc | act_regs_data_and_904_enex5 ) begin
      reg_act_regs_data_1_2_3_enexo_1 <= act_regs_data_and_124_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_45 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_904_enex5 ) begin
      reg_is_start_enexo_45 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_2_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1327_tmp | act_regs_data_and_904_enex5 ) begin
      reg_act_regs_data_1_2_sva_dfm_2_1_enexo <= and_1327_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_46 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_905_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_46 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_46 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_905_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_46 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_1_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_125_ssc | act_regs_data_and_905_enex5 ) begin
      reg_act_regs_data_1_1_3_enexo_1 <= act_regs_data_and_125_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_46 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_905_enex5 ) begin
      reg_is_start_enexo_46 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_10_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_66_ssc | act_regs_data_and_905_enex5 ) begin
      reg_act_regs_data_0_10_3_enexo <= act_regs_data_and_66_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_1_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1325_tmp | act_regs_data_and_905_enex5 ) begin
      reg_act_regs_data_1_1_sva_dfm_2_1_enexo <= and_1325_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_0_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_126_ssc | act_regs_data_and_906_enex5 ) begin
      reg_act_regs_data_1_0_3_enexo_1 <= act_regs_data_and_126_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_47 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_906_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_47 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_47 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_906_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_47 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_1_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_65_ssc | act_regs_data_and_906_enex5 ) begin
      reg_act_regs_data_0_1_3_enexo <= act_regs_data_and_65_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_47 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_906_enex5 ) begin
      reg_is_start_enexo_47 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_0_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1323_tmp | act_regs_data_and_906_enex5 ) begin
      reg_act_regs_data_1_0_sva_dfm_2_1_enexo <= and_1323_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_48 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_907_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_48 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_48 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_907_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_48 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_2_1_enexo <= 1'b1;
    end
    else if ( and_1246_tmp | act_regs_data_and_907_enex5 ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_2_1_enexo <= and_1246_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_48 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_907_enex5 ) begin
      reg_is_start_enexo_48 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_15_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1321_tmp | act_regs_data_and_907_enex5 ) begin
      reg_act_regs_data_0_15_sva_dfm_2_1_enexo <= and_1321_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_15_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_71_ssc | act_regs_data_and_907_enex5 ) begin
      reg_act_regs_data_0_15_3_enexo_1 <= act_regs_data_and_71_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_49 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_908_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_49 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_49 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_908_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_49 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_14_1_enexo <= 1'b1;
    end
    else if ( and_1243_tmp | act_regs_data_and_908_enex5 ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_14_1_enexo <= and_1243_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_49 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_908_enex5 ) begin
      reg_is_start_enexo_49 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_14_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1319_tmp | act_regs_data_and_908_enex5 ) begin
      reg_act_regs_data_0_14_sva_dfm_2_1_enexo <= and_1319_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_14_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_70_ssc | act_regs_data_and_908_enex5 ) begin
      reg_act_regs_data_0_14_3_enexo_1 <= act_regs_data_and_70_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_50 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_909_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_50 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_50 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_909_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_50 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_50 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_909_enex5 ) begin
      reg_is_start_enexo_50 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_13_1_enexo <= 1'b1;
    end
    else if ( and_1237_tmp | act_regs_data_and_909_enex5 ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_13_1_enexo <= and_1237_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_13_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_69_ssc | act_regs_data_and_909_enex5 ) begin
      reg_act_regs_data_0_13_3_enexo_1 <= act_regs_data_and_69_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_13_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1317_tmp | act_regs_data_and_909_enex5 ) begin
      reg_act_regs_data_0_13_sva_dfm_2_1_enexo <= and_1317_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_51 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_910_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_51 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_51 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_910_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_51 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_12_1_enexo <= 1'b1;
    end
    else if ( and_1231_tmp | act_regs_data_and_910_enex5 ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_12_1_enexo <= and_1231_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_51 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_910_enex5 ) begin
      reg_is_start_enexo_51 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_12_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_68_ssc | act_regs_data_and_910_enex5 ) begin
      reg_act_regs_data_0_12_3_enexo_1 <= act_regs_data_and_68_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_12_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1315_tmp | act_regs_data_and_910_enex5 ) begin
      reg_act_regs_data_0_12_sva_dfm_2_1_enexo <= and_1315_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_52 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_911_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_52 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_11_1_enexo <= 1'b1;
    end
    else if ( and_1275_tmp | act_regs_data_and_911_enex5 ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_11_1_enexo <= and_1275_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_52 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_911_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_52 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_52 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_911_enex5 ) begin
      reg_is_start_enexo_52 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_11_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_67_ssc | act_regs_data_and_911_enex5 ) begin
      reg_act_regs_data_0_11_3_enexo_1 <= act_regs_data_and_67_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_11_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1313_tmp | act_regs_data_and_911_enex5 ) begin
      reg_act_regs_data_0_11_sva_dfm_2_1_enexo <= and_1313_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_53 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_912_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_53 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_10_1_enexo <= 1'b1;
    end
    else if ( and_1268_tmp | act_regs_data_and_912_enex5 ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_10_1_enexo <= and_1268_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_53 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_912_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_53 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_53 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_912_enex5 ) begin
      reg_is_start_enexo_53 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_10_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_66_ssc | act_regs_data_and_912_enex5 ) begin
      reg_act_regs_data_0_10_3_enexo_1 <= act_regs_data_and_66_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_10_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1311_tmp | act_regs_data_and_912_enex5 ) begin
      reg_act_regs_data_0_10_sva_dfm_2_1_enexo <= and_1311_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_9_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_127_ssc | act_regs_data_and_913_enex5 ) begin
      reg_act_regs_data_0_9_3_enexo_1 <= act_regs_data_and_127_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_54 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_913_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_54 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_54 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_913_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_54 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_0_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_64_ssc | act_regs_data_and_913_enex5 ) begin
      reg_act_regs_data_0_0_3_enexo <= act_regs_data_and_64_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_54 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_913_enex5 ) begin
      reg_is_start_enexo_54 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_9_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1309_tmp | act_regs_data_and_913_enex5 ) begin
      reg_act_regs_data_0_9_sva_dfm_2_1_enexo <= and_1309_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_55 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_914_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_55 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_8_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_78_ssc | act_regs_data_and_914_enex5 ) begin
      reg_act_regs_data_0_8_3_enexo_1 <= act_regs_data_and_78_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_55 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_914_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_55 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_55 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_914_enex5 ) begin
      reg_is_start_enexo_55 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_9_1_enexo <= 1'b1;
    end
    else if ( and_1240_tmp | act_regs_data_and_914_enex5 ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_9_1_enexo <= and_1240_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_8_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1307_tmp | act_regs_data_and_914_enex5 ) begin
      reg_act_regs_data_0_8_sva_dfm_2_1_enexo <= and_1307_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_56 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_915_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_56 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_7_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_77_ssc | act_regs_data_and_915_enex5 ) begin
      reg_act_regs_data_0_7_3_enexo_1 <= act_regs_data_and_77_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_56 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_915_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_56 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_8_1_enexo <= 1'b1;
    end
    else if ( and_1234_tmp | act_regs_data_and_915_enex5 ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_8_1_enexo <= and_1234_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_56 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_915_enex5 ) begin
      reg_is_start_enexo_56 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_7_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1305_tmp | act_regs_data_and_915_enex5 ) begin
      reg_act_regs_data_0_7_sva_dfm_2_1_enexo <= and_1305_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_7_1_enexo <= 1'b1;
    end
    else if ( and_1228_tmp | act_regs_data_and_916_enex5 ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_7_1_enexo <= and_1228_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_6_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_76_ssc | act_regs_data_and_916_enex5 ) begin
      reg_act_regs_data_0_6_3_enexo_1 <= act_regs_data_and_76_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_57 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_916_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_57 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_57 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_916_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_57 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_57 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_916_enex5 ) begin
      reg_is_start_enexo_57 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_6_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1303_tmp | act_regs_data_and_916_enex5 ) begin
      reg_act_regs_data_0_6_sva_dfm_2_1_enexo <= and_1303_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_5_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_75_ssc | act_regs_data_and_917_enex5 ) begin
      reg_act_regs_data_0_5_3_enexo_1 <= act_regs_data_and_75_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_58 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_917_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_58 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_58 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_917_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_58 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_58 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_917_enex5 ) begin
      reg_is_start_enexo_58 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_6_1_enexo <= 1'b1;
    end
    else if ( and_1289_tmp | act_regs_data_and_917_enex5 ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_6_1_enexo <= and_1289_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_5_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1301_tmp | act_regs_data_and_917_enex5 ) begin
      reg_act_regs_data_0_5_sva_dfm_2_1_enexo <= and_1301_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_59 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_918_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_59 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_59 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_918_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_59 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_4_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_74_ssc | act_regs_data_and_918_enex5 ) begin
      reg_act_regs_data_0_4_3_enexo_1 <= act_regs_data_and_74_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_59 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_918_enex5 ) begin
      reg_is_start_enexo_59 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_5_1_enexo <= 1'b1;
    end
    else if ( and_1282_tmp | act_regs_data_and_918_enex5 ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_5_1_enexo <= and_1282_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_4_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1299_tmp | act_regs_data_and_918_enex5 ) begin
      reg_act_regs_data_0_4_sva_dfm_2_1_enexo <= and_1299_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_60 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_919_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_60 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_4_1_enexo <= 1'b1;
    end
    else if ( and_1254_tmp | act_regs_data_and_919_enex5 ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_4_1_enexo <= and_1254_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_60 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_919_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_60 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_3_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_73_ssc | act_regs_data_and_919_enex5 ) begin
      reg_act_regs_data_0_3_3_enexo_1 <= act_regs_data_and_73_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_60 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_919_enex5 ) begin
      reg_is_start_enexo_60 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_3_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1297_tmp | act_regs_data_and_919_enex5 ) begin
      reg_act_regs_data_0_3_sva_dfm_2_1_enexo <= and_1297_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_61 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_920_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_61 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_3_1_enexo <= 1'b1;
    end
    else if ( and_1250_tmp | act_regs_data_and_920_enex5 ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_3_1_enexo <= and_1250_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_61 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_920_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_61 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_2_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_72_ssc | act_regs_data_and_920_enex5 ) begin
      reg_act_regs_data_0_2_3_enexo_1 <= act_regs_data_and_72_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_61 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_920_enex5 ) begin
      reg_is_start_enexo_61 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_2_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1295_tmp | act_regs_data_and_920_enex5 ) begin
      reg_act_regs_data_0_2_sva_dfm_2_1_enexo <= and_1295_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_62 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_921_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_62 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_1_1_enexo <= 1'b1;
    end
    else if ( and_1261_tmp | act_regs_data_and_921_enex5 ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_1_1_enexo <= and_1261_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_62 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_921_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_62 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_1_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_65_ssc | act_regs_data_and_921_enex5 ) begin
      reg_act_regs_data_0_1_3_enexo_1 <= act_regs_data_and_65_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_62 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_921_enex5 ) begin
      reg_is_start_enexo_62 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_1_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1293_tmp | act_regs_data_and_921_enex5 ) begin
      reg_act_regs_data_0_1_sva_dfm_2_1_enexo <= and_1293_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_0_1_enexo <= 1'b1;
    end
    else if ( and_1225_tmp | act_regs_data_and_922_enex5 ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_0_1_enexo <= and_1225_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_63 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_922_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_63 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_63 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_922_enex5 )
        begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_63 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_0_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_64_ssc | act_regs_data_and_922_enex5 ) begin
      reg_act_regs_data_0_0_3_enexo_1 <= act_regs_data_and_64_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_63 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_922_enex5 ) begin
      reg_is_start_enexo_63 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_0_sva_dfm_2_1_enexo <= 1'b1;
    end
    else if ( and_1291_tmp | act_regs_data_and_922_enex5 ) begin
      reg_act_regs_data_0_0_sva_dfm_2_1_enexo <= and_1291_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_15_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_mem_banks_read_read_data_and_16_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_15_enexo <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_14_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_mem_banks_read_read_data_and_17_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_14_enexo <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_13_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_mem_banks_read_read_data_and_18_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_13_enexo <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_12_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_mem_banks_read_read_data_and_19_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_12_enexo <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_11_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_mem_banks_read_read_data_and_20_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_11_enexo <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_10_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_mem_banks_read_read_data_and_21_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_10_enexo <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_9_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_mem_banks_read_read_data_and_22_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_9_enexo <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_8_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_mem_banks_read_read_data_and_23_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_8_enexo <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_7_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_mem_banks_read_read_data_and_24_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_7_enexo <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_6_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_mem_banks_read_read_data_and_25_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_6_enexo <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_5_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_mem_banks_read_read_data_and_26_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_5_enexo <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_4_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_mem_banks_read_read_data_and_27_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_4_enexo <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_3_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_mem_banks_read_read_data_and_28_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_3_enexo <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_2_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_mem_banks_read_read_data_and_29_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_2_enexo <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_1_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_mem_banks_read_read_data_and_30_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_1_enexo <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_mem_banks_read_read_data_and_31_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_enexo <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_15_enexo_1 <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_port_read_out_data_and_16_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_15_enexo_1 <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_31_0_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_read_data_and_16_enex5 | act_port_read_out_data_and_16_enex5
        ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_31_0_enexo <= act_mem_banks_read_read_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_CheckStart_start_reg_enexo <= 1'b1;
    end
    else if ( ActUnit_CheckStart_start_reg_and_tmp | act_port_read_out_data_and_16_enex5
        ) begin
      reg_ActUnit_CheckStart_start_reg_enexo <= ActUnit_CheckStart_start_reg_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_63_32_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_read_data_and_17_enex5 | act_port_read_out_data_and_17_enex5
        ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_63_32_enexo <= act_mem_banks_read_read_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_CheckStart_start_reg_enexo_1 <= 1'b1;
    end
    else if ( ActUnit_CheckStart_start_reg_and_tmp | act_port_read_out_data_and_17_enex5
        ) begin
      reg_ActUnit_CheckStart_start_reg_enexo_1 <= ActUnit_CheckStart_start_reg_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_14_enexo_1 <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_port_read_out_data_and_17_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_14_enexo_1 <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_95_64_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_read_data_and_18_enex5 | act_port_read_out_data_and_18_enex5
        ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_95_64_enexo <= act_mem_banks_read_read_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_CheckStart_start_reg_enexo_2 <= 1'b1;
    end
    else if ( ActUnit_CheckStart_start_reg_and_tmp | act_port_read_out_data_and_18_enex5
        ) begin
      reg_ActUnit_CheckStart_start_reg_enexo_2 <= ActUnit_CheckStart_start_reg_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_13_enexo_1 <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_port_read_out_data_and_18_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_13_enexo_1 <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_CheckStart_start_reg_enexo_3 <= 1'b1;
    end
    else if ( ActUnit_CheckStart_start_reg_and_tmp | act_port_read_out_data_and_19_enex5
        ) begin
      reg_ActUnit_CheckStart_start_reg_enexo_3 <= ActUnit_CheckStart_start_reg_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_12_enexo_1 <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_port_read_out_data_and_19_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_12_enexo_1 <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_127_96_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_read_data_and_19_enex5 | act_port_read_out_data_and_19_enex5
        ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_127_96_enexo <= act_mem_banks_read_read_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_11_enexo_1 <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_port_read_out_data_and_20_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_11_enexo_1 <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_CheckStart_start_reg_enexo_4 <= 1'b1;
    end
    else if ( ActUnit_CheckStart_start_reg_and_tmp | act_port_read_out_data_and_20_enex5
        ) begin
      reg_ActUnit_CheckStart_start_reg_enexo_4 <= ActUnit_CheckStart_start_reg_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_159_128_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_read_data_and_20_enex5 | act_port_read_out_data_and_20_enex5
        ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_159_128_enexo <= act_mem_banks_read_read_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_10_enexo_1 <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_port_read_out_data_and_21_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_10_enexo_1 <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_191_160_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_read_data_and_21_enex5 | act_port_read_out_data_and_21_enex5
        ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_191_160_enexo <= act_mem_banks_read_read_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_CheckStart_start_reg_enexo_5 <= 1'b1;
    end
    else if ( ActUnit_CheckStart_start_reg_and_tmp | act_port_read_out_data_and_21_enex5
        ) begin
      reg_ActUnit_CheckStart_start_reg_enexo_5 <= ActUnit_CheckStart_start_reg_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_9_enexo_1 <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_port_read_out_data_and_22_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_9_enexo_1 <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_223_192_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_read_data_and_22_enex5 | act_port_read_out_data_and_22_enex5
        ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_223_192_enexo <= act_mem_banks_read_read_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_CheckStart_start_reg_enexo_6 <= 1'b1;
    end
    else if ( ActUnit_CheckStart_start_reg_and_tmp | act_port_read_out_data_and_22_enex5
        ) begin
      reg_ActUnit_CheckStart_start_reg_enexo_6 <= ActUnit_CheckStart_start_reg_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_8_enexo_1 <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_port_read_out_data_and_23_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_8_enexo_1 <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_CheckStart_start_reg_enexo_7 <= 1'b1;
    end
    else if ( ActUnit_CheckStart_start_reg_and_tmp | act_port_read_out_data_and_23_enex5
        ) begin
      reg_ActUnit_CheckStart_start_reg_enexo_7 <= ActUnit_CheckStart_start_reg_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_255_224_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_read_data_and_23_enex5 | act_port_read_out_data_and_23_enex5
        ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_255_224_enexo <= act_mem_banks_read_read_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_287_256_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_read_data_and_24_enex5 | act_port_read_out_data_and_24_enex5
        ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_287_256_enexo <= act_mem_banks_read_read_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_7_enexo_1 <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_port_read_out_data_and_24_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_7_enexo_1 <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_CheckStart_start_reg_enexo_8 <= 1'b1;
    end
    else if ( ActUnit_CheckStart_start_reg_and_tmp | act_port_read_out_data_and_24_enex5
        ) begin
      reg_ActUnit_CheckStart_start_reg_enexo_8 <= ActUnit_CheckStart_start_reg_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_6_enexo_1 <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_port_read_out_data_and_25_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_6_enexo_1 <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_319_288_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_read_data_and_25_enex5 | act_port_read_out_data_and_25_enex5
        ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_319_288_enexo <= act_mem_banks_read_read_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_CheckStart_start_reg_enexo_9 <= 1'b1;
    end
    else if ( ActUnit_CheckStart_start_reg_and_tmp | act_port_read_out_data_and_25_enex5
        ) begin
      reg_ActUnit_CheckStart_start_reg_enexo_9 <= ActUnit_CheckStart_start_reg_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_5_enexo_1 <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_port_read_out_data_and_26_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_5_enexo_1 <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_CheckStart_start_reg_enexo_10 <= 1'b1;
    end
    else if ( ActUnit_CheckStart_start_reg_and_tmp | act_port_read_out_data_and_26_enex5
        ) begin
      reg_ActUnit_CheckStart_start_reg_enexo_10 <= ActUnit_CheckStart_start_reg_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_351_320_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_read_data_and_26_enex5 | act_port_read_out_data_and_26_enex5
        ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_351_320_enexo <= act_mem_banks_read_read_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_4_enexo_1 <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_port_read_out_data_and_27_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_4_enexo_1 <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_383_352_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_read_data_and_27_enex5 | act_port_read_out_data_and_27_enex5
        ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_383_352_enexo <= act_mem_banks_read_read_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_CheckStart_start_reg_enexo_11 <= 1'b1;
    end
    else if ( ActUnit_CheckStart_start_reg_and_tmp | act_port_read_out_data_and_27_enex5
        ) begin
      reg_ActUnit_CheckStart_start_reg_enexo_11 <= ActUnit_CheckStart_start_reg_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_415_384_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_read_data_and_28_enex5 | act_port_read_out_data_and_28_enex5
        ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_415_384_enexo <= act_mem_banks_read_read_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_3_enexo_1 <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_port_read_out_data_and_28_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_3_enexo_1 <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_CheckStart_start_reg_enexo_12 <= 1'b1;
    end
    else if ( ActUnit_CheckStart_start_reg_and_tmp | act_port_read_out_data_and_28_enex5
        ) begin
      reg_ActUnit_CheckStart_start_reg_enexo_12 <= ActUnit_CheckStart_start_reg_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_447_416_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_read_data_and_29_enex5 | act_port_read_out_data_and_29_enex5
        ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_447_416_enexo <= act_mem_banks_read_read_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_2_enexo_1 <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_port_read_out_data_and_29_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_2_enexo_1 <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_CheckStart_start_reg_enexo_13 <= 1'b1;
    end
    else if ( ActUnit_CheckStart_start_reg_and_tmp | act_port_read_out_data_and_29_enex5
        ) begin
      reg_ActUnit_CheckStart_start_reg_enexo_13 <= ActUnit_CheckStart_start_reg_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_479_448_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_read_data_and_30_enex5 | act_port_read_out_data_and_30_enex5
        ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_479_448_enexo <= act_mem_banks_read_read_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_1_enexo_1 <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_port_read_out_data_and_30_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_1_enexo_1 <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_CheckStart_start_reg_enexo_14 <= 1'b1;
    end
    else if ( ActUnit_CheckStart_start_reg_and_tmp | act_port_read_out_data_and_30_enex5
        ) begin
      reg_ActUnit_CheckStart_start_reg_enexo_14 <= ActUnit_CheckStart_start_reg_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_enexo_1 <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_port_read_out_data_and_31_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_enexo_1 <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_CheckStart_start_reg_enexo_15 <= 1'b1;
    end
    else if ( ActUnit_CheckStart_start_reg_and_tmp | act_port_read_out_data_and_31_enex5
        ) begin
      reg_ActUnit_CheckStart_start_reg_enexo_15 <= ActUnit_CheckStart_start_reg_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_511_480_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_read_data_and_31_enex5 | act_port_read_out_data_and_31_enex5
        ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_511_480_enexo <= act_mem_banks_read_read_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_37_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_37_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_15_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_891_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_37_enex5
        ) begin
      reg_act_regs_data_1_15_2_enexo <= act_regs_data_and_891_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_15_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_875_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_37_enex5
        ) begin
      reg_act_regs_data_2_15_2_enexo <= act_regs_data_and_875_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_15_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_907_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_37_enex5
        ) begin
      reg_act_regs_data_0_15_2_enexo <= act_regs_data_and_907_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_37_enex5
        ) begin
      reg_act_config_inst_counter_enexo <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_15_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_859_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_37_enex5
        ) begin
      reg_act_regs_data_3_15_2_enexo <= act_regs_data_and_859_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_1 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_38_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_1 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_1 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_38_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_1 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_14_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_860_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_38_enex5
        ) begin
      reg_act_regs_data_3_14_2_enexo <= act_regs_data_and_860_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_14_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_908_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_38_enex5
        ) begin
      reg_act_regs_data_0_14_2_enexo <= act_regs_data_and_908_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_14_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_892_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_38_enex5
        ) begin
      reg_act_regs_data_1_14_2_enexo <= act_regs_data_and_892_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_14_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_876_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_38_enex5
        ) begin
      reg_act_regs_data_2_14_2_enexo <= act_regs_data_and_876_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_1 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_38_enex5
        ) begin
      reg_act_config_inst_counter_enexo_1 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_2 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_39_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_2 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_2 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_39_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_2 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_13_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_893_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_39_enex5
        ) begin
      reg_act_regs_data_1_13_2_enexo <= act_regs_data_and_893_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_13_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_909_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_39_enex5
        ) begin
      reg_act_regs_data_0_13_2_enexo <= act_regs_data_and_909_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_13_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_861_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_39_enex5
        ) begin
      reg_act_regs_data_3_13_2_enexo <= act_regs_data_and_861_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_13_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_877_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_39_enex5
        ) begin
      reg_act_regs_data_2_13_2_enexo <= act_regs_data_and_877_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_2 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_39_enex5
        ) begin
      reg_act_config_inst_counter_enexo_2 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_3 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_40_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_3 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_3 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_40_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_3 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_12_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_894_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_40_enex5
        ) begin
      reg_act_regs_data_1_12_2_enexo <= act_regs_data_and_894_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_12_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_878_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_40_enex5
        ) begin
      reg_act_regs_data_2_12_2_enexo <= act_regs_data_and_878_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_12_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_910_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_40_enex5
        ) begin
      reg_act_regs_data_0_12_2_enexo <= act_regs_data_and_910_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_12_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_862_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_40_enex5
        ) begin
      reg_act_regs_data_3_12_2_enexo <= act_regs_data_and_862_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_3 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_40_enex5
        ) begin
      reg_act_config_inst_counter_enexo_3 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_4 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_41_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_4 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_4 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_41_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_4 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_11_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_879_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_41_enex5
        ) begin
      reg_act_regs_data_2_11_2_enexo <= act_regs_data_and_879_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_11_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_863_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_41_enex5
        ) begin
      reg_act_regs_data_3_11_2_enexo <= act_regs_data_and_863_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_11_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_895_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_41_enex5
        ) begin
      reg_act_regs_data_1_11_2_enexo <= act_regs_data_and_895_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_11_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_911_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_41_enex5
        ) begin
      reg_act_regs_data_0_11_2_enexo <= act_regs_data_and_911_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_4 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_41_enex5
        ) begin
      reg_act_config_inst_counter_enexo_4 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_5 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_42_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_5 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_5 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_42_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_5 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_10_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_912_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_42_enex5
        ) begin
      reg_act_regs_data_0_10_2_enexo <= act_regs_data_and_912_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_10_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_896_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_42_enex5
        ) begin
      reg_act_regs_data_1_10_2_enexo <= act_regs_data_and_896_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_10_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_880_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_42_enex5
        ) begin
      reg_act_regs_data_2_10_2_enexo <= act_regs_data_and_880_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_10_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_864_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_42_enex5
        ) begin
      reg_act_regs_data_3_10_2_enexo <= act_regs_data_and_864_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_5 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_42_enex5
        ) begin
      reg_act_config_inst_counter_enexo_5 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_6 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_43_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_6 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_6 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_43_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_6 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_9_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_897_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_43_enex5
        ) begin
      reg_act_regs_data_1_9_2_enexo <= act_regs_data_and_897_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_9_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_913_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_43_enex5
        ) begin
      reg_act_regs_data_0_9_2_enexo <= act_regs_data_and_913_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_9_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_881_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_43_enex5
        ) begin
      reg_act_regs_data_2_9_2_enexo <= act_regs_data_and_881_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_9_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_865_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_43_enex5
        ) begin
      reg_act_regs_data_3_9_2_enexo <= act_regs_data_and_865_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_6 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_43_enex5
        ) begin
      reg_act_config_inst_counter_enexo_6 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_7 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_44_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_7 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_7 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_44_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_7 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_8_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_866_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_44_enex5
        ) begin
      reg_act_regs_data_3_8_2_enexo <= act_regs_data_and_866_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_8_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_898_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_44_enex5
        ) begin
      reg_act_regs_data_1_8_2_enexo <= act_regs_data_and_898_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_8_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_914_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_44_enex5
        ) begin
      reg_act_regs_data_0_8_2_enexo <= act_regs_data_and_914_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_8_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_882_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_44_enex5
        ) begin
      reg_act_regs_data_2_8_2_enexo <= act_regs_data_and_882_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_7 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_44_enex5
        ) begin
      reg_act_config_inst_counter_enexo_7 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_8 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_45_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_8 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_8 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_45_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_8 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_7_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_883_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_45_enex5
        ) begin
      reg_act_regs_data_2_7_2_enexo <= act_regs_data_and_883_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_7_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_899_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_45_enex5
        ) begin
      reg_act_regs_data_1_7_2_enexo <= act_regs_data_and_899_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_7_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_915_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_45_enex5
        ) begin
      reg_act_regs_data_0_7_2_enexo <= act_regs_data_and_915_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_7_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_867_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_45_enex5
        ) begin
      reg_act_regs_data_3_7_2_enexo <= act_regs_data_and_867_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_8 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_45_enex5
        ) begin
      reg_act_config_inst_counter_enexo_8 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_9 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_46_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_9 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_9 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_46_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_9 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_6_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_868_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_46_enex5
        ) begin
      reg_act_regs_data_3_6_2_enexo <= act_regs_data_and_868_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_6_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_900_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_46_enex5
        ) begin
      reg_act_regs_data_1_6_2_enexo <= act_regs_data_and_900_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_6_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_916_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_46_enex5
        ) begin
      reg_act_regs_data_0_6_2_enexo <= act_regs_data_and_916_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_6_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_884_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_46_enex5
        ) begin
      reg_act_regs_data_2_6_2_enexo <= act_regs_data_and_884_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_9 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_46_enex5
        ) begin
      reg_act_config_inst_counter_enexo_9 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_10 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_47_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_10 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_10 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_47_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_10 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_5_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_917_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_47_enex5
        ) begin
      reg_act_regs_data_0_5_2_enexo <= act_regs_data_and_917_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_5_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_885_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_47_enex5
        ) begin
      reg_act_regs_data_2_5_2_enexo <= act_regs_data_and_885_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_5_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_869_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_47_enex5
        ) begin
      reg_act_regs_data_3_5_2_enexo <= act_regs_data_and_869_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_5_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_901_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_47_enex5
        ) begin
      reg_act_regs_data_1_5_2_enexo <= act_regs_data_and_901_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_10 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_47_enex5
        ) begin
      reg_act_config_inst_counter_enexo_10 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_11 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_48_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_11 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_11 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_48_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_11 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_4_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_886_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_48_enex5
        ) begin
      reg_act_regs_data_2_4_2_enexo <= act_regs_data_and_886_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_4_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_870_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_48_enex5
        ) begin
      reg_act_regs_data_3_4_2_enexo <= act_regs_data_and_870_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_4_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_902_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_48_enex5
        ) begin
      reg_act_regs_data_1_4_2_enexo <= act_regs_data_and_902_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_4_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_918_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_48_enex5
        ) begin
      reg_act_regs_data_0_4_2_enexo <= act_regs_data_and_918_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_11 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_48_enex5
        ) begin
      reg_act_config_inst_counter_enexo_11 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_12 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_49_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_12 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_12 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_49_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_12 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_3_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_887_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_49_enex5
        ) begin
      reg_act_regs_data_2_3_2_enexo <= act_regs_data_and_887_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_3_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_871_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_49_enex5
        ) begin
      reg_act_regs_data_3_3_2_enexo <= act_regs_data_and_871_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_3_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_903_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_49_enex5
        ) begin
      reg_act_regs_data_1_3_2_enexo <= act_regs_data_and_903_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_3_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_919_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_49_enex5
        ) begin
      reg_act_regs_data_0_3_2_enexo <= act_regs_data_and_919_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_12 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_49_enex5
        ) begin
      reg_act_config_inst_counter_enexo_12 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_13 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_50_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_13 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_13 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_50_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_13 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_2_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_920_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_50_enex5
        ) begin
      reg_act_regs_data_0_2_2_enexo <= act_regs_data_and_920_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_2_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_888_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_50_enex5
        ) begin
      reg_act_regs_data_2_2_2_enexo <= act_regs_data_and_888_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_2_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_904_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_50_enex5
        ) begin
      reg_act_regs_data_1_2_2_enexo <= act_regs_data_and_904_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_2_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_872_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_50_enex5
        ) begin
      reg_act_regs_data_3_2_2_enexo <= act_regs_data_and_872_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_13 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_50_enex5
        ) begin
      reg_act_config_inst_counter_enexo_13 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_14 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_51_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_14 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_14 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_51_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_14 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_1_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_905_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_51_enex5
        ) begin
      reg_act_regs_data_1_1_2_enexo <= act_regs_data_and_905_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_1_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_873_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_51_enex5
        ) begin
      reg_act_regs_data_3_1_2_enexo <= act_regs_data_and_873_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_1_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_921_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_51_enex5
        ) begin
      reg_act_regs_data_0_1_2_enexo <= act_regs_data_and_921_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_1_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_889_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_51_enex5
        ) begin
      reg_act_regs_data_2_1_2_enexo <= act_regs_data_and_889_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_14 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_51_enex5
        ) begin
      reg_act_config_inst_counter_enexo_14 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_15 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_52_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_15 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_15 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_52_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_15 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_0_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_890_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_52_enex5
        ) begin
      reg_act_regs_data_2_0_2_enexo <= act_regs_data_and_890_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_0_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_874_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_52_enex5
        ) begin
      reg_act_regs_data_3_0_2_enexo <= act_regs_data_and_874_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_0_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_906_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_52_enex5
        ) begin
      reg_act_regs_data_1_0_2_enexo <= act_regs_data_and_906_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_0_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_922_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_52_enex5
        ) begin
      reg_act_regs_data_0_0_2_enexo <= act_regs_data_and_922_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_15 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_52_enex5
        ) begin
      reg_act_config_inst_counter_enexo_15 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_16 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_31_enex5 ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_16 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_16 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_31_enex5 ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_16 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_15_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_cse | Relu_for_y_qelse_and_31_enex5 ) begin
      reg_act_regs_data_3_15_enexo <= act_regs_data_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_15_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_891_enex5 | Relu_for_y_qelse_and_31_enex5 ) begin
      reg_act_regs_data_1_15_2_enexo_1 <= act_regs_data_and_891_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_15_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_875_enex5 | Relu_for_y_qelse_and_31_enex5 ) begin
      reg_act_regs_data_2_15_2_enexo_1 <= act_regs_data_and_875_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_15_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_907_enex5 | Relu_for_y_qelse_and_31_enex5 ) begin
      reg_act_regs_data_0_15_2_enexo_1 <= act_regs_data_and_907_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_16 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_31_enex5 ) begin
      reg_act_config_inst_counter_enexo_16 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_15_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_859_enex5 | Relu_for_y_qelse_and_31_enex5 ) begin
      reg_act_regs_data_3_15_2_enexo_1 <= act_regs_data_and_859_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_17 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_32_enex5 ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_17 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_17 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_32_enex5 ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_17 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_14_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_cse | Relu_for_y_qelse_and_32_enex5 ) begin
      reg_act_regs_data_1_14_enexo <= act_regs_data_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_14_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_860_enex5 | Relu_for_y_qelse_and_32_enex5 ) begin
      reg_act_regs_data_3_14_2_enexo_1 <= act_regs_data_and_860_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_14_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_908_enex5 | Relu_for_y_qelse_and_32_enex5 ) begin
      reg_act_regs_data_0_14_2_enexo_1 <= act_regs_data_and_908_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_14_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_892_enex5 | Relu_for_y_qelse_and_32_enex5 ) begin
      reg_act_regs_data_1_14_2_enexo_1 <= act_regs_data_and_892_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_14_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_876_enex5 | Relu_for_y_qelse_and_32_enex5 ) begin
      reg_act_regs_data_2_14_2_enexo_1 <= act_regs_data_and_876_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_17 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_32_enex5 ) begin
      reg_act_config_inst_counter_enexo_17 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_18 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_33_enex5 ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_18 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_18 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_33_enex5 ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_18 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_13_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_893_enex5 | Relu_for_y_qelse_and_33_enex5 ) begin
      reg_act_regs_data_1_13_2_enexo_1 <= act_regs_data_and_893_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_13_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_cse | Relu_for_y_qelse_and_33_enex5 ) begin
      reg_act_regs_data_1_13_enexo <= act_regs_data_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_13_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_909_enex5 | Relu_for_y_qelse_and_33_enex5 ) begin
      reg_act_regs_data_0_13_2_enexo_1 <= act_regs_data_and_909_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_13_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_861_enex5 | Relu_for_y_qelse_and_33_enex5 ) begin
      reg_act_regs_data_3_13_2_enexo_1 <= act_regs_data_and_861_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_13_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_877_enex5 | Relu_for_y_qelse_and_33_enex5 ) begin
      reg_act_regs_data_2_13_2_enexo_1 <= act_regs_data_and_877_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_18 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_33_enex5 ) begin
      reg_act_config_inst_counter_enexo_18 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_19 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_34_enex5 ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_19 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_19 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_34_enex5 ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_19 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_12_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_cse | Relu_for_y_qelse_and_34_enex5 ) begin
      reg_act_regs_data_1_12_enexo <= act_regs_data_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_12_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_894_enex5 | Relu_for_y_qelse_and_34_enex5 ) begin
      reg_act_regs_data_1_12_2_enexo_1 <= act_regs_data_and_894_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_12_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_878_enex5 | Relu_for_y_qelse_and_34_enex5 ) begin
      reg_act_regs_data_2_12_2_enexo_1 <= act_regs_data_and_878_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_12_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_910_enex5 | Relu_for_y_qelse_and_34_enex5 ) begin
      reg_act_regs_data_0_12_2_enexo_1 <= act_regs_data_and_910_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_12_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_862_enex5 | Relu_for_y_qelse_and_34_enex5 ) begin
      reg_act_regs_data_3_12_2_enexo_1 <= act_regs_data_and_862_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_19 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_34_enex5 ) begin
      reg_act_config_inst_counter_enexo_19 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_20 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_35_enex5 ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_20 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_20 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_35_enex5 ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_20 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_11_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_cse | Relu_for_y_qelse_and_35_enex5 ) begin
      reg_act_regs_data_1_11_enexo <= act_regs_data_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_11_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_879_enex5 | Relu_for_y_qelse_and_35_enex5 ) begin
      reg_act_regs_data_2_11_2_enexo_1 <= act_regs_data_and_879_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_11_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_863_enex5 | Relu_for_y_qelse_and_35_enex5 ) begin
      reg_act_regs_data_3_11_2_enexo_1 <= act_regs_data_and_863_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_11_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_895_enex5 | Relu_for_y_qelse_and_35_enex5 ) begin
      reg_act_regs_data_1_11_2_enexo_1 <= act_regs_data_and_895_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_11_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_911_enex5 | Relu_for_y_qelse_and_35_enex5 ) begin
      reg_act_regs_data_0_11_2_enexo_1 <= act_regs_data_and_911_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_20 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_35_enex5 ) begin
      reg_act_config_inst_counter_enexo_20 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_21 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_36_enex5 ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_21 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_21 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_36_enex5 ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_21 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_10_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_912_enex5 | Relu_for_y_qelse_and_36_enex5 ) begin
      reg_act_regs_data_0_10_2_enexo_1 <= act_regs_data_and_912_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_10_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_cse | Relu_for_y_qelse_and_36_enex5 ) begin
      reg_act_regs_data_2_10_enexo <= act_regs_data_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_10_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_896_enex5 | Relu_for_y_qelse_and_36_enex5 ) begin
      reg_act_regs_data_1_10_2_enexo_1 <= act_regs_data_and_896_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_10_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_880_enex5 | Relu_for_y_qelse_and_36_enex5 ) begin
      reg_act_regs_data_2_10_2_enexo_1 <= act_regs_data_and_880_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_10_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_864_enex5 | Relu_for_y_qelse_and_36_enex5 ) begin
      reg_act_regs_data_3_10_2_enexo_1 <= act_regs_data_and_864_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_21 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_36_enex5 ) begin
      reg_act_config_inst_counter_enexo_21 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_22 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_37_enex5 ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_22 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_22 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_37_enex5 ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_22 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_9_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_cse | Relu_for_y_qelse_and_37_enex5 ) begin
      reg_act_regs_data_0_9_enexo <= act_regs_data_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_9_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_897_enex5 | Relu_for_y_qelse_and_37_enex5 ) begin
      reg_act_regs_data_1_9_2_enexo_1 <= act_regs_data_and_897_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_9_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_913_enex5 | Relu_for_y_qelse_and_37_enex5 ) begin
      reg_act_regs_data_0_9_2_enexo_1 <= act_regs_data_and_913_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_9_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_881_enex5 | Relu_for_y_qelse_and_37_enex5 ) begin
      reg_act_regs_data_2_9_2_enexo_1 <= act_regs_data_and_881_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_9_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_865_enex5 | Relu_for_y_qelse_and_37_enex5 ) begin
      reg_act_regs_data_3_9_2_enexo_1 <= act_regs_data_and_865_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_22 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_37_enex5 ) begin
      reg_act_config_inst_counter_enexo_22 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_23 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_38_enex5 ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_23 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_23 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_38_enex5 ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_23 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_8_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_cse | Relu_for_y_qelse_and_38_enex5 ) begin
      reg_act_regs_data_0_8_enexo <= act_regs_data_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_8_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_866_enex5 | Relu_for_y_qelse_and_38_enex5 ) begin
      reg_act_regs_data_3_8_2_enexo_1 <= act_regs_data_and_866_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_8_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_898_enex5 | Relu_for_y_qelse_and_38_enex5 ) begin
      reg_act_regs_data_1_8_2_enexo_1 <= act_regs_data_and_898_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_8_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_914_enex5 | Relu_for_y_qelse_and_38_enex5 ) begin
      reg_act_regs_data_0_8_2_enexo_1 <= act_regs_data_and_914_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_8_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_882_enex5 | Relu_for_y_qelse_and_38_enex5 ) begin
      reg_act_regs_data_2_8_2_enexo_1 <= act_regs_data_and_882_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_23 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_38_enex5 ) begin
      reg_act_config_inst_counter_enexo_23 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_24 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_39_enex5 ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_24 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_24 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_39_enex5 ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_24 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_7_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_883_enex5 | Relu_for_y_qelse_and_39_enex5 ) begin
      reg_act_regs_data_2_7_2_enexo_1 <= act_regs_data_and_883_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_7_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_cse | Relu_for_y_qelse_and_39_enex5 ) begin
      reg_act_regs_data_1_7_enexo <= act_regs_data_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_7_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_899_enex5 | Relu_for_y_qelse_and_39_enex5 ) begin
      reg_act_regs_data_1_7_2_enexo_1 <= act_regs_data_and_899_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_7_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_915_enex5 | Relu_for_y_qelse_and_39_enex5 ) begin
      reg_act_regs_data_0_7_2_enexo_1 <= act_regs_data_and_915_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_7_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_867_enex5 | Relu_for_y_qelse_and_39_enex5 ) begin
      reg_act_regs_data_3_7_2_enexo_1 <= act_regs_data_and_867_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_24 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_39_enex5 ) begin
      reg_act_config_inst_counter_enexo_24 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_25 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_40_enex5 ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_25 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_25 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_40_enex5 ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_25 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_6_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_cse | Relu_for_y_qelse_and_40_enex5 ) begin
      reg_act_regs_data_2_6_enexo <= act_regs_data_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_6_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_868_enex5 | Relu_for_y_qelse_and_40_enex5 ) begin
      reg_act_regs_data_3_6_2_enexo_1 <= act_regs_data_and_868_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_6_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_900_enex5 | Relu_for_y_qelse_and_40_enex5 ) begin
      reg_act_regs_data_1_6_2_enexo_1 <= act_regs_data_and_900_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_6_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_916_enex5 | Relu_for_y_qelse_and_40_enex5 ) begin
      reg_act_regs_data_0_6_2_enexo_1 <= act_regs_data_and_916_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_6_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_884_enex5 | Relu_for_y_qelse_and_40_enex5 ) begin
      reg_act_regs_data_2_6_2_enexo_1 <= act_regs_data_and_884_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_25 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_40_enex5 ) begin
      reg_act_config_inst_counter_enexo_25 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_26 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_41_enex5 ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_26 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_26 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_41_enex5 ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_26 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_5_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_917_enex5 | Relu_for_y_qelse_and_41_enex5 ) begin
      reg_act_regs_data_0_5_2_enexo_1 <= act_regs_data_and_917_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_5_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_885_enex5 | Relu_for_y_qelse_and_41_enex5 ) begin
      reg_act_regs_data_2_5_2_enexo_1 <= act_regs_data_and_885_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_5_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_cse | Relu_for_y_qelse_and_41_enex5 ) begin
      reg_act_regs_data_3_5_enexo <= act_regs_data_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_5_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_869_enex5 | Relu_for_y_qelse_and_41_enex5 ) begin
      reg_act_regs_data_3_5_2_enexo_1 <= act_regs_data_and_869_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_5_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_901_enex5 | Relu_for_y_qelse_and_41_enex5 ) begin
      reg_act_regs_data_1_5_2_enexo_1 <= act_regs_data_and_901_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_26 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_41_enex5 ) begin
      reg_act_config_inst_counter_enexo_26 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_27 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_42_enex5 ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_27 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_27 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_42_enex5 ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_27 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_4_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_cse | Relu_for_y_qelse_and_42_enex5 ) begin
      reg_act_regs_data_1_4_enexo <= act_regs_data_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_4_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_886_enex5 | Relu_for_y_qelse_and_42_enex5 ) begin
      reg_act_regs_data_2_4_2_enexo_1 <= act_regs_data_and_886_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_4_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_870_enex5 | Relu_for_y_qelse_and_42_enex5 ) begin
      reg_act_regs_data_3_4_2_enexo_1 <= act_regs_data_and_870_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_4_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_902_enex5 | Relu_for_y_qelse_and_42_enex5 ) begin
      reg_act_regs_data_1_4_2_enexo_1 <= act_regs_data_and_902_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_4_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_918_enex5 | Relu_for_y_qelse_and_42_enex5 ) begin
      reg_act_regs_data_0_4_2_enexo_1 <= act_regs_data_and_918_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_27 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_42_enex5 ) begin
      reg_act_config_inst_counter_enexo_27 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_28 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_43_enex5 ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_28 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_28 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_43_enex5 ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_28 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_cse | Relu_for_y_qelse_and_43_enex5 ) begin
      reg_act_regs_data_0_3_enexo <= act_regs_data_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_3_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_887_enex5 | Relu_for_y_qelse_and_43_enex5 ) begin
      reg_act_regs_data_2_3_2_enexo_1 <= act_regs_data_and_887_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_3_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_871_enex5 | Relu_for_y_qelse_and_43_enex5 ) begin
      reg_act_regs_data_3_3_2_enexo_1 <= act_regs_data_and_871_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_3_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_903_enex5 | Relu_for_y_qelse_and_43_enex5 ) begin
      reg_act_regs_data_1_3_2_enexo_1 <= act_regs_data_and_903_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_3_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_919_enex5 | Relu_for_y_qelse_and_43_enex5 ) begin
      reg_act_regs_data_0_3_2_enexo_1 <= act_regs_data_and_919_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_28 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_43_enex5 ) begin
      reg_act_config_inst_counter_enexo_28 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_29 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_44_enex5 ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_29 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_29 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_44_enex5 ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_29 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_cse | Relu_for_y_qelse_and_44_enex5 ) begin
      reg_act_regs_data_1_2_enexo <= act_regs_data_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_2_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_920_enex5 | Relu_for_y_qelse_and_44_enex5 ) begin
      reg_act_regs_data_0_2_2_enexo_1 <= act_regs_data_and_920_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_2_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_888_enex5 | Relu_for_y_qelse_and_44_enex5 ) begin
      reg_act_regs_data_2_2_2_enexo_1 <= act_regs_data_and_888_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_2_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_904_enex5 | Relu_for_y_qelse_and_44_enex5 ) begin
      reg_act_regs_data_1_2_2_enexo_1 <= act_regs_data_and_904_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_2_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_872_enex5 | Relu_for_y_qelse_and_44_enex5 ) begin
      reg_act_regs_data_3_2_2_enexo_1 <= act_regs_data_and_872_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_29 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_44_enex5 ) begin
      reg_act_config_inst_counter_enexo_29 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_30 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_45_enex5 ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_30 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_30 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_45_enex5 ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_30 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_cse | Relu_for_y_qelse_and_45_enex5 ) begin
      reg_act_regs_data_0_1_enexo <= act_regs_data_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_1_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_905_enex5 | Relu_for_y_qelse_and_45_enex5 ) begin
      reg_act_regs_data_1_1_2_enexo_1 <= act_regs_data_and_905_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_1_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_873_enex5 | Relu_for_y_qelse_and_45_enex5 ) begin
      reg_act_regs_data_3_1_2_enexo_1 <= act_regs_data_and_873_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_1_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_921_enex5 | Relu_for_y_qelse_and_45_enex5 ) begin
      reg_act_regs_data_0_1_2_enexo_1 <= act_regs_data_and_921_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_1_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_889_enex5 | Relu_for_y_qelse_and_45_enex5 ) begin
      reg_act_regs_data_2_1_2_enexo_1 <= act_regs_data_and_889_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_30 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_45_enex5 ) begin
      reg_act_config_inst_counter_enexo_30 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_31 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_46_enex5 ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_31 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_31 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_46_enex5 ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_31 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_cse | Relu_for_y_qelse_and_46_enex5 ) begin
      reg_act_regs_data_2_0_enexo <= act_regs_data_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_0_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_890_enex5 | Relu_for_y_qelse_and_46_enex5 ) begin
      reg_act_regs_data_2_0_2_enexo_1 <= act_regs_data_and_890_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_0_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_874_enex5 | Relu_for_y_qelse_and_46_enex5 ) begin
      reg_act_regs_data_3_0_2_enexo_1 <= act_regs_data_and_874_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_0_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_906_enex5 | Relu_for_y_qelse_and_46_enex5 ) begin
      reg_act_regs_data_1_0_2_enexo_1 <= act_regs_data_and_906_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_0_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_922_enex5 | Relu_for_y_qelse_and_46_enex5 ) begin
      reg_act_regs_data_0_0_2_enexo_1 <= act_regs_data_and_922_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_31 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_46_enex5 ) begin
      reg_act_config_inst_counter_enexo_31 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_32 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_15_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_32 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_32 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_15_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_32 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_2_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_920_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_15_enex5
        ) begin
      reg_act_regs_data_0_2_2_enexo_2 <= act_regs_data_and_920_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_2_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_888_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_15_enex5
        ) begin
      reg_act_regs_data_2_2_2_enexo_2 <= act_regs_data_and_888_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_2_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_904_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_15_enex5
        ) begin
      reg_act_regs_data_1_2_2_enexo_2 <= act_regs_data_and_904_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_2_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_872_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_15_enex5
        ) begin
      reg_act_regs_data_3_2_2_enexo_2 <= act_regs_data_and_872_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_32 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_15_enex5
        ) begin
      reg_act_config_inst_counter_enexo_32 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_33 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_16_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_33 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_33 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_16_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_33 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_3_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_887_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_16_enex5
        ) begin
      reg_act_regs_data_2_3_2_enexo_2 <= act_regs_data_and_887_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_3_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_871_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_16_enex5
        ) begin
      reg_act_regs_data_3_3_2_enexo_2 <= act_regs_data_and_871_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_3_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_903_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_16_enex5
        ) begin
      reg_act_regs_data_1_3_2_enexo_2 <= act_regs_data_and_903_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_3_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_919_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_16_enex5
        ) begin
      reg_act_regs_data_0_3_2_enexo_2 <= act_regs_data_and_919_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_33 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_16_enex5
        ) begin
      reg_act_config_inst_counter_enexo_33 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_34 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | ActUnit_RunInst_switch_lp_and_815_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_34 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_34 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | ActUnit_RunInst_switch_lp_and_815_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_34 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_0_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_890_enex5 | ActUnit_RunInst_switch_lp_and_815_enex5
        ) begin
      reg_act_regs_data_2_0_2_enexo_2 <= act_regs_data_and_890_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_0_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_874_enex5 | ActUnit_RunInst_switch_lp_and_815_enex5
        ) begin
      reg_act_regs_data_3_0_2_enexo_2 <= act_regs_data_and_874_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_0_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_906_enex5 | ActUnit_RunInst_switch_lp_and_815_enex5
        ) begin
      reg_act_regs_data_1_0_2_enexo_2 <= act_regs_data_and_906_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_0_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_922_enex5 | ActUnit_RunInst_switch_lp_and_815_enex5
        ) begin
      reg_act_regs_data_0_0_2_enexo_2 <= act_regs_data_and_922_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_34 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | ActUnit_RunInst_switch_lp_and_815_enex5
        ) begin
      reg_act_config_inst_counter_enexo_34 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_35 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_17_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_35 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_35 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_17_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_35 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_1_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_905_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_17_enex5
        ) begin
      reg_act_regs_data_1_1_2_enexo_2 <= act_regs_data_and_905_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_1_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_873_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_17_enex5
        ) begin
      reg_act_regs_data_3_1_2_enexo_2 <= act_regs_data_and_873_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_1_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_921_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_17_enex5
        ) begin
      reg_act_regs_data_0_1_2_enexo_2 <= act_regs_data_and_921_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_1_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_889_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_17_enex5
        ) begin
      reg_act_regs_data_2_1_2_enexo_2 <= act_regs_data_and_889_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_35 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_17_enex5
        ) begin
      reg_act_config_inst_counter_enexo_35 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_36 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_18_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_36 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_36 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_18_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_36 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_4_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_886_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_18_enex5
        ) begin
      reg_act_regs_data_2_4_2_enexo_2 <= act_regs_data_and_886_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_4_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_870_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_18_enex5
        ) begin
      reg_act_regs_data_3_4_2_enexo_2 <= act_regs_data_and_870_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_4_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_902_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_18_enex5
        ) begin
      reg_act_regs_data_1_4_2_enexo_2 <= act_regs_data_and_902_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_4_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_918_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_18_enex5
        ) begin
      reg_act_regs_data_0_4_2_enexo_2 <= act_regs_data_and_918_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_36 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_18_enex5
        ) begin
      reg_act_config_inst_counter_enexo_36 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_37 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_19_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_37 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_37 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_19_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_37 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_5_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_917_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_19_enex5
        ) begin
      reg_act_regs_data_0_5_2_enexo_2 <= act_regs_data_and_917_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_5_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_885_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_19_enex5
        ) begin
      reg_act_regs_data_2_5_2_enexo_2 <= act_regs_data_and_885_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_5_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_869_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_19_enex5
        ) begin
      reg_act_regs_data_3_5_2_enexo_2 <= act_regs_data_and_869_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_5_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_901_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_19_enex5
        ) begin
      reg_act_regs_data_1_5_2_enexo_2 <= act_regs_data_and_901_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_37 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_19_enex5
        ) begin
      reg_act_config_inst_counter_enexo_37 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_38 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_20_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_38 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_38 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_20_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_38 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_6_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_868_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_20_enex5
        ) begin
      reg_act_regs_data_3_6_2_enexo_2 <= act_regs_data_and_868_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_6_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_900_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_20_enex5
        ) begin
      reg_act_regs_data_1_6_2_enexo_2 <= act_regs_data_and_900_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_6_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_916_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_20_enex5
        ) begin
      reg_act_regs_data_0_6_2_enexo_2 <= act_regs_data_and_916_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_6_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_884_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_20_enex5
        ) begin
      reg_act_regs_data_2_6_2_enexo_2 <= act_regs_data_and_884_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_38 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_20_enex5
        ) begin
      reg_act_config_inst_counter_enexo_38 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_39 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_21_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_39 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_39 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_21_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_39 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_7_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_883_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_21_enex5
        ) begin
      reg_act_regs_data_2_7_2_enexo_2 <= act_regs_data_and_883_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_7_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_899_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_21_enex5
        ) begin
      reg_act_regs_data_1_7_2_enexo_2 <= act_regs_data_and_899_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_7_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_915_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_21_enex5
        ) begin
      reg_act_regs_data_0_7_2_enexo_2 <= act_regs_data_and_915_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_7_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_867_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_21_enex5
        ) begin
      reg_act_regs_data_3_7_2_enexo_2 <= act_regs_data_and_867_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_39 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_21_enex5
        ) begin
      reg_act_config_inst_counter_enexo_39 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_40 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_22_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_40 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_40 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_22_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_40 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_8_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_866_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_22_enex5
        ) begin
      reg_act_regs_data_3_8_2_enexo_2 <= act_regs_data_and_866_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_8_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_898_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_22_enex5
        ) begin
      reg_act_regs_data_1_8_2_enexo_2 <= act_regs_data_and_898_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_8_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_914_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_22_enex5
        ) begin
      reg_act_regs_data_0_8_2_enexo_2 <= act_regs_data_and_914_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_8_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_882_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_22_enex5
        ) begin
      reg_act_regs_data_2_8_2_enexo_2 <= act_regs_data_and_882_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_40 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_22_enex5
        ) begin
      reg_act_config_inst_counter_enexo_40 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_41 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_23_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_41 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_41 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_23_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_41 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_9_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_897_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_23_enex5
        ) begin
      reg_act_regs_data_1_9_2_enexo_2 <= act_regs_data_and_897_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_9_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_913_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_23_enex5
        ) begin
      reg_act_regs_data_0_9_2_enexo_2 <= act_regs_data_and_913_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_9_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_881_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_23_enex5
        ) begin
      reg_act_regs_data_2_9_2_enexo_2 <= act_regs_data_and_881_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_9_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_865_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_23_enex5
        ) begin
      reg_act_regs_data_3_9_2_enexo_2 <= act_regs_data_and_865_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_41 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_23_enex5
        ) begin
      reg_act_config_inst_counter_enexo_41 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_42 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_24_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_42 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_42 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_24_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_42 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_10_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_912_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_24_enex5
        ) begin
      reg_act_regs_data_0_10_2_enexo_2 <= act_regs_data_and_912_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_10_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_896_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_24_enex5
        ) begin
      reg_act_regs_data_1_10_2_enexo_2 <= act_regs_data_and_896_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_10_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_880_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_24_enex5
        ) begin
      reg_act_regs_data_2_10_2_enexo_2 <= act_regs_data_and_880_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_10_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_864_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_24_enex5
        ) begin
      reg_act_regs_data_3_10_2_enexo_2 <= act_regs_data_and_864_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_42 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_24_enex5
        ) begin
      reg_act_config_inst_counter_enexo_42 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_43 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_25_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_43 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_43 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_25_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_43 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_11_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_879_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_25_enex5
        ) begin
      reg_act_regs_data_2_11_2_enexo_2 <= act_regs_data_and_879_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_11_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_863_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_25_enex5
        ) begin
      reg_act_regs_data_3_11_2_enexo_2 <= act_regs_data_and_863_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_11_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_895_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_25_enex5
        ) begin
      reg_act_regs_data_1_11_2_enexo_2 <= act_regs_data_and_895_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_11_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_911_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_25_enex5
        ) begin
      reg_act_regs_data_0_11_2_enexo_2 <= act_regs_data_and_911_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_43 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_25_enex5
        ) begin
      reg_act_config_inst_counter_enexo_43 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_44 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_26_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_44 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_44 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_26_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_44 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_12_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_894_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_26_enex5
        ) begin
      reg_act_regs_data_1_12_2_enexo_2 <= act_regs_data_and_894_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_12_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_878_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_26_enex5
        ) begin
      reg_act_regs_data_2_12_2_enexo_2 <= act_regs_data_and_878_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_12_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_910_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_26_enex5
        ) begin
      reg_act_regs_data_0_12_2_enexo_2 <= act_regs_data_and_910_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_12_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_862_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_26_enex5
        ) begin
      reg_act_regs_data_3_12_2_enexo_2 <= act_regs_data_and_862_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_44 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_26_enex5
        ) begin
      reg_act_config_inst_counter_enexo_44 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_45 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_27_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_45 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_45 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_27_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_45 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_13_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_893_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_27_enex5
        ) begin
      reg_act_regs_data_1_13_2_enexo_2 <= act_regs_data_and_893_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_13_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_909_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_27_enex5
        ) begin
      reg_act_regs_data_0_13_2_enexo_2 <= act_regs_data_and_909_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_13_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_861_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_27_enex5
        ) begin
      reg_act_regs_data_3_13_2_enexo_2 <= act_regs_data_and_861_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_13_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_877_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_27_enex5
        ) begin
      reg_act_regs_data_2_13_2_enexo_2 <= act_regs_data_and_877_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_45 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_27_enex5
        ) begin
      reg_act_config_inst_counter_enexo_45 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_46 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_28_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_46 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_46 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_28_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_46 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_14_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_860_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_28_enex5
        ) begin
      reg_act_regs_data_3_14_2_enexo_2 <= act_regs_data_and_860_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_14_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_908_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_28_enex5
        ) begin
      reg_act_regs_data_0_14_2_enexo_2 <= act_regs_data_and_908_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_14_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_892_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_28_enex5
        ) begin
      reg_act_regs_data_1_14_2_enexo_2 <= act_regs_data_and_892_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_14_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_876_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_28_enex5
        ) begin
      reg_act_regs_data_2_14_2_enexo_2 <= act_regs_data_and_876_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_46 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_28_enex5
        ) begin
      reg_act_config_inst_counter_enexo_46 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_47 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_29_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_47 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_47 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_29_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_47 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_15_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_891_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_29_enex5
        ) begin
      reg_act_regs_data_1_15_2_enexo_2 <= act_regs_data_and_891_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_15_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_875_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_29_enex5
        ) begin
      reg_act_regs_data_2_15_2_enexo_2 <= act_regs_data_and_875_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_15_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_907_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_29_enex5
        ) begin
      reg_act_regs_data_0_15_2_enexo_2 <= act_regs_data_and_907_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_47 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_29_enex5
        ) begin
      reg_act_config_inst_counter_enexo_47 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_15_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_859_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_29_enex5
        ) begin
      reg_act_regs_data_3_15_2_enexo_2 <= act_regs_data_and_859_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_48 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_48 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_48 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_48 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_2_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_920_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_enex5
        ) begin
      reg_act_regs_data_0_2_2_enexo_3 <= act_regs_data_and_920_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_2_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_888_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_enex5
        ) begin
      reg_act_regs_data_2_2_2_enexo_3 <= act_regs_data_and_888_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_2_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_904_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_enex5
        ) begin
      reg_act_regs_data_1_2_2_enexo_3 <= act_regs_data_and_904_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_2_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_872_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_enex5
        ) begin
      reg_act_regs_data_3_2_2_enexo_3 <= act_regs_data_and_872_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_48 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_enex5
        ) begin
      reg_act_config_inst_counter_enexo_48 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_49 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_15_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_49 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_49 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_15_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_49 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_11_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_879_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_15_enex5
        ) begin
      reg_act_regs_data_2_11_2_enexo_3 <= act_regs_data_and_879_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_11_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_863_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_15_enex5
        ) begin
      reg_act_regs_data_3_11_2_enexo_3 <= act_regs_data_and_863_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_11_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_895_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_15_enex5
        ) begin
      reg_act_regs_data_1_11_2_enexo_3 <= act_regs_data_and_895_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_11_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_911_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_15_enex5
        ) begin
      reg_act_regs_data_0_11_2_enexo_3 <= act_regs_data_and_911_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_49 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_15_enex5
        ) begin
      reg_act_config_inst_counter_enexo_49 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_50 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | ActUnit_RunInst_switch_lp_and_816_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_50 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_50 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | ActUnit_RunInst_switch_lp_and_816_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_50 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_0_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_890_enex5 | ActUnit_RunInst_switch_lp_and_816_enex5
        ) begin
      reg_act_regs_data_2_0_2_enexo_3 <= act_regs_data_and_890_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_0_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_874_enex5 | ActUnit_RunInst_switch_lp_and_816_enex5
        ) begin
      reg_act_regs_data_3_0_2_enexo_3 <= act_regs_data_and_874_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_0_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_906_enex5 | ActUnit_RunInst_switch_lp_and_816_enex5
        ) begin
      reg_act_regs_data_1_0_2_enexo_3 <= act_regs_data_and_906_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_0_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_922_enex5 | ActUnit_RunInst_switch_lp_and_816_enex5
        ) begin
      reg_act_regs_data_0_0_2_enexo_3 <= act_regs_data_and_922_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_50 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | ActUnit_RunInst_switch_lp_and_816_enex5
        ) begin
      reg_act_config_inst_counter_enexo_50 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_51 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_16_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_51 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_51 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_16_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_51 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_1_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_905_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_16_enex5
        ) begin
      reg_act_regs_data_1_1_2_enexo_3 <= act_regs_data_and_905_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_1_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_873_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_16_enex5
        ) begin
      reg_act_regs_data_3_1_2_enexo_3 <= act_regs_data_and_873_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_1_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_921_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_16_enex5
        ) begin
      reg_act_regs_data_0_1_2_enexo_3 <= act_regs_data_and_921_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_1_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_889_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_16_enex5
        ) begin
      reg_act_regs_data_2_1_2_enexo_3 <= act_regs_data_and_889_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_51 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_16_enex5
        ) begin
      reg_act_config_inst_counter_enexo_51 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_52 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_17_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_52 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_52 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_17_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_52 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_3_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_887_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_17_enex5
        ) begin
      reg_act_regs_data_2_3_2_enexo_3 <= act_regs_data_and_887_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_3_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_871_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_17_enex5
        ) begin
      reg_act_regs_data_3_3_2_enexo_3 <= act_regs_data_and_871_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_3_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_903_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_17_enex5
        ) begin
      reg_act_regs_data_1_3_2_enexo_3 <= act_regs_data_and_903_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_3_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_919_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_17_enex5
        ) begin
      reg_act_regs_data_0_3_2_enexo_3 <= act_regs_data_and_919_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_52 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_17_enex5
        ) begin
      reg_act_config_inst_counter_enexo_52 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_53 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_18_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_53 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_53 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_18_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_53 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_4_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_886_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_18_enex5
        ) begin
      reg_act_regs_data_2_4_2_enexo_3 <= act_regs_data_and_886_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_4_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_870_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_18_enex5
        ) begin
      reg_act_regs_data_3_4_2_enexo_3 <= act_regs_data_and_870_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_4_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_902_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_18_enex5
        ) begin
      reg_act_regs_data_1_4_2_enexo_3 <= act_regs_data_and_902_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_4_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_918_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_18_enex5
        ) begin
      reg_act_regs_data_0_4_2_enexo_3 <= act_regs_data_and_918_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_53 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_18_enex5
        ) begin
      reg_act_config_inst_counter_enexo_53 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_54 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_19_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_54 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_54 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_19_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_54 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_5_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_917_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_19_enex5
        ) begin
      reg_act_regs_data_0_5_2_enexo_3 <= act_regs_data_and_917_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_5_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_885_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_19_enex5
        ) begin
      reg_act_regs_data_2_5_2_enexo_3 <= act_regs_data_and_885_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_5_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_869_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_19_enex5
        ) begin
      reg_act_regs_data_3_5_2_enexo_3 <= act_regs_data_and_869_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_5_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_901_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_19_enex5
        ) begin
      reg_act_regs_data_1_5_2_enexo_3 <= act_regs_data_and_901_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_54 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_19_enex5
        ) begin
      reg_act_config_inst_counter_enexo_54 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_55 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_20_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_55 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_55 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_20_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_55 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_6_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_868_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_20_enex5
        ) begin
      reg_act_regs_data_3_6_2_enexo_3 <= act_regs_data_and_868_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_6_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_900_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_20_enex5
        ) begin
      reg_act_regs_data_1_6_2_enexo_3 <= act_regs_data_and_900_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_6_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_916_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_20_enex5
        ) begin
      reg_act_regs_data_0_6_2_enexo_3 <= act_regs_data_and_916_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_6_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_884_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_20_enex5
        ) begin
      reg_act_regs_data_2_6_2_enexo_3 <= act_regs_data_and_884_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_55 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_20_enex5
        ) begin
      reg_act_config_inst_counter_enexo_55 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_56 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_21_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_56 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_56 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_21_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_56 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_7_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_883_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_21_enex5
        ) begin
      reg_act_regs_data_2_7_2_enexo_3 <= act_regs_data_and_883_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_7_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_899_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_21_enex5
        ) begin
      reg_act_regs_data_1_7_2_enexo_3 <= act_regs_data_and_899_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_7_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_915_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_21_enex5
        ) begin
      reg_act_regs_data_0_7_2_enexo_3 <= act_regs_data_and_915_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_7_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_867_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_21_enex5
        ) begin
      reg_act_regs_data_3_7_2_enexo_3 <= act_regs_data_and_867_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_56 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_21_enex5
        ) begin
      reg_act_config_inst_counter_enexo_56 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_57 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_22_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_57 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_57 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_22_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_57 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_8_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_866_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_22_enex5
        ) begin
      reg_act_regs_data_3_8_2_enexo_3 <= act_regs_data_and_866_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_8_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_898_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_22_enex5
        ) begin
      reg_act_regs_data_1_8_2_enexo_3 <= act_regs_data_and_898_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_8_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_914_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_22_enex5
        ) begin
      reg_act_regs_data_0_8_2_enexo_3 <= act_regs_data_and_914_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_8_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_882_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_22_enex5
        ) begin
      reg_act_regs_data_2_8_2_enexo_3 <= act_regs_data_and_882_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_57 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_22_enex5
        ) begin
      reg_act_config_inst_counter_enexo_57 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_58 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_23_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_58 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_58 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_23_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_58 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_9_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_897_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_23_enex5
        ) begin
      reg_act_regs_data_1_9_2_enexo_3 <= act_regs_data_and_897_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_9_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_913_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_23_enex5
        ) begin
      reg_act_regs_data_0_9_2_enexo_3 <= act_regs_data_and_913_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_9_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_881_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_23_enex5
        ) begin
      reg_act_regs_data_2_9_2_enexo_3 <= act_regs_data_and_881_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_9_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_865_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_23_enex5
        ) begin
      reg_act_regs_data_3_9_2_enexo_3 <= act_regs_data_and_865_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_58 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_23_enex5
        ) begin
      reg_act_config_inst_counter_enexo_58 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_59 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_24_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_59 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_59 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_24_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_59 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_10_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_912_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_24_enex5
        ) begin
      reg_act_regs_data_0_10_2_enexo_3 <= act_regs_data_and_912_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_10_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_896_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_24_enex5
        ) begin
      reg_act_regs_data_1_10_2_enexo_3 <= act_regs_data_and_896_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_10_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_880_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_24_enex5
        ) begin
      reg_act_regs_data_2_10_2_enexo_3 <= act_regs_data_and_880_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_10_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_864_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_24_enex5
        ) begin
      reg_act_regs_data_3_10_2_enexo_3 <= act_regs_data_and_864_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_59 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_24_enex5
        ) begin
      reg_act_config_inst_counter_enexo_59 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_60 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_25_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_60 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_60 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_25_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_60 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_12_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_894_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_25_enex5
        ) begin
      reg_act_regs_data_1_12_2_enexo_3 <= act_regs_data_and_894_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_12_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_878_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_25_enex5
        ) begin
      reg_act_regs_data_2_12_2_enexo_3 <= act_regs_data_and_878_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_12_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_910_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_25_enex5
        ) begin
      reg_act_regs_data_0_12_2_enexo_3 <= act_regs_data_and_910_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_12_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_862_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_25_enex5
        ) begin
      reg_act_regs_data_3_12_2_enexo_3 <= act_regs_data_and_862_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_60 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_25_enex5
        ) begin
      reg_act_config_inst_counter_enexo_60 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_61 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_26_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_61 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_61 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_26_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_61 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_13_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_893_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_26_enex5
        ) begin
      reg_act_regs_data_1_13_2_enexo_3 <= act_regs_data_and_893_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_13_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_909_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_26_enex5
        ) begin
      reg_act_regs_data_0_13_2_enexo_3 <= act_regs_data_and_909_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_13_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_861_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_26_enex5
        ) begin
      reg_act_regs_data_3_13_2_enexo_3 <= act_regs_data_and_861_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_13_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_877_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_26_enex5
        ) begin
      reg_act_regs_data_2_13_2_enexo_3 <= act_regs_data_and_877_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_61 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_26_enex5
        ) begin
      reg_act_config_inst_counter_enexo_61 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_62 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_27_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_62 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_62 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_27_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_62 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_14_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_860_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_27_enex5
        ) begin
      reg_act_regs_data_3_14_2_enexo_3 <= act_regs_data_and_860_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_14_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_908_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_27_enex5
        ) begin
      reg_act_regs_data_0_14_2_enexo_3 <= act_regs_data_and_908_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_14_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_892_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_27_enex5
        ) begin
      reg_act_regs_data_1_14_2_enexo_3 <= act_regs_data_and_892_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_14_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_876_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_27_enex5
        ) begin
      reg_act_regs_data_2_14_2_enexo_3 <= act_regs_data_and_876_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_62 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_27_enex5
        ) begin
      reg_act_config_inst_counter_enexo_62 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_63 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_28_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_63 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_63 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_28_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_63 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_15_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_891_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_28_enex5
        ) begin
      reg_act_regs_data_1_15_2_enexo_3 <= act_regs_data_and_891_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_15_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_875_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_28_enex5
        ) begin
      reg_act_regs_data_2_15_2_enexo_3 <= act_regs_data_and_875_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_15_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_907_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_28_enex5
        ) begin
      reg_act_regs_data_0_15_2_enexo_3 <= act_regs_data_and_907_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_63 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_28_enex5
        ) begin
      reg_act_config_inst_counter_enexo_63 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_15_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_859_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_28_enex5
        ) begin
      reg_act_regs_data_3_15_2_enexo_3 <= act_regs_data_and_859_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_64 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | ActUnit_RunInst_curr_inst_and_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_64 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_64 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | ActUnit_RunInst_curr_inst_and_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_64 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_64 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | ActUnit_RunInst_curr_inst_and_enex5
        ) begin
      reg_act_config_inst_counter_enexo_64 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_65 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | ActUnit_RunInst_switch_lp_and_817_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_65 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_65 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | ActUnit_RunInst_switch_lp_and_817_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_65 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_0_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_890_enex5 | ActUnit_RunInst_switch_lp_and_817_enex5
        ) begin
      reg_act_regs_data_2_0_2_enexo_4 <= act_regs_data_and_890_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_0_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_874_enex5 | ActUnit_RunInst_switch_lp_and_817_enex5
        ) begin
      reg_act_regs_data_3_0_2_enexo_4 <= act_regs_data_and_874_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_0_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_906_enex5 | ActUnit_RunInst_switch_lp_and_817_enex5
        ) begin
      reg_act_regs_data_1_0_2_enexo_4 <= act_regs_data_and_906_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_0_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_922_enex5 | ActUnit_RunInst_switch_lp_and_817_enex5
        ) begin
      reg_act_regs_data_0_0_2_enexo_4 <= act_regs_data_and_922_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_65 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | ActUnit_RunInst_switch_lp_and_817_enex5
        ) begin
      reg_act_config_inst_counter_enexo_65 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_66 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_3_for_and_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_66 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_66 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_3_for_and_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_66 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_1_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_905_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_enex5
        ) begin
      reg_act_regs_data_1_1_2_enexo_4 <= act_regs_data_and_905_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_1_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_873_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_enex5
        ) begin
      reg_act_regs_data_3_1_2_enexo_4 <= act_regs_data_and_873_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_1_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_921_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_enex5
        ) begin
      reg_act_regs_data_0_1_2_enexo_4 <= act_regs_data_and_921_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_1_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_889_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_enex5
        ) begin
      reg_act_regs_data_2_1_2_enexo_4 <= act_regs_data_and_889_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_66 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_3_for_and_enex5
        ) begin
      reg_act_config_inst_counter_enexo_66 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_67 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_3_for_and_15_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_67 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_67 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_3_for_and_15_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_67 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_2_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_920_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_15_enex5
        ) begin
      reg_act_regs_data_0_2_2_enexo_4 <= act_regs_data_and_920_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_2_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_888_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_15_enex5
        ) begin
      reg_act_regs_data_2_2_2_enexo_4 <= act_regs_data_and_888_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_2_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_904_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_15_enex5
        ) begin
      reg_act_regs_data_1_2_2_enexo_4 <= act_regs_data_and_904_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_2_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_872_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_15_enex5
        ) begin
      reg_act_regs_data_3_2_2_enexo_4 <= act_regs_data_and_872_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_67 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_3_for_and_15_enex5
        ) begin
      reg_act_config_inst_counter_enexo_67 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_68 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_3_for_and_16_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_68 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_68 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_3_for_and_16_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_68 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_3_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_887_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_16_enex5
        ) begin
      reg_act_regs_data_2_3_2_enexo_4 <= act_regs_data_and_887_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_3_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_871_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_16_enex5
        ) begin
      reg_act_regs_data_3_3_2_enexo_4 <= act_regs_data_and_871_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_3_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_903_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_16_enex5
        ) begin
      reg_act_regs_data_1_3_2_enexo_4 <= act_regs_data_and_903_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_3_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_919_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_16_enex5
        ) begin
      reg_act_regs_data_0_3_2_enexo_4 <= act_regs_data_and_919_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_68 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_3_for_and_16_enex5
        ) begin
      reg_act_config_inst_counter_enexo_68 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_69 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_3_for_and_17_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_69 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_69 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_3_for_and_17_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_69 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_4_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_886_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_17_enex5
        ) begin
      reg_act_regs_data_2_4_2_enexo_4 <= act_regs_data_and_886_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_4_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_870_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_17_enex5
        ) begin
      reg_act_regs_data_3_4_2_enexo_4 <= act_regs_data_and_870_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_4_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_902_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_17_enex5
        ) begin
      reg_act_regs_data_1_4_2_enexo_4 <= act_regs_data_and_902_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_4_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_918_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_17_enex5
        ) begin
      reg_act_regs_data_0_4_2_enexo_4 <= act_regs_data_and_918_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_69 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_3_for_and_17_enex5
        ) begin
      reg_act_config_inst_counter_enexo_69 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_70 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_3_for_and_18_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_70 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_70 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_3_for_and_18_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_70 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_5_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_917_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_18_enex5
        ) begin
      reg_act_regs_data_0_5_2_enexo_4 <= act_regs_data_and_917_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_5_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_885_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_18_enex5
        ) begin
      reg_act_regs_data_2_5_2_enexo_4 <= act_regs_data_and_885_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_5_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_869_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_18_enex5
        ) begin
      reg_act_regs_data_3_5_2_enexo_4 <= act_regs_data_and_869_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_5_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_901_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_18_enex5
        ) begin
      reg_act_regs_data_1_5_2_enexo_4 <= act_regs_data_and_901_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_70 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_3_for_and_18_enex5
        ) begin
      reg_act_config_inst_counter_enexo_70 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_71 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_3_for_and_19_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_71 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_71 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_3_for_and_19_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_71 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_6_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_868_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_19_enex5
        ) begin
      reg_act_regs_data_3_6_2_enexo_4 <= act_regs_data_and_868_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_6_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_900_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_19_enex5
        ) begin
      reg_act_regs_data_1_6_2_enexo_4 <= act_regs_data_and_900_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_6_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_916_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_19_enex5
        ) begin
      reg_act_regs_data_0_6_2_enexo_4 <= act_regs_data_and_916_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_6_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_884_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_19_enex5
        ) begin
      reg_act_regs_data_2_6_2_enexo_4 <= act_regs_data_and_884_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_71 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_3_for_and_19_enex5
        ) begin
      reg_act_config_inst_counter_enexo_71 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_72 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_3_for_and_20_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_72 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_72 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_3_for_and_20_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_72 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_7_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_883_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_20_enex5
        ) begin
      reg_act_regs_data_2_7_2_enexo_4 <= act_regs_data_and_883_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_7_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_899_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_20_enex5
        ) begin
      reg_act_regs_data_1_7_2_enexo_4 <= act_regs_data_and_899_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_7_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_915_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_20_enex5
        ) begin
      reg_act_regs_data_0_7_2_enexo_4 <= act_regs_data_and_915_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_7_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_867_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_20_enex5
        ) begin
      reg_act_regs_data_3_7_2_enexo_4 <= act_regs_data_and_867_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_72 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_3_for_and_20_enex5
        ) begin
      reg_act_config_inst_counter_enexo_72 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_73 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_3_for_and_21_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_73 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_73 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_3_for_and_21_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_73 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_8_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_866_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_21_enex5
        ) begin
      reg_act_regs_data_3_8_2_enexo_4 <= act_regs_data_and_866_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_8_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_898_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_21_enex5
        ) begin
      reg_act_regs_data_1_8_2_enexo_4 <= act_regs_data_and_898_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_8_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_914_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_21_enex5
        ) begin
      reg_act_regs_data_0_8_2_enexo_4 <= act_regs_data_and_914_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_8_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_882_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_21_enex5
        ) begin
      reg_act_regs_data_2_8_2_enexo_4 <= act_regs_data_and_882_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_73 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_3_for_and_21_enex5
        ) begin
      reg_act_config_inst_counter_enexo_73 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_74 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_3_for_and_22_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_74 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_74 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_3_for_and_22_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_74 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_11_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_879_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_22_enex5
        ) begin
      reg_act_regs_data_2_11_2_enexo_4 <= act_regs_data_and_879_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_11_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_863_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_22_enex5
        ) begin
      reg_act_regs_data_3_11_2_enexo_4 <= act_regs_data_and_863_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_11_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_895_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_22_enex5
        ) begin
      reg_act_regs_data_1_11_2_enexo_4 <= act_regs_data_and_895_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_11_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_911_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_22_enex5
        ) begin
      reg_act_regs_data_0_11_2_enexo_4 <= act_regs_data_and_911_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_74 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_3_for_and_22_enex5
        ) begin
      reg_act_config_inst_counter_enexo_74 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_75 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_3_for_and_23_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_75 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_75 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_3_for_and_23_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_75 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_12_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_894_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_23_enex5
        ) begin
      reg_act_regs_data_1_12_2_enexo_4 <= act_regs_data_and_894_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_12_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_878_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_23_enex5
        ) begin
      reg_act_regs_data_2_12_2_enexo_4 <= act_regs_data_and_878_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_12_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_910_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_23_enex5
        ) begin
      reg_act_regs_data_0_12_2_enexo_4 <= act_regs_data_and_910_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_12_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_862_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_23_enex5
        ) begin
      reg_act_regs_data_3_12_2_enexo_4 <= act_regs_data_and_862_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_75 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_3_for_and_23_enex5
        ) begin
      reg_act_config_inst_counter_enexo_75 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_76 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_3_for_and_24_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_76 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_76 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_3_for_and_24_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_76 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_13_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_893_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_24_enex5
        ) begin
      reg_act_regs_data_1_13_2_enexo_4 <= act_regs_data_and_893_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_13_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_909_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_24_enex5
        ) begin
      reg_act_regs_data_0_13_2_enexo_4 <= act_regs_data_and_909_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_13_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_861_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_24_enex5
        ) begin
      reg_act_regs_data_3_13_2_enexo_4 <= act_regs_data_and_861_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_13_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_877_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_24_enex5
        ) begin
      reg_act_regs_data_2_13_2_enexo_4 <= act_regs_data_and_877_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_76 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_3_for_and_24_enex5
        ) begin
      reg_act_config_inst_counter_enexo_76 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_77 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_3_for_and_25_enex5
        ) begin
      reg_act_config_inst_regs_1_sva_dfm_5_enexo_77 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_77 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_3_for_and_25_enex5
        ) begin
      reg_act_config_inst_regs_17_sva_dfm_6_enexo_77 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_14_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_860_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_25_enex5
        ) begin
      reg_act_regs_data_3_14_2_enexo_4 <= act_regs_data_and_860_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_14_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_908_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_25_enex5
        ) begin
      reg_act_regs_data_0_14_2_enexo_4 <= act_regs_data_and_908_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_14_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_892_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_25_enex5
        ) begin
      reg_act_regs_data_1_14_2_enexo_4 <= act_regs_data_and_892_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_14_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_876_enex5 | nv_scvector_cctor_nv_scvector_3_for_and_25_enex5
        ) begin
      reg_act_regs_data_2_14_2_enexo_4 <= act_regs_data_and_876_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_77 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_3_for_and_25_enex5
        ) begin
      reg_act_config_inst_counter_enexo_77 <= act_config_inst_counter_and_tmp;
    end
  end
  assign and_843_nl = and_dcpl_553 & and_dcpl_789 & while_asn_262_itm;
  assign while_else_1_while_else_1_nand_1_nl = ~(act_config_InstIncr_if_act_config_InstIncr_if_if_nor_tmp
      & act_config_InstIncr_act_config_InstIncr_if_and_svs_1 & is_incr_lpi_1_dfm_1);
  assign nl_operator_8_false_acc_nl = act_config_output_counter_sva_dfm_3 + 8'b00000001;
  assign operator_8_false_acc_nl = nl_operator_8_false_acc_nl[7:0];
  assign act_config_InstIncr_if_not_nl = ~ act_config_InstIncr_if_act_config_InstIncr_if_if_nor_mdf_sva;
  assign act_config_InstIncr_if_act_config_InstIncr_if_and_1_nl = MUX_v_8_2_2(8'b00000000,
      operator_8_false_acc_nl, act_config_InstIncr_if_not_nl);
  assign nl_operator_5_false_acc_nl = act_config_inst_counter_sva_dfm_3 + 5'b00001;
  assign operator_5_false_acc_nl = nl_operator_5_false_acc_nl[4:0];
  assign act_config_InstIncr_if_not_7_nl = ~ act_config_InstIncr_act_config_InstIncr_if_and_svs_1;
  assign act_config_InstIncr_act_config_InstIncr_and_1_nl = MUX_v_5_2_2(5'b00000,
      operator_5_false_acc_nl, act_config_InstIncr_if_not_7_nl);
  assign and_880_nl = nor_61_cse & and_dcpl_829;
  assign nor_678_nl = ~((act_config_inst_regs_0_sva_dfm_5[7:4]!=4'b0010));
  assign nor_679_nl = ~((act_config_inst_regs_1_sva_dfm_5[7:4]!=4'b0010));
  assign mux_291_nl = MUX_s_1_2_2(nor_678_nl, nor_679_nl, act_config_inst_counter_sva[0]);
  assign nor_680_nl = ~((act_config_inst_regs_2_sva_dfm_5[7:4]!=4'b0010));
  assign nor_681_nl = ~((act_config_inst_regs_3_sva_dfm_5[7:4]!=4'b0010));
  assign mux_290_nl = MUX_s_1_2_2(nor_680_nl, nor_681_nl, act_config_inst_counter_sva[0]);
  assign mux_292_nl = MUX_s_1_2_2(mux_291_nl, mux_290_nl, act_config_inst_counter_sva[1]);
  assign nor_682_nl = ~((act_config_inst_regs_4_sva_dfm_5[7:4]!=4'b0010));
  assign nor_683_nl = ~((act_config_inst_regs_5_sva_dfm_5[7:4]!=4'b0010));
  assign mux_288_nl = MUX_s_1_2_2(nor_682_nl, nor_683_nl, act_config_inst_counter_sva[0]);
  assign nor_684_nl = ~((act_config_inst_regs_6_sva_dfm_5[7:4]!=4'b0010));
  assign nor_685_nl = ~((act_config_inst_regs_7_sva_dfm_5[7:4]!=4'b0010));
  assign mux_287_nl = MUX_s_1_2_2(nor_684_nl, nor_685_nl, act_config_inst_counter_sva[0]);
  assign mux_289_nl = MUX_s_1_2_2(mux_288_nl, mux_287_nl, act_config_inst_counter_sva[1]);
  assign mux_293_nl = MUX_s_1_2_2(mux_292_nl, mux_289_nl, act_config_inst_counter_sva[2]);
  assign nor_686_nl = ~((act_config_inst_regs_8_sva_dfm_5[7:4]!=4'b0010));
  assign nor_687_nl = ~((act_config_inst_regs_9_sva_dfm_5[7:4]!=4'b0010));
  assign mux_284_nl = MUX_s_1_2_2(nor_686_nl, nor_687_nl, act_config_inst_counter_sva[0]);
  assign nor_688_nl = ~((act_config_inst_regs_10_sva_dfm_5[7:4]!=4'b0010));
  assign nor_689_nl = ~((act_config_inst_regs_11_sva_dfm_5[7:4]!=4'b0010));
  assign mux_283_nl = MUX_s_1_2_2(nor_688_nl, nor_689_nl, act_config_inst_counter_sva[0]);
  assign mux_285_nl = MUX_s_1_2_2(mux_284_nl, mux_283_nl, act_config_inst_counter_sva[1]);
  assign nor_690_nl = ~((act_config_inst_regs_12_sva_dfm_5[7:4]!=4'b0010));
  assign nor_691_nl = ~((act_config_inst_regs_13_sva_dfm_5[7:4]!=4'b0010));
  assign mux_281_nl = MUX_s_1_2_2(nor_690_nl, nor_691_nl, act_config_inst_counter_sva[0]);
  assign nor_692_nl = ~((act_config_inst_regs_14_sva_dfm_5[7:4]!=4'b0010));
  assign nor_693_nl = ~((act_config_inst_regs_15_sva_dfm_5[7:4]!=4'b0010));
  assign mux_280_nl = MUX_s_1_2_2(nor_692_nl, nor_693_nl, act_config_inst_counter_sva[0]);
  assign mux_282_nl = MUX_s_1_2_2(mux_281_nl, mux_280_nl, act_config_inst_counter_sva[1]);
  assign mux_286_nl = MUX_s_1_2_2(mux_285_nl, mux_282_nl, act_config_inst_counter_sva[2]);
  assign mux_294_nl = MUX_s_1_2_2(mux_293_nl, mux_286_nl, act_config_inst_counter_sva[3]);
  assign nor_694_nl = ~((act_config_inst_regs_16_sva_dfm_6[7:4]!=4'b0010));
  assign nor_695_nl = ~((act_config_inst_regs_17_sva_dfm_6[7:4]!=4'b0010));
  assign mux_276_nl = MUX_s_1_2_2(nor_694_nl, nor_695_nl, act_config_inst_counter_sva[0]);
  assign nor_696_nl = ~((act_config_inst_regs_18_sva_dfm_6[7:4]!=4'b0010));
  assign nor_697_nl = ~((act_config_inst_regs_19_sva_dfm_6[7:4]!=4'b0010));
  assign mux_275_nl = MUX_s_1_2_2(nor_696_nl, nor_697_nl, act_config_inst_counter_sva[0]);
  assign mux_277_nl = MUX_s_1_2_2(mux_276_nl, mux_275_nl, act_config_inst_counter_sva[1]);
  assign nor_698_nl = ~((act_config_inst_regs_20_sva_dfm_6[7:4]!=4'b0010));
  assign nor_699_nl = ~((act_config_inst_regs_21_sva_dfm_6[7:4]!=4'b0010));
  assign mux_273_nl = MUX_s_1_2_2(nor_698_nl, nor_699_nl, act_config_inst_counter_sva[0]);
  assign nor_700_nl = ~((act_config_inst_regs_22_sva_dfm_6[7:4]!=4'b0010));
  assign nor_701_nl = ~((act_config_inst_regs_23_sva_dfm_6[7:4]!=4'b0010));
  assign mux_272_nl = MUX_s_1_2_2(nor_700_nl, nor_701_nl, act_config_inst_counter_sva[0]);
  assign mux_274_nl = MUX_s_1_2_2(mux_273_nl, mux_272_nl, act_config_inst_counter_sva[1]);
  assign mux_278_nl = MUX_s_1_2_2(mux_277_nl, mux_274_nl, act_config_inst_counter_sva[2]);
  assign nor_702_nl = ~((act_config_inst_regs_24_sva_dfm_6[7:4]!=4'b0010));
  assign nor_703_nl = ~((act_config_inst_regs_25_sva_dfm_6[7:4]!=4'b0010));
  assign mux_269_nl = MUX_s_1_2_2(nor_702_nl, nor_703_nl, act_config_inst_counter_sva[0]);
  assign nor_704_nl = ~((act_config_inst_regs_26_sva_dfm_6[7:4]!=4'b0010));
  assign nor_705_nl = ~((act_config_inst_regs_27_sva_dfm_6[7:4]!=4'b0010));
  assign mux_268_nl = MUX_s_1_2_2(nor_704_nl, nor_705_nl, act_config_inst_counter_sva[0]);
  assign mux_270_nl = MUX_s_1_2_2(mux_269_nl, mux_268_nl, act_config_inst_counter_sva[1]);
  assign nor_706_nl = ~((act_config_inst_regs_28_sva_dfm_6[7:4]!=4'b0010));
  assign nor_707_nl = ~((act_config_inst_regs_29_sva_dfm_6[7:4]!=4'b0010));
  assign mux_266_nl = MUX_s_1_2_2(nor_706_nl, nor_707_nl, act_config_inst_counter_sva[0]);
  assign nor_708_nl = ~((act_config_inst_regs_30_sva_dfm_6[7:4]!=4'b0010));
  assign nor_709_nl = ~((act_config_inst_regs_31_sva_dfm_6[7:4]!=4'b0010));
  assign mux_nl = MUX_s_1_2_2(nor_708_nl, nor_709_nl, act_config_inst_counter_sva[0]);
  assign mux_267_nl = MUX_s_1_2_2(mux_266_nl, mux_nl, act_config_inst_counter_sva[1]);
  assign mux_271_nl = MUX_s_1_2_2(mux_270_nl, mux_267_nl, act_config_inst_counter_sva[2]);
  assign mux_279_nl = MUX_s_1_2_2(mux_278_nl, mux_271_nl, act_config_inst_counter_sva[3]);
  assign mux_295_nl = MUX_s_1_2_2(mux_294_nl, mux_279_nl, act_config_inst_counter_sva[4]);
  assign and_1426_nl = is_start_sva & mux_295_nl;
  assign nor_nl = ~(is_start_sva | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11:9]!=3'b100)
      | (~(rva_in_PopNB_mioi_return_rsc_z_mxwt & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[8])
      & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)));
  assign mux_296_nl = MUX_s_1_2_2(and_1426_nl, nor_nl, fsm_output[1]);
  assign ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_13_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      rva_out_reg_data_159_128_sva_dfm_3, ActUnit_DecodeAxiRead_unequal_tmp_1);
  assign ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_12_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      rva_out_reg_data_191_160_sva_dfm_3, ActUnit_DecodeAxiRead_unequal_tmp_1);
  assign ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_11_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      rva_out_reg_data_223_192_sva_dfm_3, ActUnit_DecodeAxiRead_unequal_tmp_1);
  assign ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_10_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      rva_out_reg_data_255_224_sva_dfm_3, ActUnit_DecodeAxiRead_unequal_tmp_1);
  assign ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_9_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      rva_out_reg_data_287_256_sva_dfm_3, ActUnit_DecodeAxiRead_unequal_tmp_1);
  assign ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_8_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      rva_out_reg_data_319_288_sva_dfm_3, ActUnit_DecodeAxiRead_unequal_tmp_1);
  assign ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_7_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      rva_out_reg_data_351_320_sva_dfm_3, ActUnit_DecodeAxiRead_unequal_tmp_1);
  assign ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_6_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      rva_out_reg_data_383_352_sva_dfm_3, ActUnit_DecodeAxiRead_unequal_tmp_1);
  assign ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_5_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      rva_out_reg_data_415_384_sva_dfm_3, ActUnit_DecodeAxiRead_unequal_tmp_1);
  assign ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_4_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      rva_out_reg_data_447_416_sva_dfm_3, ActUnit_DecodeAxiRead_unequal_tmp_1);
  assign ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_3_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      rva_out_reg_data_479_448_sva_dfm_3, ActUnit_DecodeAxiRead_unequal_tmp_1);
  assign ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      rva_out_reg_data_511_480_sva_dfm_3, ActUnit_DecodeAxiRead_unequal_tmp_1);
  assign mux_252_nl = MUX_v_8_2_2(act_config_inst_regs_28_sva_dfm_6, act_config_inst_regs_12_sva_dfm_5,
      and_dcpl_916);
  assign not_1290_nl = ~ or_dcpl_639;
  assign and_1111_nl = MUX_v_8_2_2(8'b00000000, mux_252_nl, not_1290_nl);
  assign mux_253_nl = MUX_v_8_2_2(act_config_inst_regs_29_sva_dfm_6, act_config_inst_regs_13_sva_dfm_5,
      and_dcpl_916);
  assign not_1292_nl = ~ or_dcpl_639;
  assign and_1113_nl = MUX_v_8_2_2(8'b00000000, mux_253_nl, not_1292_nl);
  assign mux_254_nl = MUX_v_8_2_2(act_config_inst_regs_30_sva_dfm_6, act_config_inst_regs_14_sva_dfm_5,
      and_dcpl_916);
  assign not_1294_nl = ~ or_dcpl_639;
  assign and_1115_nl = MUX_v_8_2_2(8'b00000000, mux_254_nl, not_1294_nl);
  assign mux_255_nl = MUX_v_8_2_2(act_config_inst_regs_31_sva_dfm_6, act_config_inst_regs_15_sva_dfm_5,
      and_dcpl_916);
  assign not_1296_nl = ~ or_dcpl_639;
  assign and_1117_nl = MUX_v_8_2_2(8'b00000000, mux_255_nl, not_1296_nl);
  assign mux_256_nl = MUX_v_8_2_2(act_config_inst_regs_18_sva_dfm_6, act_config_inst_regs_2_sva_dfm_5,
      and_dcpl_916);
  assign not_1298_nl = ~ or_dcpl_639;
  assign and_1119_nl = MUX_v_8_2_2(8'b00000000, mux_256_nl, not_1298_nl);
  assign mux_257_nl = MUX_v_8_2_2(act_config_inst_regs_21_sva_dfm_6, act_config_inst_regs_5_sva_dfm_5,
      and_dcpl_916);
  assign not_1300_nl = ~ or_dcpl_639;
  assign and_1121_nl = MUX_v_8_2_2(8'b00000000, mux_257_nl, not_1300_nl);
  assign mux_258_nl = MUX_v_8_2_2(act_config_inst_regs_23_sva_dfm_6, act_config_inst_regs_7_sva_dfm_5,
      and_dcpl_916);
  assign not_1302_nl = ~ or_dcpl_639;
  assign and_1123_nl = MUX_v_8_2_2(8'b00000000, mux_258_nl, not_1302_nl);
  assign mux_259_nl = MUX_v_8_2_2(act_config_inst_regs_25_sva_dfm_6, act_config_inst_regs_9_sva_dfm_5,
      and_dcpl_916);
  assign not_1304_nl = ~ or_dcpl_639;
  assign and_1125_nl = MUX_v_8_2_2(8'b00000000, mux_259_nl, not_1304_nl);
  assign mux_260_nl = MUX_v_8_2_2(act_config_inst_regs_26_sva_dfm_6, act_config_inst_regs_10_sva_dfm_5,
      and_dcpl_916);
  assign not_1306_nl = ~ or_dcpl_639;
  assign and_1127_nl = MUX_v_8_2_2(8'b00000000, mux_260_nl, not_1306_nl);
  assign mux_261_nl = MUX_v_8_2_2(act_config_inst_regs_27_sva_dfm_6, act_config_inst_regs_11_sva_dfm_5,
      and_dcpl_916);
  assign not_1308_nl = ~ or_dcpl_639;
  assign and_1129_nl = MUX_v_8_2_2(8'b00000000, mux_261_nl, not_1308_nl);
  assign mux_262_nl = MUX_v_2_2_2((act_config_inst_regs_19_sva_dfm_6[7:6]), (act_config_inst_regs_3_sva_dfm_5[7:6]),
      and_dcpl_916);
  assign not_1310_nl = ~ or_dcpl_639;
  assign and_1131_nl = MUX_v_2_2_2(2'b00, mux_262_nl, not_1310_nl);
  assign mux_263_nl = MUX_v_7_2_2((act_config_inst_regs_17_sva_dfm_6[7:1]), (act_config_inst_regs_1_sva_dfm_5[7:1]),
      and_dcpl_916);
  assign not_1312_nl = ~ or_dcpl_639;
  assign and_1133_nl = MUX_v_7_2_2(7'b0000000, mux_263_nl, not_1312_nl);
  assign mux_264_nl = MUX_v_7_2_2((act_config_inst_regs_16_sva_dfm_6[7:1]), (act_config_inst_regs_0_sva_dfm_5[7:1]),
      and_dcpl_916);
  assign not_1314_nl = ~ or_dcpl_639;
  assign and_1135_nl = MUX_v_7_2_2(7'b0000000, mux_264_nl, not_1314_nl);
  assign mux_265_nl = MUX_v_3_2_2((act_config_inst_regs_22_sva_dfm_6[7:5]), (act_config_inst_regs_6_sva_dfm_5[7:5]),
      and_dcpl_916);
  assign not_1316_nl = ~ or_dcpl_639;
  assign and_1137_nl = MUX_v_3_2_2(3'b000, mux_265_nl, not_1316_nl);
  assign ActUnit_RunInst_switch_lp_mux_1_nl = MUX_s_1_2_2(ActUnit_RunInst_switch_lp_equal_tmp_1_mx0w0,
      ActUnit_RunInst_switch_lp_and_32_tmp, and_dcpl_557);
  assign ActUnit_RunInst_switch_lp_mux_2_nl = MUX_s_1_2_2(ActUnit_RunInst_switch_lp_equal_tmp_2_mx0w0,
      ActUnit_RunInst_switch_lp_equal_tmp_2, or_dcpl_442);
  assign ActUnit_RunInst_switch_lp_mux_4_nl = MUX_s_1_2_2(ActUnit_RunInst_switch_lp_equal_tmp_3_mx0w0,
      ActUnit_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva,
      and_dcpl_557);
  assign ActUnit_RunInst_switch_lp_mux_5_nl = MUX_s_1_2_2(ActUnit_RunInst_switch_lp_equal_tmp_4_mx0w0,
      ActUnit_RunInst_switch_lp_equal_tmp_4, or_dcpl_442);
  assign ActUnit_RunInst_switch_lp_mux_7_nl = MUX_s_1_2_2(ActUnit_RunInst_switch_lp_equal_tmp_5_mx0w0,
      ActUnit_RunInst_switch_lp_equal_tmp_5, or_dcpl_442);
  assign ActUnit_RunInst_switch_lp_mux_9_nl = MUX_s_1_2_2(ActUnit_RunInst_switch_lp_equal_tmp_6_mx0w0,
      ActUnit_RunInst_switch_lp_equal_tmp_6, or_dcpl_442);
  assign ActUnit_RunInst_switch_lp_mux_11_nl = MUX_s_1_2_2(ActUnit_RunInst_switch_lp_equal_tmp_7_mx0w0,
      ActUnit_RunInst_switch_lp_equal_tmp_7, or_dcpl_442);
  assign ActUnit_RunInst_switch_lp_mux_13_nl = MUX_s_1_2_2(ActUnit_RunInst_switch_lp_equal_tmp_8_mx0w0,
      ActUnit_RunInst_switch_lp_equal_tmp_8, or_dcpl_442);
  assign nv_scvector_cctor_nv_scvector_4_for_not_14_nl = ~ nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31;
  assign nv_scvector_cctor_nv_scvector_4_for_not_13_nl = ~ nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31;
  assign nv_scvector_cctor_nv_scvector_4_for_not_12_nl = ~ nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31;
  assign nv_scvector_cctor_nv_scvector_4_for_not_11_nl = ~ nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31;
  assign nv_scvector_cctor_nv_scvector_4_for_not_10_nl = ~ nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31;
  assign nv_scvector_cctor_nv_scvector_4_for_not_9_nl = ~ nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31;
  assign nv_scvector_cctor_nv_scvector_4_for_not_8_nl = ~ nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31;
  assign nv_scvector_cctor_nv_scvector_4_for_not_7_nl = ~ nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31;
  assign nv_scvector_cctor_nv_scvector_4_for_not_6_nl = ~ nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31;
  assign nv_scvector_cctor_nv_scvector_4_for_not_5_nl = ~ nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31;
  assign nv_scvector_cctor_nv_scvector_4_for_not_4_nl = ~ nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31;
  assign nv_scvector_cctor_nv_scvector_4_for_not_3_nl = ~ nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31;
  assign nv_scvector_cctor_nv_scvector_4_for_not_2_nl = ~ nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31;
  assign nv_scvector_cctor_nv_scvector_4_for_not_1_nl = ~ nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31;
  assign nv_scvector_cctor_nv_scvector_4_for_not_nl = ~ nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_slc_act_regs_data_32_31_0_1_ncse_sva_1_31;
  assign ActUnit_RunInst_switch_lp_not_1_nl = ~ ActUnit_RunInst_case_11_nv_scvector_cctor_data_0_sva_1_31;
  assign ActUnit_RunInst_switch_lp_or_3_nl = ActUnit_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva_mx0c3
      | and_dcpl_849;
  assign ActUnit_PushOutput_if_for_i_not_nl = ~ ActUnit_PushOutput_if_for_i_4_0_sva_3_0_mx0c0;
  assign nor_232_nl = ~((fsm_output[1:0]!=2'b01));
  assign mux_213_nl = MUX_s_1_2_2(nor_139_cse, nor_232_nl, fsm_output[4]);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_68_nl = act_regs_data_0_9_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_67_0;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_141_nl = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      act_regs_data_0_9_sva_dfm_2_30_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_67_0);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_4_nl = act_regs_data_1_0_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_71_0;
  assign act_regs_data_mux1h_74_nl = MUX1HOT_s_1_4_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_31,
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_4_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_0_1_sva_dfm_2_31, {and_dcpl_557 , and_dcpl_852 , act_regs_data_and_406_ssc
      , act_regs_data_and_407_ssc});
  assign act_regs_data_mux1h_575_nl = MUX1HOT_v_31_4_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_30_0,
      act_regs_data_1_0_sva_dfm_2_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
      act_regs_data_0_1_sva_dfm_2_30_0, {and_dcpl_557 , and_dcpl_852 , act_regs_data_and_406_ssc
      , act_regs_data_and_407_ssc});
  assign not_3696_nl = ~ or_dcpl_652;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_11_nl = act_regs_data_1_1_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_71_0;
  assign act_regs_data_mux1h_79_nl = MUX1HOT_s_1_4_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_31,
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_11_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_0_10_sva_dfm_2_31, {and_dcpl_557 , and_dcpl_852 , act_regs_data_and_408_ssc
      , act_regs_data_and_409_ssc});
  assign act_regs_data_mux1h_567_nl = MUX1HOT_v_31_4_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_30_0,
      act_regs_data_1_1_sva_dfm_2_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
      act_regs_data_0_10_sva_dfm_2_30_0, {and_dcpl_557 , and_dcpl_852 , act_regs_data_and_408_ssc
      , act_regs_data_and_409_ssc});
  assign not_3697_nl = ~ or_dcpl_652;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_73_nl = act_regs_data_1_10_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_71_0;
  assign act_regs_data_mux1h_84_nl = MUX1HOT_s_1_4_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_31,
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_73_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_0_11_sva_dfm_2_31, {and_dcpl_557 , and_dcpl_852 , act_regs_data_and_410_ssc
      , act_regs_data_and_411_ssc});
  assign act_regs_data_mux1h_566_nl = MUX1HOT_v_31_4_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_30_0,
      act_regs_data_1_10_sva_dfm_2_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
      act_regs_data_0_11_sva_dfm_2_30_0, {and_dcpl_557 , and_dcpl_852 , act_regs_data_and_410_ssc
      , act_regs_data_and_411_ssc});
  assign not_3698_nl = ~ or_dcpl_652;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_80_nl = act_regs_data_1_11_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_71_0;
  assign act_regs_data_mux1h_89_nl = MUX1HOT_s_1_4_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_31,
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_80_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_0_12_sva_dfm_2_31, {and_dcpl_557 , and_dcpl_852 , act_regs_data_and_412_ssc
      , act_regs_data_and_413_ssc});
  assign act_regs_data_mux1h_565_nl = MUX1HOT_v_31_4_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_30_0,
      act_regs_data_1_11_sva_dfm_2_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
      act_regs_data_0_12_sva_dfm_2_30_0, {and_dcpl_557 , and_dcpl_852 , act_regs_data_and_412_ssc
      , act_regs_data_and_413_ssc});
  assign not_3699_nl = ~ or_dcpl_652;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_87_nl = act_regs_data_1_12_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_71_0;
  assign act_regs_data_mux1h_94_nl = MUX1HOT_s_1_4_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_31,
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_87_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_0_13_sva_dfm_2_31, {and_dcpl_557 , and_dcpl_852 , act_regs_data_and_414_ssc
      , act_regs_data_and_415_ssc});
  assign act_regs_data_mux1h_564_nl = MUX1HOT_v_31_4_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_30_0,
      act_regs_data_1_12_sva_dfm_2_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
      act_regs_data_0_13_sva_dfm_2_30_0, {and_dcpl_557 , and_dcpl_852 , act_regs_data_and_414_ssc
      , act_regs_data_and_415_ssc});
  assign not_3700_nl = ~ or_dcpl_652;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_94_nl = act_regs_data_1_13_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_71_0;
  assign act_regs_data_mux1h_99_nl = MUX1HOT_s_1_4_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_31,
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_94_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_0_14_sva_dfm_2_31, {and_dcpl_557 , and_dcpl_852 , act_regs_data_and_416_ssc
      , act_regs_data_and_417_ssc});
  assign act_regs_data_mux1h_563_nl = MUX1HOT_v_31_4_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_30_0,
      act_regs_data_1_13_sva_dfm_2_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
      act_regs_data_0_14_sva_dfm_2_30_0, {and_dcpl_557 , and_dcpl_852 , act_regs_data_and_416_ssc
      , act_regs_data_and_417_ssc});
  assign not_3701_nl = ~ or_dcpl_652;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_101_nl = act_regs_data_1_14_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_71_0;
  assign act_regs_data_mux1h_104_nl = MUX1HOT_s_1_4_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_31,
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_101_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_0_15_sva_dfm_2_31, {and_dcpl_557 , and_dcpl_852 , act_regs_data_and_418_ssc
      , act_regs_data_and_419_ssc});
  assign act_regs_data_mux1h_562_nl = MUX1HOT_v_31_4_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_30_0,
      act_regs_data_1_14_sva_dfm_2_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
      act_regs_data_0_15_sva_dfm_2_30_0, {and_dcpl_557 , and_dcpl_852 , act_regs_data_and_418_ssc
      , act_regs_data_and_419_ssc});
  assign not_3702_nl = ~ or_dcpl_652;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_108_nl = act_regs_data_1_15_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_71_0;
  assign act_regs_data_mux1h_109_nl = MUX1HOT_s_1_4_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_31,
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_108_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_0_2_sva_dfm_2_31, {and_dcpl_557 , and_dcpl_852 , act_regs_data_and_420_ssc
      , act_regs_data_and_421_ssc});
  assign act_regs_data_mux1h_574_nl = MUX1HOT_v_31_4_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_30_0,
      act_regs_data_1_15_sva_dfm_2_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
      act_regs_data_0_2_sva_dfm_2_30_0, {and_dcpl_557 , and_dcpl_852 , act_regs_data_and_420_ssc
      , act_regs_data_and_421_ssc});
  assign not_3703_nl = ~ or_dcpl_652;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_18_nl = act_regs_data_1_2_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_71_0;
  assign act_regs_data_mux1h_114_nl = MUX1HOT_s_1_4_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_31,
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_18_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_0_3_sva_dfm_2_31, {and_dcpl_557 , and_dcpl_852 , act_regs_data_and_422_ssc
      , act_regs_data_and_423_ssc});
  assign act_regs_data_mux1h_573_nl = MUX1HOT_v_31_4_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_30_0,
      act_regs_data_1_2_sva_dfm_2_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
      act_regs_data_0_3_sva_dfm_2_30_0, {and_dcpl_557 , and_dcpl_852 , act_regs_data_and_422_ssc
      , act_regs_data_and_423_ssc});
  assign not_3704_nl = ~ or_dcpl_652;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_25_nl = act_regs_data_1_3_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_71_0;
  assign act_regs_data_mux1h_119_nl = MUX1HOT_s_1_4_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_31,
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_25_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_0_4_sva_dfm_2_31, {and_dcpl_557 , and_dcpl_852 , act_regs_data_and_424_ssc
      , act_regs_data_and_425_ssc});
  assign act_regs_data_mux1h_572_nl = MUX1HOT_v_31_4_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_30_0,
      act_regs_data_1_3_sva_dfm_2_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
      act_regs_data_0_4_sva_dfm_2_30_0, {and_dcpl_557 , and_dcpl_852 , act_regs_data_and_424_ssc
      , act_regs_data_and_425_ssc});
  assign not_3705_nl = ~ or_dcpl_652;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_32_nl = act_regs_data_1_4_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_71_0;
  assign act_regs_data_mux1h_124_nl = MUX1HOT_s_1_4_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_31,
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_32_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_0_5_sva_dfm_2_31, {and_dcpl_557 , and_dcpl_852 , act_regs_data_and_426_ssc
      , act_regs_data_and_427_ssc});
  assign act_regs_data_mux1h_571_nl = MUX1HOT_v_31_4_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_30_0,
      act_regs_data_1_4_sva_dfm_2_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
      act_regs_data_0_5_sva_dfm_2_30_0, {and_dcpl_557 , and_dcpl_852 , act_regs_data_and_426_ssc
      , act_regs_data_and_427_ssc});
  assign not_3706_nl = ~ or_dcpl_652;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_39_nl = act_regs_data_1_5_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_71_0;
  assign act_regs_data_mux1h_129_nl = MUX1HOT_s_1_4_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_31,
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_39_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_0_6_sva_dfm_2_31, {and_dcpl_557 , and_dcpl_852 , act_regs_data_and_428_ssc
      , act_regs_data_and_429_ssc});
  assign act_regs_data_mux1h_570_nl = MUX1HOT_v_31_4_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_30_0,
      act_regs_data_1_5_sva_dfm_2_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
      act_regs_data_0_6_sva_dfm_2_30_0, {and_dcpl_557 , and_dcpl_852 , act_regs_data_and_428_ssc
      , act_regs_data_and_429_ssc});
  assign not_3707_nl = ~ or_dcpl_652;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_46_nl = act_regs_data_1_6_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_71_0;
  assign act_regs_data_mux1h_134_nl = MUX1HOT_s_1_4_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_31,
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_46_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_0_7_sva_dfm_2_31, {and_dcpl_557 , and_dcpl_852 , act_regs_data_and_430_ssc
      , act_regs_data_and_431_ssc});
  assign act_regs_data_mux1h_569_nl = MUX1HOT_v_31_4_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_30_0,
      act_regs_data_1_6_sva_dfm_2_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
      act_regs_data_0_7_sva_dfm_2_30_0, {and_dcpl_557 , and_dcpl_852 , act_regs_data_and_430_ssc
      , act_regs_data_and_431_ssc});
  assign not_3708_nl = ~ or_dcpl_652;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_53_nl = act_regs_data_1_7_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_71_0;
  assign act_regs_data_mux1h_139_nl = MUX1HOT_s_1_4_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_31,
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_53_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_0_8_sva_dfm_2_31, {and_dcpl_557 , and_dcpl_852 , act_regs_data_and_432_ssc
      , act_regs_data_and_433_ssc});
  assign act_regs_data_mux1h_568_nl = MUX1HOT_v_31_4_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_30_0,
      act_regs_data_1_7_sva_dfm_2_30_0, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:0]),
      act_regs_data_0_8_sva_dfm_2_30_0, {and_dcpl_557 , and_dcpl_852 , act_regs_data_and_432_ssc
      , act_regs_data_and_433_ssc});
  assign not_3709_nl = ~ or_dcpl_652;
  assign ActUnit_RunInst_case_2_for_ActUnit_RunInst_case_2_for_and_nl = ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_31
      & ActUnit_RunInst_case_2_for_and_27_seb;
  assign Gelu_for_Gelu_for_and_11_nl = (z_out_28_1[27]) & (~ Gelu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & (~ Gelu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_6_nl = act_regs_data_0_0_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_67_0;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_and_34_nl = (~ Gelu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & and_dcpl_900;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_and_35_nl = Gelu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & and_dcpl_900;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_90_nl = MUX1HOT_v_31_5_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_30_0,
      ({{3{z_out_28_1[27]}}, z_out_28_1}), nv_scvector_cctor_nv_scvector_6_for_12_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0,
      ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_2_30_0, act_regs_data_0_0_sva_dfm_2_30_0,
      {and_dcpl_557 , ActUnit_PushOutput_if_output_port_reg_data_data_and_34_nl ,
      ActUnit_PushOutput_if_output_port_reg_data_data_and_35_nl , and_dcpl_832 ,
      and_dcpl_852});
  assign nor_771_nl = ~(and_dcpl_1229 | (Gelu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
      & and_dcpl_900) | ((~ ActUnit_RunInst_case_2_for_and_27_seb) & and_dcpl_557));
  assign nor_340_nl = ~(and_dcpl_906 | or_996_tmp);
  assign and_1140_nl = and_dcpl_906 & (~ or_996_tmp);
  assign mux_217_nl = MUX_s_1_2_2((~ or_tmp_317), or_1097_cse, fsm_output[4]);
  assign ActUnit_DecodeAxiRead_else_mux_1_nl = MUX_s_1_2_2(ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0,
      ActUnit_DecodeAxiRead_else_unequal_tmp, or_dcpl_301);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_5_nl = (~ ActUnit_DecodeAxiRead_else_mux_1_nl)
      & ActUnit_DecodeAxiRead_unequal_tmp_1 & (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      & rva_in_PopNB_mioi_return_rsc_z_mxwt;
  assign act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_24_nl
      = act_config_inst_regs_16_sva_0 & act_config_ActConfigRead_else_else_not_21;
  assign act_config_ActConfigRead_else_mux_19_nl = MUX_s_1_2_2(act_config_inst_regs_0_sva_0,
      act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_24_nl,
      act_config_ActConfigRead_else_unequal_tmp_1);
  assign act_config_ActConfigRead_mux_19_nl = MUX_s_1_2_2(act_config_is_valid_sva,
      act_config_ActConfigRead_else_mux_19_nl, act_config_ActConfigRead_unequal_tmp_1);
  assign ActUnit_DecodeAxiRead_mux_33_nl = MUX_s_1_2_2(act_config_ActConfigRead_mux_19_nl,
      ActUnit_PushOutput_if_for_and_stg_2_7_sva, ActUnit_DecodeAxiRead_unequal_tmp_1);
  assign ActUnit_DecodeAxi_if_mux_91_nl = MUX_s_1_2_2(ActUnit_DecodeAxiRead_mux_33_nl,
      ActUnit_PushOutput_if_for_and_stg_2_7_sva, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt);
  assign ActUnit_DecodeAxi_mux_93_nl = MUX_s_1_2_2(ActUnit_PushOutput_if_for_and_stg_2_7_sva,
      ActUnit_DecodeAxi_if_mux_91_nl, rva_in_PopNB_mioi_return_rsc_z_mxwt);
  assign act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_18_nl
      = act_config_inst_regs_17_sva_0 & act_config_ActConfigRead_else_else_not_21;
  assign act_config_ActConfigRead_else_mux_17_nl = MUX_s_1_2_2(act_config_inst_regs_1_sva_0,
      act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_18_nl,
      act_config_ActConfigRead_else_unequal_tmp_1);
  assign act_config_ActConfigRead_mux_17_nl = MUX_s_1_2_2(act_config_is_zero_first_sva,
      act_config_ActConfigRead_else_mux_17_nl, act_config_ActConfigRead_unequal_tmp_1);
  assign ActUnit_DecodeAxiRead_mux_31_nl = MUX_s_1_2_2(act_config_ActConfigRead_mux_17_nl,
      Gelu_for_and_2_cse_sva, ActUnit_DecodeAxiRead_unequal_tmp_1);
  assign ActUnit_DecodeAxi_if_mux_89_nl = MUX_s_1_2_2(ActUnit_DecodeAxiRead_mux_31_nl,
      Gelu_for_and_2_cse_sva, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt);
  assign ActUnit_DecodeAxi_mux_94_nl = MUX_s_1_2_2(Gelu_for_and_2_cse_sva, ActUnit_DecodeAxi_if_mux_89_nl,
      rva_in_PopNB_mioi_return_rsc_z_mxwt);
  assign act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_20_nl
      = MUX_v_6_2_2(6'b000000, (act_config_inst_regs_19_sva_dfm_6[5:0]), act_config_ActConfigRead_else_else_not_21);
  assign act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_21_nl
      = MUX_v_8_2_2(8'b00000000, act_config_inst_regs_20_sva_dfm_6, act_config_ActConfigRead_else_else_not_21);
  assign act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_22_nl
      = MUX_v_5_2_2(5'b00000, (act_config_inst_regs_22_sva_dfm_6[4:0]), act_config_ActConfigRead_else_else_not_21);
  assign act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_23_nl
      = MUX_v_8_2_2(8'b00000000, act_config_inst_regs_24_sva_dfm_6, act_config_ActConfigRead_else_else_not_21);
  assign or_997_nl = and_dcpl_908 | ActUnit_DecodeAxiRead_unequal_tmp_1;
  assign act_config_ActConfigWrite_mux_1_nl = MUX_s_1_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[8]),
      act_config_is_zero_first_sva, act_config_ActConfigRead_unequal_tmp_1);
  assign ActUnit_DecodeAxiWrite_mux_4_nl = MUX_s_1_2_2(act_config_ActConfigWrite_mux_1_nl,
      act_config_is_zero_first_sva, ActUnit_DecodeAxiRead_unequal_tmp_1);
  assign ActUnit_DecodeAxiWrite_if_mux_5_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[3:2]),
      (act_config_inst_regs_16_sva_dfm_6[3:2]), not_tmp_347);
  assign ActUnit_DecodeAxiWrite_if_mux_7_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[11:10]),
      (act_config_inst_regs_17_sva_dfm_6[3:2]), not_tmp_347);
  assign ActUnit_DecodeAxiWrite_if_mux_9_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[19:18]),
      (act_config_inst_regs_18_sva_dfm_6[3:2]), not_tmp_347);
  assign ActUnit_DecodeAxiWrite_if_mux_11_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[27:26]),
      (act_config_inst_regs_19_sva_dfm_6[3:2]), not_tmp_347);
  assign ActUnit_DecodeAxiWrite_if_mux_13_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[35:34]),
      (act_config_inst_regs_20_sva_dfm_6[3:2]), not_tmp_347);
  assign ActUnit_DecodeAxiWrite_if_mux_15_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[43:42]),
      (act_config_inst_regs_21_sva_dfm_6[3:2]), not_tmp_347);
  assign ActUnit_DecodeAxiWrite_if_mux_17_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[51:50]),
      (act_config_inst_regs_22_sva_dfm_6[3:2]), not_tmp_347);
  assign ActUnit_DecodeAxiWrite_if_mux_19_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[59:58]),
      (act_config_inst_regs_23_sva_dfm_6[3:2]), not_tmp_347);
  assign ActUnit_DecodeAxiWrite_if_mux_21_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[67:66]),
      (act_config_inst_regs_24_sva_dfm_6[3:2]), not_tmp_347);
  assign ActUnit_DecodeAxiWrite_if_mux_23_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[75:74]),
      (act_config_inst_regs_25_sva_dfm_6[3:2]), not_tmp_347);
  assign ActUnit_DecodeAxiWrite_if_mux_25_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[83:82]),
      (act_config_inst_regs_26_sva_dfm_6[3:2]), not_tmp_347);
  assign ActUnit_DecodeAxiWrite_if_mux_27_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[91:90]),
      (act_config_inst_regs_27_sva_dfm_6[3:2]), not_tmp_347);
  assign ActUnit_DecodeAxiWrite_if_mux_29_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[99:98]),
      (act_config_inst_regs_28_sva_dfm_6[3:2]), not_tmp_347);
  assign ActUnit_DecodeAxiWrite_if_mux_31_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[107:106]),
      (act_config_inst_regs_29_sva_dfm_6[3:2]), not_tmp_347);
  assign ActUnit_DecodeAxiWrite_if_mux_33_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[115:114]),
      (act_config_inst_regs_30_sva_dfm_6[3:2]), not_tmp_347);
  assign ActUnit_DecodeAxiWrite_if_mux_35_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[123:122]),
      (act_config_inst_regs_31_sva_dfm_6[3:2]), not_tmp_347);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_69_nl = act_regs_data_3_9_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_65_0;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_174_nl = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      act_regs_data_3_9_sva_dfm_2_30_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_65_0);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_104_nl = act_regs_data_3_14_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_65_0;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_173_nl = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      act_regs_data_3_14_sva_dfm_2_30_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_65_0);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_97_nl = act_regs_data_3_13_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_65_0;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_171_nl = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      act_regs_data_3_13_sva_dfm_2_30_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_65_0);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_90_nl = act_regs_data_3_12_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_65_0;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_169_nl = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      act_regs_data_3_12_sva_dfm_2_30_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_65_0);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_83_nl = act_regs_data_3_11_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_65_0;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_167_nl = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      act_regs_data_3_11_sva_dfm_2_30_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_65_0);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_76_nl = act_regs_data_3_10_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_65_0;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_165_nl = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      act_regs_data_3_10_sva_dfm_2_30_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_65_0);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_12_nl = act_regs_data_3_1_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_65_0;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_163_nl = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      act_regs_data_3_1_sva_dfm_2_30_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_65_0);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_62_nl = act_regs_data_3_8_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_65_0;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_161_nl = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      act_regs_data_3_8_sva_dfm_2_30_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_65_0);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_54_nl = act_regs_data_3_7_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_65_0;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_159_nl = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      act_regs_data_3_7_sva_dfm_2_30_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_65_0);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_47_nl = act_regs_data_3_6_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_65_0;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_157_nl = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      act_regs_data_3_6_sva_dfm_2_30_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_65_0);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_40_nl = act_regs_data_3_5_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_65_0;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_155_nl = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      act_regs_data_3_5_sva_dfm_2_30_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_65_0);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_33_nl = act_regs_data_3_4_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_65_0;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_153_nl = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      act_regs_data_3_4_sva_dfm_2_30_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_65_0);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_26_nl = act_regs_data_3_3_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_65_0;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_151_nl = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      act_regs_data_3_3_sva_dfm_2_30_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_65_0);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_19_nl = act_regs_data_3_2_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_65_0;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_149_nl = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      act_regs_data_3_2_sva_dfm_2_30_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_65_0);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_111_nl = act_regs_data_3_15_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_65_0;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_147_nl = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      act_regs_data_3_15_sva_dfm_2_30_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_65_0);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_5_nl = act_regs_data_3_0_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_65_0;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_145_nl = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      act_regs_data_3_0_sva_dfm_2_30_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_65_0);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_67_nl = act_regs_data_2_9_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_69_0;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_143_nl = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      act_regs_data_2_9_sva_dfm_2_30_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_69_0);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_102_nl = act_regs_data_2_14_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_69_0;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_142_nl = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      act_regs_data_2_14_sva_dfm_2_30_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_69_0);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_95_nl = act_regs_data_2_13_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_69_0;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_144_nl = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      act_regs_data_2_13_sva_dfm_2_30_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_69_0);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_88_nl = act_regs_data_2_12_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_69_0;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_146_nl = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      act_regs_data_2_12_sva_dfm_2_30_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_69_0);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_81_nl = act_regs_data_2_11_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_69_0;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_148_nl = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      act_regs_data_2_11_sva_dfm_2_30_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_69_0);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_74_nl = act_regs_data_2_10_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_69_0;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_150_nl = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      act_regs_data_2_10_sva_dfm_2_30_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_69_0);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_10_nl = act_regs_data_2_1_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_69_0;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_152_nl = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      act_regs_data_2_1_sva_dfm_2_30_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_69_0);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_60_nl = act_regs_data_2_8_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_69_0;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_154_nl = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      act_regs_data_2_8_sva_dfm_2_30_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_69_0);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_52_nl = act_regs_data_2_7_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_69_0;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_156_nl = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      act_regs_data_2_7_sva_dfm_2_30_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_69_0);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_45_nl = act_regs_data_2_6_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_69_0;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_158_nl = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      act_regs_data_2_6_sva_dfm_2_30_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_69_0);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_38_nl = act_regs_data_2_5_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_69_0;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_160_nl = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      act_regs_data_2_5_sva_dfm_2_30_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_69_0);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_31_nl = act_regs_data_2_4_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_69_0;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_162_nl = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      act_regs_data_2_4_sva_dfm_2_30_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_69_0);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_24_nl = act_regs_data_2_3_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_69_0;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_164_nl = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      act_regs_data_2_3_sva_dfm_2_30_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_69_0);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_17_nl = act_regs_data_2_2_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_69_0;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_166_nl = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      act_regs_data_2_2_sva_dfm_2_30_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_69_0);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_109_nl = act_regs_data_2_15_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_69_0;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_168_nl = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      act_regs_data_2_15_sva_dfm_2_30_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_69_0);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_3_nl = act_regs_data_2_0_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_69_0;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_170_nl = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      act_regs_data_2_0_sva_dfm_2_30_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_69_0);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_66_nl = act_regs_data_1_9_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_71_0;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_172_nl = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      act_regs_data_1_9_sva_dfm_2_30_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_71_0);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_59_nl = act_regs_data_1_8_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_71_0;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_175_nl = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      act_regs_data_1_8_sva_dfm_2_30_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_71_0);
  assign ActUnit_DecodeAxiRead_else_mux_3_nl = MUX_s_1_2_2(ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0,
      ActUnit_DecodeAxiWrite_else_unequal_tmp, or_dcpl_304);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_23_nl = (~ ActUnit_DecodeAxiRead_else_mux_3_nl)
      & ActUnit_DecodeAxiRead_unequal_tmp_1 & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & rva_in_PopNB_mioi_return_rsc_z_mxwt;
  assign while_and_64_nl = act_config_InstIncr_act_config_InstIncr_if_and_svs_1 &
      is_incr_lpi_1_dfm_1 & is_start_sva;
  assign Silu_for_else_mux_1_nl = MUX_v_31_2_2(({{2{z_out_3_29_1[28]}}, z_out_3_29_1}),
      nv_scvector_cctor_nv_scvector_5_for_2_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0,
      Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs);
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_not_34_nl = ~ Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs;
  assign Silu_for_Silu_for_and_nl = (Silu_for_1_else_else_acc_itm_29_1[28]) & (~
      Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      & (~ Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_48_nl = act_regs_data_0_6_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_67_0;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_10_nl = MUX1HOT_s_1_3_2(Silu_for_Silu_for_and_nl,
      ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_2_31, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_48_nl,
      {and_dcpl_592 , and_dcpl_832 , and_dcpl_852});
  assign mux_222_nl = MUX_s_1_2_2((~ (fsm_output[3])), (fsm_output[3]), and_1046_cse);
  assign mux_223_nl = MUX_s_1_2_2(mux_222_nl, or_1097_cse, fsm_output[4]);
  assign ActUnit_PushOutput_if_output_port_reg_data_data_and_36_nl = (~ Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      & and_dcpl_592;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_and_37_nl = Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
      & and_dcpl_592;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_83_nl = MUX1HOT_v_31_4_2(({{2{Silu_for_1_else_else_acc_itm_29_1[28]}},
      Silu_for_1_else_else_acc_itm_29_1}), ActUnit_RunInst_case_14_nv_scvector_cctor_data_0_sva_30_0,
      ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_2_30_0, act_regs_data_0_6_sva_dfm_2_30_0,
      {ActUnit_PushOutput_if_output_port_reg_data_data_and_36_nl , ActUnit_PushOutput_if_output_port_reg_data_data_and_37_nl
      , and_dcpl_832 , and_dcpl_852});
  assign nor_772_nl = ~(or_dcpl_655 | (and_dcpl_592 & Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs));
  assign Silu_for_else_mux_3_nl = MUX_v_31_2_2(({{2{z_out_4_29_1[28]}}, z_out_4_29_1}),
      nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0,
      Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs);
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_not_36_nl = ~ Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs;
  assign Silu_for_else_mux_2_nl = MUX_v_31_2_2(({{2{z_out_3_29_1[28]}}, z_out_3_29_1}),
      nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0,
      Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs);
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_not_35_nl = ~ Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs;
  assign Silu_for_else_mux_5_nl = MUX_v_31_2_2(({{2{z_out_4_29_1[28]}}, z_out_4_29_1}),
      nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0,
      Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs);
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_not_38_nl = ~ Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs;
  assign Silu_for_else_mux_4_nl = MUX_v_31_2_2(({{2{z_out_3_29_1[28]}}, z_out_3_29_1}),
      nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0,
      Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs);
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_not_37_nl = ~ Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs;
  assign or_993_nl = (fsm_output[0]) | (fsm_output[2]) | (~ (fsm_output[3]));
  assign or_994_nl = (~ (fsm_output[0])) | (~ (fsm_output[2])) | (fsm_output[3]);
  assign mux_227_nl = MUX_s_1_2_2(or_993_nl, or_994_nl, fsm_output[1]);
  assign Silu_for_else_mux_7_nl = MUX_v_31_2_2(({{2{z_out_3_29_1[28]}}, z_out_3_29_1}),
      nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0,
      Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs);
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_not_40_nl = ~ Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs;
  assign Silu_for_else_mux_6_nl = MUX_v_31_2_2(({{2{z_out_4_29_1[28]}}, z_out_4_29_1}),
      nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0,
      Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs);
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_not_39_nl = ~ Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs;
  assign Silu_for_else_mux_8_nl = MUX_v_31_2_2(({{2{z_out_4_29_1[28]}}, z_out_4_29_1}),
      nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0,
      Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs);
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_not_41_nl = ~ Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs;
  assign Gelu_for_Gelu_for_and_1_nl = (z_out_1_28_1[27]) & (~ Gelu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & (~ Gelu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_89_nl = act_regs_data_0_12_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_67_0;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_15_nl = MUX1HOT_s_1_3_2(Gelu_for_Gelu_for_and_1_nl,
      ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_2_31, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_89_nl,
      {and_dcpl_576 , and_dcpl_832 , and_dcpl_852});
  assign ActUnit_PushOutput_if_output_port_reg_data_data_and_38_nl = (~ Gelu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & and_dcpl_576;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_and_39_nl = Gelu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & and_dcpl_576;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_78_nl = MUX1HOT_v_31_4_2(({{3{z_out_1_28_1[27]}},
      z_out_1_28_1}), nv_scvector_cctor_nv_scvector_6_for_2_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0,
      ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_2_30_0, act_regs_data_0_12_sva_dfm_2_30_0,
      {ActUnit_PushOutput_if_output_port_reg_data_data_and_38_nl , ActUnit_PushOutput_if_output_port_reg_data_data_and_39_nl
      , and_dcpl_832 , and_dcpl_852});
  assign nor_773_nl = ~(or_dcpl_655 | (Gelu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
      & and_dcpl_576));
  assign Silu_for_Silu_for_and_9_nl = (z_out_3_29_1[28]) & (~ Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      & (~ Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_55_nl = act_regs_data_0_7_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_67_0;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_20_nl = MUX1HOT_s_1_3_2(Silu_for_Silu_for_and_9_nl,
      ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_2_31, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_55_nl,
      {and_dcpl_576 , and_dcpl_832 , and_dcpl_852});
  assign ActUnit_PushOutput_if_output_port_reg_data_data_and_40_nl = (~ Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      & and_dcpl_576;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_and_41_nl = Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
      & and_dcpl_576;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_82_nl = MUX1HOT_v_31_4_2(({{2{z_out_3_29_1[28]}},
      z_out_3_29_1}), nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0,
      ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_2_30_0, act_regs_data_0_7_sva_dfm_2_30_0,
      {ActUnit_PushOutput_if_output_port_reg_data_data_and_40_nl , ActUnit_PushOutput_if_output_port_reg_data_data_and_41_nl
      , and_dcpl_832 , and_dcpl_852});
  assign nor_774_nl = ~(or_dcpl_655 | (and_dcpl_576 & Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs));
  assign Gelu_for_Gelu_for_and_nl = (z_out_2_28_1[27]) & (~ Gelu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & (~ Gelu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs);
  assign Gelu_for_else_mux_nl = MUX_v_31_2_2(({{3{z_out_2_28_1[27]}}, z_out_2_28_1}),
      ActUnit_RunInst_case_15_nv_scvector_cctor_data_0_sva_30_0, Gelu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs);
  assign operator_32_8_true_AC_TRN_AC_WRAP_3_not_34_nl = ~ Gelu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs;
  assign Gelu_for_Gelu_for_and_19_nl = MUX_v_31_2_2(31'b0000000000000000000000000000000,
      Gelu_for_else_mux_nl, operator_32_8_true_AC_TRN_AC_WRAP_3_not_34_nl);
  assign Silu_for_else_mux_11_nl = MUX_v_31_2_2(({{2{z_out_3_29_1[28]}}, z_out_3_29_1}),
      nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0,
      Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs);
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_not_42_nl = ~ Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs;
  assign Gelu_for_Gelu_for_and_2_nl = (z_out_1_28_1[27]) & (~ Gelu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & (~ Gelu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_96_nl = act_regs_data_0_13_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_67_0;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_25_nl = MUX1HOT_s_1_3_2(Gelu_for_Gelu_for_and_2_nl,
      ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_2_31, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_96_nl,
      {and_dcpl_578 , and_dcpl_832 , and_dcpl_852});
  assign ActUnit_PushOutput_if_output_port_reg_data_data_and_42_nl = (~ Gelu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & and_dcpl_578;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_and_43_nl = Gelu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & and_dcpl_578;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_77_nl = MUX1HOT_v_31_4_2(({{3{z_out_1_28_1[27]}},
      z_out_1_28_1}), nv_scvector_cctor_nv_scvector_6_for_3_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0,
      ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_2_30_0, act_regs_data_0_13_sva_dfm_2_30_0,
      {ActUnit_PushOutput_if_output_port_reg_data_data_and_42_nl , ActUnit_PushOutput_if_output_port_reg_data_data_and_43_nl
      , and_dcpl_832 , and_dcpl_852});
  assign nor_775_nl = ~(or_dcpl_655 | (Gelu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
      & and_dcpl_578));
  assign Silu_for_Silu_for_and_10_nl = (z_out_4_29_1[28]) & (~ Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      & (~ Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_61_nl = act_regs_data_0_8_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_67_0;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_30_nl = MUX1HOT_s_1_3_2(Silu_for_Silu_for_and_10_nl,
      ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_2_31, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_61_nl,
      {and_dcpl_578 , and_dcpl_832 , and_dcpl_852});
  assign ActUnit_PushOutput_if_output_port_reg_data_data_and_44_nl = (~ Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      & and_dcpl_578;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_and_45_nl = Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
      & and_dcpl_578;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_81_nl = MUX1HOT_v_31_4_2(({{2{z_out_4_29_1[28]}},
      z_out_4_29_1}), nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0,
      ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_2_30_0, act_regs_data_0_8_sva_dfm_2_30_0,
      {ActUnit_PushOutput_if_output_port_reg_data_data_and_44_nl , ActUnit_PushOutput_if_output_port_reg_data_data_and_45_nl
      , and_dcpl_832 , and_dcpl_852});
  assign nor_776_nl = ~(or_dcpl_655 | (and_dcpl_578 & Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs));
  assign Silu_for_else_mux_13_nl = MUX_v_31_2_2(({{2{z_out_3_29_1[28]}}, z_out_3_29_1}),
      nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0,
      Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs);
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_not_44_nl = ~ Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs;
  assign Silu_for_else_mux_12_nl = MUX_v_31_2_2(({{2{z_out_4_29_1[28]}}, z_out_4_29_1}),
      nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0,
      Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs);
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_not_43_nl = ~ Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs;
  assign Gelu_for_Gelu_for_and_3_nl = (z_out_1_28_1[27]) & (~ Gelu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & (~ Gelu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_103_nl = act_regs_data_0_14_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_67_0;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_35_nl = MUX1HOT_s_1_3_2(Gelu_for_Gelu_for_and_3_nl,
      ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_2_31, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_103_nl,
      {and_dcpl_1006 , and_dcpl_832 , and_dcpl_852});
  assign ActUnit_PushOutput_if_output_port_reg_data_data_and_46_nl = (~ Gelu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & and_dcpl_1006;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_and_47_nl = Gelu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & and_dcpl_1006;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_76_nl = MUX1HOT_v_31_4_2(({{3{z_out_1_28_1[27]}},
      z_out_1_28_1}), nv_scvector_cctor_nv_scvector_6_for_4_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0,
      ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_2_30_0, act_regs_data_0_14_sva_dfm_2_30_0,
      {ActUnit_PushOutput_if_output_port_reg_data_data_and_46_nl , ActUnit_PushOutput_if_output_port_reg_data_data_and_47_nl
      , and_dcpl_832 , and_dcpl_852});
  assign nor_777_nl = ~(or_dcpl_655 | (Gelu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs
      & and_dcpl_1006));
  assign Gelu_for_Gelu_for_and_4_nl = (z_out_2_28_1[27]) & (~ Gelu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & (~ Gelu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_110_nl = act_regs_data_0_15_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_67_0;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_40_nl = MUX1HOT_s_1_3_2(Gelu_for_Gelu_for_and_4_nl,
      ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_2_31, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_110_nl,
      {and_dcpl_1006 , and_dcpl_832 , and_dcpl_852});
  assign ActUnit_PushOutput_if_output_port_reg_data_data_and_48_nl = (~ Gelu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & and_dcpl_1006;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_and_49_nl = Gelu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & and_dcpl_1006;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_88_nl = MUX1HOT_v_31_4_2(({{3{z_out_2_28_1[27]}},
      z_out_2_28_1}), nv_scvector_cctor_nv_scvector_6_for_5_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0,
      ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_2_30_0, act_regs_data_0_15_sva_dfm_2_30_0,
      {ActUnit_PushOutput_if_output_port_reg_data_data_and_48_nl , ActUnit_PushOutput_if_output_port_reg_data_data_and_49_nl
      , and_dcpl_832 , and_dcpl_852});
  assign nor_778_nl = ~(or_dcpl_655 | (and_dcpl_1006 & Gelu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs));
  assign Silu_for_else_mux_15_nl = MUX_v_31_2_2(({{2{z_out_3_29_1[28]}}, z_out_3_29_1}),
      nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0,
      Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs);
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_not_46_nl = ~ Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs;
  assign Silu_for_else_mux_14_nl = MUX_v_31_2_2(({{2{z_out_4_29_1[28]}}, z_out_4_29_1}),
      nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0,
      Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs);
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_not_45_nl = ~ Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_7_svs;
  assign Gelu_for_Gelu_for_and_5_nl = (z_out_1_28_1[27]) & (~ Gelu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & (~ Gelu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_20_nl = act_regs_data_0_2_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_67_0;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_45_nl = MUX1HOT_s_1_3_2(Gelu_for_Gelu_for_and_5_nl,
      ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_2_31, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_20_nl,
      {and_dcpl_900 , and_dcpl_832 , and_dcpl_852});
  assign ActUnit_PushOutput_if_output_port_reg_data_data_and_50_nl = (~ Gelu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & and_dcpl_900;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_and_51_nl = Gelu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & and_dcpl_900;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_87_nl = MUX1HOT_v_31_4_2(({{3{z_out_1_28_1[27]}},
      z_out_1_28_1}), nv_scvector_cctor_nv_scvector_6_for_6_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0,
      ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_2_30_0, act_regs_data_0_2_sva_dfm_2_30_0,
      {ActUnit_PushOutput_if_output_port_reg_data_data_and_50_nl , ActUnit_PushOutput_if_output_port_reg_data_data_and_51_nl
      , and_dcpl_832 , and_dcpl_852});
  assign nor_779_nl = ~(or_dcpl_655 | (and_dcpl_900 & Gelu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs));
  assign Gelu_for_Gelu_for_and_6_nl = (z_out_2_28_1[27]) & (~ Gelu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & (~ Gelu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_27_nl = act_regs_data_0_3_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_67_0;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_50_nl = MUX1HOT_s_1_3_2(Gelu_for_Gelu_for_and_6_nl,
      ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_2_31, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_27_nl,
      {and_dcpl_900 , and_dcpl_832 , and_dcpl_852});
  assign ActUnit_PushOutput_if_output_port_reg_data_data_and_52_nl = (~ Gelu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & and_dcpl_900;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_and_53_nl = Gelu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & and_dcpl_900;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_86_nl = MUX1HOT_v_31_4_2(({{3{z_out_2_28_1[27]}},
      z_out_2_28_1}), nv_scvector_cctor_nv_scvector_6_for_7_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0,
      ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_2_30_0, act_regs_data_0_3_sva_dfm_2_30_0,
      {ActUnit_PushOutput_if_output_port_reg_data_data_and_52_nl , ActUnit_PushOutput_if_output_port_reg_data_data_and_53_nl
      , and_dcpl_832 , and_dcpl_852});
  assign nor_780_nl = ~(or_dcpl_655 | (and_dcpl_900 & Gelu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs));
  assign Gelu_for_Gelu_for_and_12_nl = (Gelu_for_13_else_else_acc_itm_28_1[27]) &
      (~ Gelu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & (~ Gelu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_13_nl = act_regs_data_0_1_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_67_0;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_55_nl = MUX1HOT_s_1_3_2(Gelu_for_Gelu_for_and_12_nl,
      ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_2_31, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_13_nl,
      {and_dcpl_1007 , and_dcpl_832 , and_dcpl_852});
  assign ActUnit_PushOutput_if_output_port_reg_data_data_and_54_nl = (~ Gelu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & and_dcpl_1007;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_and_55_nl = Gelu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & and_dcpl_1007;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_89_nl = MUX1HOT_v_31_4_2(({{3{Gelu_for_13_else_else_acc_itm_28_1[27]}},
      Gelu_for_13_else_else_acc_itm_28_1}), nv_scvector_cctor_nv_scvector_6_for_13_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0,
      ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_2_30_0, act_regs_data_0_1_sva_dfm_2_30_0,
      {ActUnit_PushOutput_if_output_port_reg_data_data_and_54_nl , ActUnit_PushOutput_if_output_port_reg_data_data_and_55_nl
      , and_dcpl_832 , and_dcpl_852});
  assign nor_781_nl = ~(or_dcpl_655 | (and_dcpl_1007 & Gelu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs));
  assign Gelu_for_Gelu_for_and_13_nl = (z_out_2_28_1[27]) & (~ Gelu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & (~ Gelu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_75_nl = act_regs_data_0_10_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_67_0;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_60_nl = MUX1HOT_s_1_3_2(Gelu_for_Gelu_for_and_13_nl,
      ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_2_31, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_75_nl,
      {and_dcpl_1007 , and_dcpl_832 , and_dcpl_852});
  assign ActUnit_PushOutput_if_output_port_reg_data_data_and_56_nl = (~ Gelu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & and_dcpl_1007;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_and_57_nl = Gelu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & and_dcpl_1007;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_80_nl = MUX1HOT_v_31_4_2(({{3{z_out_2_28_1[27]}},
      z_out_2_28_1}), nv_scvector_cctor_nv_scvector_6_for_14_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0,
      ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_2_30_0, act_regs_data_0_10_sva_dfm_2_30_0,
      {ActUnit_PushOutput_if_output_port_reg_data_data_and_56_nl , ActUnit_PushOutput_if_output_port_reg_data_data_and_57_nl
      , and_dcpl_832 , and_dcpl_852});
  assign nor_782_nl = ~(or_dcpl_655 | (and_dcpl_1007 & Gelu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs));
  assign Gelu_for_Gelu_for_and_14_nl = (z_out_1_28_1[27]) & (~ Gelu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & (~ Gelu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_82_nl = act_regs_data_0_11_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_67_0;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_65_nl = MUX1HOT_s_1_3_2(Gelu_for_Gelu_for_and_14_nl,
      ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_2_31, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_82_nl,
      {and_dcpl_1007 , and_dcpl_832 , and_dcpl_852});
  assign ActUnit_PushOutput_if_output_port_reg_data_data_and_58_nl = (~ Gelu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & and_dcpl_1007;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_and_59_nl = Gelu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & and_dcpl_1007;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_79_nl = MUX1HOT_v_31_4_2(({{3{z_out_1_28_1[27]}},
      z_out_1_28_1}), nv_scvector_cctor_nv_scvector_6_for_15_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0,
      ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_2_30_0, act_regs_data_0_11_sva_dfm_2_30_0,
      {ActUnit_PushOutput_if_output_port_reg_data_data_and_58_nl , ActUnit_PushOutput_if_output_port_reg_data_data_and_59_nl
      , and_dcpl_832 , and_dcpl_852});
  assign nor_783_nl = ~(or_dcpl_655 | (and_dcpl_1007 & Gelu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs));
  assign Gelu_for_Gelu_for_and_7_nl = (Gelu_for_8_else_else_acc_itm_28_1[27]) & (~
      Gelu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & (~ Gelu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_34_nl = act_regs_data_0_4_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_67_0;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_70_nl = MUX1HOT_s_1_3_2(Gelu_for_Gelu_for_and_7_nl,
      ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_2_31, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_34_nl,
      {and_dcpl_1007 , and_dcpl_832 , and_dcpl_852});
  assign ActUnit_PushOutput_if_output_port_reg_data_data_and_60_nl = (~ Gelu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & and_dcpl_1007;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_and_61_nl = Gelu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & and_dcpl_1007;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_85_nl = MUX1HOT_v_31_4_2(({{3{Gelu_for_8_else_else_acc_itm_28_1[27]}},
      Gelu_for_8_else_else_acc_itm_28_1}), nv_scvector_cctor_nv_scvector_6_for_8_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0,
      ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_2_30_0, act_regs_data_0_4_sva_dfm_2_30_0,
      {ActUnit_PushOutput_if_output_port_reg_data_data_and_60_nl , ActUnit_PushOutput_if_output_port_reg_data_data_and_61_nl
      , and_dcpl_832 , and_dcpl_852});
  assign nor_784_nl = ~(or_dcpl_655 | (and_dcpl_1007 & Gelu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs));
  assign Gelu_for_Gelu_for_and_8_nl = (z_out_28_1[27]) & (~ Gelu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & (~ Gelu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_41_nl = act_regs_data_0_5_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_exs_67_0;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_75_nl = MUX1HOT_s_1_3_2(Gelu_for_Gelu_for_and_8_nl,
      ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_2_31, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_41_nl,
      {and_dcpl_1007 , and_dcpl_832 , and_dcpl_852});
  assign ActUnit_PushOutput_if_output_port_reg_data_data_and_62_nl = (~ Gelu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & and_dcpl_1007;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_and_63_nl = Gelu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & and_dcpl_1007;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_84_nl = MUX1HOT_v_31_4_2(({{3{z_out_28_1[27]}},
      z_out_28_1}), nv_scvector_cctor_nv_scvector_6_for_9_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0,
      ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_2_30_0, act_regs_data_0_5_sva_dfm_2_30_0,
      {ActUnit_PushOutput_if_output_port_reg_data_data_and_62_nl , ActUnit_PushOutput_if_output_port_reg_data_data_and_63_nl
      , and_dcpl_832 , and_dcpl_852});
  assign nor_785_nl = ~(or_dcpl_655 | (and_dcpl_1007 & Gelu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_3_slc_operator_32_8_true_AC_TRN_AC_WRAP_3_acc_8_svs));
  assign while_while_mux1h_84_nl = MUX1HOT_s_1_6_2(act_regs_data_0_0_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[31]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_1_exs_5_30_0[30]), ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_31,
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_31, {while_asn_1383
      , while_asn_1385 , while_asn_1387 , while_asn_1389 , while_asn_1393 , while_asn_1395});
  assign while_and_273_nl = while_while_mux1h_84_nl & (~ while_asn_1391);
  assign while_while_mux1h_85_nl = MUX1HOT_s_1_6_2(act_regs_data_0_1_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[63]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_2_exs_5_30_0[30]), Silu_for_y_2_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_31,
      {while_asn_1383 , while_asn_1385 , while_asn_1387 , while_asn_1389 , while_asn_1393
      , while_asn_1395});
  assign while_and_272_nl = while_while_mux1h_85_nl & (~ while_asn_1391);
  assign while_while_mux1h_86_nl = MUX1HOT_s_1_6_2(act_regs_data_0_2_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[95]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_3_exs_5_30_0[30]), Silu_for_y_3_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_31,
      {while_asn_1383 , while_asn_1385 , while_asn_1387 , while_asn_1389 , while_asn_1393
      , while_asn_1395});
  assign while_and_271_nl = while_while_mux1h_86_nl & (~ while_asn_1391);
  assign while_while_mux1h_87_nl = MUX1HOT_s_1_6_2(act_regs_data_0_3_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[127]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_4_exs_5_30_0[30]), Silu_for_y_4_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_31,
      {while_asn_1383 , while_asn_1385 , while_asn_1387 , while_asn_1389 , while_asn_1393
      , while_asn_1395});
  assign while_and_270_nl = while_while_mux1h_87_nl & (~ while_asn_1391);
  assign while_while_mux1h_88_nl = MUX1HOT_s_1_6_2(act_regs_data_0_4_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[159]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_5_exs_5_30_0[30]), Silu_for_y_5_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_31,
      {while_asn_1383 , while_asn_1385 , while_asn_1387 , while_asn_1389 , while_asn_1393
      , while_asn_1395});
  assign while_and_269_nl = while_while_mux1h_88_nl & (~ while_asn_1391);
  assign while_while_mux1h_89_nl = MUX1HOT_s_1_6_2(act_regs_data_0_5_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[191]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_6_exs_5_30_0[30]), Silu_for_y_6_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_31,
      {while_asn_1383 , while_asn_1385 , while_asn_1387 , while_asn_1389 , while_asn_1393
      , while_asn_1395});
  assign while_and_268_nl = while_while_mux1h_89_nl & (~ while_asn_1391);
  assign while_while_mux1h_90_nl = MUX1HOT_s_1_6_2(act_regs_data_0_6_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[223]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_7_exs_5_30_0[30]), Silu_for_y_7_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_31,
      {while_asn_1383 , while_asn_1385 , while_asn_1387 , while_asn_1389 , while_asn_1393
      , while_asn_1395});
  assign while_and_267_nl = while_while_mux1h_90_nl & (~ while_asn_1391);
  assign while_while_mux1h_91_nl = MUX1HOT_s_1_6_2(act_regs_data_0_7_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[255]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_8_exs_5_30_0[30]), Silu_for_y_8_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_31,
      {while_asn_1383 , while_asn_1385 , while_asn_1387 , while_asn_1389 , while_asn_1393
      , while_asn_1395});
  assign while_and_266_nl = while_while_mux1h_91_nl & (~ while_asn_1391);
  assign while_while_mux1h_92_nl = MUX1HOT_s_1_6_2(act_regs_data_0_8_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[287]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_9_exs_5_30_0[30]), Silu_for_y_9_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_31,
      {while_asn_1383 , while_asn_1385 , while_asn_1387 , while_asn_1389 , while_asn_1393
      , while_asn_1395});
  assign while_and_265_nl = while_while_mux1h_92_nl & (~ while_asn_1391);
  assign while_while_mux1h_93_nl = MUX1HOT_s_1_6_2(act_regs_data_0_9_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[319]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_10_exs_5_30_0[30]), ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_31,
      Gelu_for_y_10_lpi_1_dfm_2_31, {while_asn_1383 , while_asn_1385 , while_asn_1387
      , while_asn_1389 , while_asn_1393 , while_asn_1395});
  assign while_and_264_nl = while_while_mux1h_93_nl & (~ while_asn_1391);
  assign while_while_mux1h_94_nl = MUX1HOT_s_1_6_2(act_regs_data_0_10_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[351]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_11_exs_5_30_0[30]), ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_31,
      Gelu_for_y_11_lpi_1_dfm_2_31, {while_asn_1383 , while_asn_1385 , while_asn_1387
      , while_asn_1389 , while_asn_1393 , while_asn_1395});
  assign while_and_263_nl = while_while_mux1h_94_nl & (~ while_asn_1391);
  assign while_while_mux1h_95_nl = MUX1HOT_s_1_6_2(act_regs_data_0_11_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[383]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_12_exs_5_30_0[30]), Silu_for_y_12_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_31,
      {while_asn_1383 , while_asn_1385 , while_asn_1387 , while_asn_1389 , while_asn_1393
      , while_asn_1395});
  assign while_and_262_nl = while_while_mux1h_95_nl & (~ while_asn_1391);
  assign while_while_mux1h_96_nl = MUX1HOT_s_1_6_2(act_regs_data_0_12_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[415]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_13_exs_5_30_0[30]), Silu_for_y_13_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_1_sva_31,
      {while_asn_1383 , while_asn_1385 , while_asn_1387 , while_asn_1389 , while_asn_1393
      , while_asn_1395});
  assign while_and_261_nl = while_while_mux1h_96_nl & (~ while_asn_1391);
  assign while_while_mux1h_97_nl = MUX1HOT_s_1_6_2(act_regs_data_0_13_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[447]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_14_exs_5_30_0[30]), Silu_for_y_14_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_31,
      {while_asn_1383 , while_asn_1385 , while_asn_1387 , while_asn_1389 , while_asn_1393
      , while_asn_1395});
  assign while_and_260_nl = while_while_mux1h_97_nl & (~ while_asn_1391);
  assign while_while_mux1h_98_nl = MUX1HOT_s_1_6_2(act_regs_data_0_14_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[479]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_15_exs_5_30_0[30]), Silu_for_y_15_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_31,
      {while_asn_1383 , while_asn_1385 , while_asn_1387 , while_asn_1389 , while_asn_1393
      , while_asn_1395});
  assign while_and_259_nl = while_while_mux1h_98_nl & (~ while_asn_1391);
  assign while_while_mux1h_99_nl = MUX1HOT_s_1_6_2(act_regs_data_0_15_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[511]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_16_exs_5_30_0[30]), Silu_for_y_lpi_1_dfm_1_31, Gelu_for_y_lpi_1_dfm_2_31,
      {while_asn_1383 , while_asn_1385 , while_asn_1387 , while_asn_1389 , while_asn_1393
      , while_asn_1395});
  assign while_and_258_nl = while_while_mux1h_99_nl & (~ while_asn_1391);
  assign while_while_mux1h_100_nl = MUX1HOT_s_1_6_2(act_regs_data_1_0_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[31]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_1_exs_5_30_0[30]), ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_31,
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_31, {while_asn_1369
      , while_asn_1371 , while_asn_1373 , while_asn_1375 , while_asn_1379 , while_asn_1381});
  assign while_and_257_nl = while_while_mux1h_100_nl & (~ while_asn_1377);
  assign while_while_mux1h_101_nl = MUX1HOT_s_1_6_2(act_regs_data_1_1_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[63]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_2_exs_5_30_0[30]), Silu_for_y_2_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_31,
      {while_asn_1369 , while_asn_1371 , while_asn_1373 , while_asn_1375 , while_asn_1379
      , while_asn_1381});
  assign while_and_256_nl = while_while_mux1h_101_nl & (~ while_asn_1377);
  assign while_while_mux1h_102_nl = MUX1HOT_s_1_6_2(act_regs_data_1_2_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[95]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_3_exs_5_30_0[30]), Silu_for_y_3_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_31,
      {while_asn_1369 , while_asn_1371 , while_asn_1373 , while_asn_1375 , while_asn_1379
      , while_asn_1381});
  assign while_and_255_nl = while_while_mux1h_102_nl & (~ while_asn_1377);
  assign while_while_mux1h_103_nl = MUX1HOT_s_1_6_2(act_regs_data_1_3_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[127]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_4_exs_5_30_0[30]), Silu_for_y_4_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_31,
      {while_asn_1369 , while_asn_1371 , while_asn_1373 , while_asn_1375 , while_asn_1379
      , while_asn_1381});
  assign while_and_254_nl = while_while_mux1h_103_nl & (~ while_asn_1377);
  assign while_while_mux1h_104_nl = MUX1HOT_s_1_6_2(act_regs_data_1_4_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[159]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_5_exs_5_30_0[30]), Silu_for_y_5_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_31,
      {while_asn_1369 , while_asn_1371 , while_asn_1373 , while_asn_1375 , while_asn_1379
      , while_asn_1381});
  assign while_and_253_nl = while_while_mux1h_104_nl & (~ while_asn_1377);
  assign while_while_mux1h_105_nl = MUX1HOT_s_1_6_2(act_regs_data_1_5_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[191]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_6_exs_5_30_0[30]), Silu_for_y_6_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_31,
      {while_asn_1369 , while_asn_1371 , while_asn_1373 , while_asn_1375 , while_asn_1379
      , while_asn_1381});
  assign while_and_252_nl = while_while_mux1h_105_nl & (~ while_asn_1377);
  assign while_while_mux1h_106_nl = MUX1HOT_s_1_6_2(act_regs_data_1_6_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[223]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_7_exs_5_30_0[30]), Silu_for_y_7_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_31,
      {while_asn_1369 , while_asn_1371 , while_asn_1373 , while_asn_1375 , while_asn_1379
      , while_asn_1381});
  assign while_and_251_nl = while_while_mux1h_106_nl & (~ while_asn_1377);
  assign while_while_mux1h_107_nl = MUX1HOT_s_1_6_2(act_regs_data_1_7_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[255]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_8_exs_5_30_0[30]), Silu_for_y_8_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_31,
      {while_asn_1369 , while_asn_1371 , while_asn_1373 , while_asn_1375 , while_asn_1379
      , while_asn_1381});
  assign while_and_250_nl = while_while_mux1h_107_nl & (~ while_asn_1377);
  assign while_while_mux1h_108_nl = MUX1HOT_s_1_6_2(act_regs_data_1_8_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[287]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_9_exs_5_30_0[30]), Silu_for_y_9_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_31,
      {while_asn_1369 , while_asn_1371 , while_asn_1373 , while_asn_1375 , while_asn_1379
      , while_asn_1381});
  assign while_and_249_nl = while_while_mux1h_108_nl & (~ while_asn_1377);
  assign while_while_mux1h_109_nl = MUX1HOT_s_1_6_2(act_regs_data_1_9_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[319]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_10_exs_5_30_0[30]), ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_31,
      Gelu_for_y_10_lpi_1_dfm_2_31, {while_asn_1369 , while_asn_1371 , while_asn_1373
      , while_asn_1375 , while_asn_1379 , while_asn_1381});
  assign while_and_248_nl = while_while_mux1h_109_nl & (~ while_asn_1377);
  assign while_while_mux1h_110_nl = MUX1HOT_s_1_6_2(act_regs_data_1_10_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[351]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_11_exs_5_30_0[30]), ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_31,
      Gelu_for_y_11_lpi_1_dfm_2_31, {while_asn_1369 , while_asn_1371 , while_asn_1373
      , while_asn_1375 , while_asn_1379 , while_asn_1381});
  assign while_and_247_nl = while_while_mux1h_110_nl & (~ while_asn_1377);
  assign while_while_mux1h_111_nl = MUX1HOT_s_1_6_2(act_regs_data_1_11_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[383]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_12_exs_5_30_0[30]), Silu_for_y_12_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_31,
      {while_asn_1369 , while_asn_1371 , while_asn_1373 , while_asn_1375 , while_asn_1379
      , while_asn_1381});
  assign while_and_246_nl = while_while_mux1h_111_nl & (~ while_asn_1377);
  assign while_while_mux1h_112_nl = MUX1HOT_s_1_6_2(act_regs_data_1_12_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[415]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_13_exs_5_30_0[30]), Silu_for_y_13_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_1_sva_31,
      {while_asn_1369 , while_asn_1371 , while_asn_1373 , while_asn_1375 , while_asn_1379
      , while_asn_1381});
  assign while_and_245_nl = while_while_mux1h_112_nl & (~ while_asn_1377);
  assign while_while_mux1h_113_nl = MUX1HOT_s_1_6_2(act_regs_data_1_13_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[447]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_14_exs_5_30_0[30]), Silu_for_y_14_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_31,
      {while_asn_1369 , while_asn_1371 , while_asn_1373 , while_asn_1375 , while_asn_1379
      , while_asn_1381});
  assign while_and_244_nl = while_while_mux1h_113_nl & (~ while_asn_1377);
  assign while_while_mux1h_114_nl = MUX1HOT_s_1_6_2(act_regs_data_1_14_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[479]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_15_exs_5_30_0[30]), Silu_for_y_15_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_31,
      {while_asn_1369 , while_asn_1371 , while_asn_1373 , while_asn_1375 , while_asn_1379
      , while_asn_1381});
  assign while_and_243_nl = while_while_mux1h_114_nl & (~ while_asn_1377);
  assign while_while_mux1h_115_nl = MUX1HOT_s_1_6_2(act_regs_data_1_15_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[511]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_16_exs_5_30_0[30]), Silu_for_y_lpi_1_dfm_1_31, Gelu_for_y_lpi_1_dfm_2_31,
      {while_asn_1369 , while_asn_1371 , while_asn_1373 , while_asn_1375 , while_asn_1379
      , while_asn_1381});
  assign while_and_242_nl = while_while_mux1h_115_nl & (~ while_asn_1377);
  assign while_while_mux1h_116_nl = MUX1HOT_s_1_6_2(act_regs_data_2_0_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[31]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_1_exs_5_30_0[30]), ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_31,
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_31, {while_asn_1355
      , while_asn_1357 , while_asn_1359 , while_asn_1361 , while_asn_1365 , while_asn_1367});
  assign while_and_241_nl = while_while_mux1h_116_nl & (~ while_asn_1363);
  assign while_while_mux1h_117_nl = MUX1HOT_s_1_6_2(act_regs_data_2_1_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[63]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_2_exs_5_30_0[30]), Silu_for_y_2_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_31,
      {while_asn_1355 , while_asn_1357 , while_asn_1359 , while_asn_1361 , while_asn_1365
      , while_asn_1367});
  assign while_and_240_nl = while_while_mux1h_117_nl & (~ while_asn_1363);
  assign while_while_mux1h_118_nl = MUX1HOT_s_1_6_2(act_regs_data_2_2_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[95]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_3_exs_5_30_0[30]), Silu_for_y_3_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_31,
      {while_asn_1355 , while_asn_1357 , while_asn_1359 , while_asn_1361 , while_asn_1365
      , while_asn_1367});
  assign while_and_239_nl = while_while_mux1h_118_nl & (~ while_asn_1363);
  assign while_while_mux1h_119_nl = MUX1HOT_s_1_6_2(act_regs_data_2_3_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[127]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_4_exs_5_30_0[30]), Silu_for_y_4_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_31,
      {while_asn_1355 , while_asn_1357 , while_asn_1359 , while_asn_1361 , while_asn_1365
      , while_asn_1367});
  assign while_and_238_nl = while_while_mux1h_119_nl & (~ while_asn_1363);
  assign while_while_mux1h_120_nl = MUX1HOT_s_1_6_2(act_regs_data_2_4_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[159]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_5_exs_5_30_0[30]), Silu_for_y_5_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_31,
      {while_asn_1355 , while_asn_1357 , while_asn_1359 , while_asn_1361 , while_asn_1365
      , while_asn_1367});
  assign while_and_237_nl = while_while_mux1h_120_nl & (~ while_asn_1363);
  assign while_while_mux1h_121_nl = MUX1HOT_s_1_6_2(act_regs_data_2_5_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[191]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_6_exs_5_30_0[30]), Silu_for_y_6_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_31,
      {while_asn_1355 , while_asn_1357 , while_asn_1359 , while_asn_1361 , while_asn_1365
      , while_asn_1367});
  assign while_and_236_nl = while_while_mux1h_121_nl & (~ while_asn_1363);
  assign while_while_mux1h_122_nl = MUX1HOT_s_1_6_2(act_regs_data_2_6_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[223]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_7_exs_5_30_0[30]), Silu_for_y_7_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_31,
      {while_asn_1355 , while_asn_1357 , while_asn_1359 , while_asn_1361 , while_asn_1365
      , while_asn_1367});
  assign while_and_235_nl = while_while_mux1h_122_nl & (~ while_asn_1363);
  assign while_while_mux1h_123_nl = MUX1HOT_s_1_6_2(act_regs_data_2_7_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[255]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_8_exs_5_30_0[30]), Silu_for_y_8_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_31,
      {while_asn_1355 , while_asn_1357 , while_asn_1359 , while_asn_1361 , while_asn_1365
      , while_asn_1367});
  assign while_and_234_nl = while_while_mux1h_123_nl & (~ while_asn_1363);
  assign while_while_mux1h_124_nl = MUX1HOT_s_1_6_2(act_regs_data_2_8_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[287]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_9_exs_5_30_0[30]), Silu_for_y_9_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_31,
      {while_asn_1355 , while_asn_1357 , while_asn_1359 , while_asn_1361 , while_asn_1365
      , while_asn_1367});
  assign while_and_233_nl = while_while_mux1h_124_nl & (~ while_asn_1363);
  assign while_while_mux1h_125_nl = MUX1HOT_s_1_6_2(act_regs_data_2_9_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[319]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_10_exs_5_30_0[30]), ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_31,
      Gelu_for_y_10_lpi_1_dfm_2_31, {while_asn_1355 , while_asn_1357 , while_asn_1359
      , while_asn_1361 , while_asn_1365 , while_asn_1367});
  assign while_and_232_nl = while_while_mux1h_125_nl & (~ while_asn_1363);
  assign while_while_mux1h_126_nl = MUX1HOT_s_1_6_2(act_regs_data_2_10_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[351]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_11_exs_5_30_0[30]), ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_31,
      Gelu_for_y_11_lpi_1_dfm_2_31, {while_asn_1355 , while_asn_1357 , while_asn_1359
      , while_asn_1361 , while_asn_1365 , while_asn_1367});
  assign while_and_231_nl = while_while_mux1h_126_nl & (~ while_asn_1363);
  assign while_while_mux1h_127_nl = MUX1HOT_s_1_6_2(act_regs_data_2_11_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[383]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_12_exs_5_30_0[30]), Silu_for_y_12_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_31,
      {while_asn_1355 , while_asn_1357 , while_asn_1359 , while_asn_1361 , while_asn_1365
      , while_asn_1367});
  assign while_and_230_nl = while_while_mux1h_127_nl & (~ while_asn_1363);
  assign while_while_mux1h_128_nl = MUX1HOT_s_1_6_2(act_regs_data_2_12_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[415]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_13_exs_5_30_0[30]), Silu_for_y_13_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_1_sva_31,
      {while_asn_1355 , while_asn_1357 , while_asn_1359 , while_asn_1361 , while_asn_1365
      , while_asn_1367});
  assign while_and_229_nl = while_while_mux1h_128_nl & (~ while_asn_1363);
  assign while_while_mux1h_129_nl = MUX1HOT_s_1_6_2(act_regs_data_2_13_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[447]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_14_exs_5_30_0[30]), Silu_for_y_14_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_31,
      {while_asn_1355 , while_asn_1357 , while_asn_1359 , while_asn_1361 , while_asn_1365
      , while_asn_1367});
  assign while_and_228_nl = while_while_mux1h_129_nl & (~ while_asn_1363);
  assign while_while_mux1h_130_nl = MUX1HOT_s_1_6_2(act_regs_data_2_14_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[479]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_15_exs_5_30_0[30]), Silu_for_y_15_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_31,
      {while_asn_1355 , while_asn_1357 , while_asn_1359 , while_asn_1361 , while_asn_1365
      , while_asn_1367});
  assign while_and_227_nl = while_while_mux1h_130_nl & (~ while_asn_1363);
  assign while_while_mux1h_131_nl = MUX1HOT_s_1_6_2(act_regs_data_2_15_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[511]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_16_exs_5_30_0[30]), Silu_for_y_lpi_1_dfm_1_31, Gelu_for_y_lpi_1_dfm_2_31,
      {while_asn_1355 , while_asn_1357 , while_asn_1359 , while_asn_1361 , while_asn_1365
      , while_asn_1367});
  assign while_and_226_nl = while_while_mux1h_131_nl & (~ while_asn_1363);
  assign while_while_mux1h_132_nl = MUX1HOT_s_1_6_2(act_regs_data_3_0_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[31]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_1_exs_5_30_0[30]), ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_31,
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_31, {while_asn_1341
      , while_asn_1343 , while_asn_1345 , while_asn_1347 , while_asn_1351 , while_asn_1353});
  assign while_and_225_nl = while_while_mux1h_132_nl & (~ while_asn_1349);
  assign while_while_mux1h_133_nl = MUX1HOT_s_1_6_2(act_regs_data_3_1_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[63]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_2_exs_5_30_0[30]), Silu_for_y_2_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_31,
      {while_asn_1341 , while_asn_1343 , while_asn_1345 , while_asn_1347 , while_asn_1351
      , while_asn_1353});
  assign while_and_224_nl = while_while_mux1h_133_nl & (~ while_asn_1349);
  assign while_while_mux1h_134_nl = MUX1HOT_s_1_6_2(act_regs_data_3_2_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[95]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_3_exs_5_30_0[30]), Silu_for_y_3_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_31,
      {while_asn_1341 , while_asn_1343 , while_asn_1345 , while_asn_1347 , while_asn_1351
      , while_asn_1353});
  assign while_and_223_nl = while_while_mux1h_134_nl & (~ while_asn_1349);
  assign while_while_mux1h_135_nl = MUX1HOT_s_1_6_2(act_regs_data_3_3_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[127]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_4_exs_5_30_0[30]), Silu_for_y_4_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_31,
      {while_asn_1341 , while_asn_1343 , while_asn_1345 , while_asn_1347 , while_asn_1351
      , while_asn_1353});
  assign while_and_222_nl = while_while_mux1h_135_nl & (~ while_asn_1349);
  assign while_while_mux1h_136_nl = MUX1HOT_s_1_6_2(act_regs_data_3_4_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[159]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_5_exs_5_30_0[30]), Silu_for_y_5_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_31,
      {while_asn_1341 , while_asn_1343 , while_asn_1345 , while_asn_1347 , while_asn_1351
      , while_asn_1353});
  assign while_and_221_nl = while_while_mux1h_136_nl & (~ while_asn_1349);
  assign while_while_mux1h_137_nl = MUX1HOT_s_1_6_2(act_regs_data_3_5_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[191]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_6_exs_5_30_0[30]), Silu_for_y_6_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_31,
      {while_asn_1341 , while_asn_1343 , while_asn_1345 , while_asn_1347 , while_asn_1351
      , while_asn_1353});
  assign while_and_220_nl = while_while_mux1h_137_nl & (~ while_asn_1349);
  assign while_while_mux1h_138_nl = MUX1HOT_s_1_6_2(act_regs_data_3_6_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[223]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_7_exs_5_30_0[30]), Silu_for_y_7_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_31,
      {while_asn_1341 , while_asn_1343 , while_asn_1345 , while_asn_1347 , while_asn_1351
      , while_asn_1353});
  assign while_and_219_nl = while_while_mux1h_138_nl & (~ while_asn_1349);
  assign while_while_mux1h_139_nl = MUX1HOT_s_1_6_2(act_regs_data_3_7_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[255]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_8_exs_5_30_0[30]), Silu_for_y_8_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_31,
      {while_asn_1341 , while_asn_1343 , while_asn_1345 , while_asn_1347 , while_asn_1351
      , while_asn_1353});
  assign while_and_218_nl = while_while_mux1h_139_nl & (~ while_asn_1349);
  assign while_while_mux1h_140_nl = MUX1HOT_s_1_6_2(act_regs_data_3_8_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[287]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_9_exs_5_30_0[30]), Silu_for_y_9_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_31,
      {while_asn_1341 , while_asn_1343 , while_asn_1345 , while_asn_1347 , while_asn_1351
      , while_asn_1353});
  assign while_and_217_nl = while_while_mux1h_140_nl & (~ while_asn_1349);
  assign while_while_mux1h_141_nl = MUX1HOT_s_1_6_2(act_regs_data_3_9_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[319]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_10_exs_5_30_0[30]), ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_31,
      Gelu_for_y_10_lpi_1_dfm_2_31, {while_asn_1341 , while_asn_1343 , while_asn_1345
      , while_asn_1347 , while_asn_1351 , while_asn_1353});
  assign while_and_216_nl = while_while_mux1h_141_nl & (~ while_asn_1349);
  assign while_while_mux1h_142_nl = MUX1HOT_s_1_6_2(act_regs_data_3_10_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[351]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_11_exs_5_30_0[30]), ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_31,
      Gelu_for_y_11_lpi_1_dfm_2_31, {while_asn_1341 , while_asn_1343 , while_asn_1345
      , while_asn_1347 , while_asn_1351 , while_asn_1353});
  assign while_and_215_nl = while_while_mux1h_142_nl & (~ while_asn_1349);
  assign while_while_mux1h_143_nl = MUX1HOT_s_1_6_2(act_regs_data_3_11_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[383]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_12_exs_5_30_0[30]), Silu_for_y_12_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_31,
      {while_asn_1341 , while_asn_1343 , while_asn_1345 , while_asn_1347 , while_asn_1351
      , while_asn_1353});
  assign while_and_214_nl = while_while_mux1h_143_nl & (~ while_asn_1349);
  assign while_while_mux1h_144_nl = MUX1HOT_s_1_6_2(act_regs_data_3_12_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[415]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_13_exs_5_30_0[30]), Silu_for_y_13_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_1_sva_31,
      {while_asn_1341 , while_asn_1343 , while_asn_1345 , while_asn_1347 , while_asn_1351
      , while_asn_1353});
  assign while_and_213_nl = while_while_mux1h_144_nl & (~ while_asn_1349);
  assign while_while_mux1h_145_nl = MUX1HOT_s_1_6_2(act_regs_data_3_13_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[447]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_14_exs_5_30_0[30]), Silu_for_y_14_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_31,
      {while_asn_1341 , while_asn_1343 , while_asn_1345 , while_asn_1347 , while_asn_1351
      , while_asn_1353});
  assign while_and_212_nl = while_while_mux1h_145_nl & (~ while_asn_1349);
  assign while_while_mux1h_146_nl = MUX1HOT_s_1_6_2(act_regs_data_3_14_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[479]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_15_exs_5_30_0[30]), Silu_for_y_15_lpi_1_dfm_1_31, ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_31,
      {while_asn_1341 , while_asn_1343 , while_asn_1345 , while_asn_1347 , while_asn_1351
      , while_asn_1353});
  assign while_and_211_nl = while_while_mux1h_146_nl & (~ while_asn_1349);
  assign while_while_mux1h_147_nl = MUX1HOT_s_1_6_2(act_regs_data_3_15_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[511]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      (Tanh_for_16_exs_5_30_0[30]), Silu_for_y_lpi_1_dfm_1_31, Gelu_for_y_lpi_1_dfm_2_31,
      {while_asn_1341 , while_asn_1343 , while_asn_1345 , while_asn_1347 , while_asn_1351
      , while_asn_1353});
  assign while_and_nl = while_while_mux1h_147_nl & (~ while_asn_1349);
  assign or_399_nl = (~ act_config_InstIncr_if_equal_1_tmp) | (operator_6_false_acc_tmp[6:5]!=2'b00);
  assign mux_82_nl = MUX_s_1_2_2(is_start_sva, (~ is_start_sva), or_399_nl);
  assign act_config_InstIncr_if_act_config_InstIncr_if_and_nl = act_config_is_zero_first_sva_dfm_4
      & (~ act_config_InstIncr_if_act_config_InstIncr_if_if_nor_tmp);
  assign act_config_InstIncr_mux_2_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_config_InstIncr_if_act_config_InstIncr_if_and_nl, act_config_InstIncr_act_config_InstIncr_if_and_svs_1);
  assign nor_768_nl = ~((~ (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[0])) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[8]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[9]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[10]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])));
  assign or_1509_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[0]) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[8]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[9]) | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11]))
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[10]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]));
  assign mux_578_nl = MUX_s_1_2_2(nor_768_nl, or_1509_nl, act_config_is_valid_sva);
  assign and_1143_nl = and_dcpl_1001 & (fsm_output[2:0]==3'b011);
  assign and_1146_nl = and_dcpl_1013 & and_dcpl_563;
  assign and_1148_nl = and_dcpl_1013 & (fsm_output[1:0]==2'b01);
  assign Gelu_for_else_else_mux1h_10_nl = MUX1HOT_v_26_3_2((nv_scvector_cctor_nv_scvector_6_for_12_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_6_for_9_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_6_for_16_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      {and_1143_nl , and_1146_nl , and_1148_nl});
  assign nl_Gelu_for_12_else_else_acc_rg_1_nl = conv_s2u_28_29(Tanh_for_1_else_else_mul_cmp_13_z[72:45])
      + conv_s2u_26_29(Gelu_for_else_else_mux1h_10_nl);
  assign Gelu_for_12_else_else_acc_rg_1_nl = nl_Gelu_for_12_else_else_acc_rg_1_nl[28:0];
  assign z_out_28_1 = readslicef_29_28_1(Gelu_for_12_else_else_acc_rg_1_nl);
  assign and_1162_nl = and_dcpl_1028 & and_dcpl_1021;
  assign Gelu_for_else_else_mux1h_12_nl = MUX1HOT_v_26_6_2((nv_scvector_cctor_nv_scvector_6_for_2_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_6_for_3_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_6_for_4_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_6_for_6_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_6_for_15_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_6_for_10_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      {and_1152_cse , and_1154_cse , and_1156_cse , and_1158_cse , and_1161_cse ,
      and_1162_nl});
  assign nl_Gelu_for_10_else_else_acc_rg_1_nl = conv_s2u_28_29(Tanh_for_1_else_else_mul_cmp_12_z[72:45])
      + conv_s2u_26_29(Gelu_for_else_else_mux1h_12_nl);
  assign Gelu_for_10_else_else_acc_rg_1_nl = nl_Gelu_for_10_else_else_acc_rg_1_nl[28:0];
  assign z_out_1_28_1 = readslicef_29_28_1(Gelu_for_10_else_else_acc_rg_1_nl);
  assign and_1175_nl = and_dcpl_1028 & (fsm_output[1:0]==2'b01);
  assign Gelu_for_else_else_mux1h_14_nl = MUX1HOT_v_26_5_2((ActUnit_RunInst_case_15_nv_scvector_cctor_data_0_sva_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_6_for_5_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_6_for_7_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_6_for_14_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      (nv_scvector_cctor_nv_scvector_6_for_11_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[25:0]),
      {and_1152_cse , and_1156_cse , and_1158_cse , and_1161_cse , and_1175_nl});
  assign nl_Gelu_for_11_else_else_acc_rg_1_nl = conv_s2u_28_29(Tanh_for_1_else_else_mul_cmp_z[72:45])
      + conv_s2u_26_29(Gelu_for_else_else_mux1h_14_nl);
  assign Gelu_for_11_else_else_acc_rg_1_nl = nl_Gelu_for_11_else_else_acc_rg_1_nl[28:0];
  assign z_out_2_28_1 = readslicef_29_28_1(Gelu_for_11_else_else_acc_rg_1_nl);
  assign and_1179_nl = and_dcpl_1046 & and_dcpl_563;
  assign Silu_for_else_else_mux1h_1_nl = MUX1HOT_v_27_8_2((nv_scvector_cctor_nv_scvector_5_for_2_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[26:0]),
      (nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[26:0]),
      (nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[26:0]),
      (nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[26:0]),
      (nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[26:0]),
      (nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[26:0]),
      (nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[26:0]),
      (nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[26:0]),
      {and_1179_nl , and_1181_cse , and_1183_cse , and_1185_cse , and_1152_cse ,
      and_1154_cse , and_1190_cse , and_1191_cse});
  assign nl_Silu_for_10_else_else_acc_rg_1_nl = conv_s2u_29_30(Tanh_for_1_else_else_mul_1_cmp_1_z[53:25])
      + conv_s2u_27_30(Silu_for_else_else_mux1h_1_nl);
  assign Silu_for_10_else_else_acc_rg_1_nl = nl_Silu_for_10_else_else_acc_rg_1_nl[29:0];
  assign z_out_3_29_1 = readslicef_30_29_1(Silu_for_10_else_else_acc_rg_1_nl);
  assign Silu_for_else_else_mux1h_3_nl = MUX1HOT_v_27_7_2((nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[26:0]),
      (nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[26:0]),
      (nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[26:0]),
      (nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[26:0]),
      (nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[26:0]),
      (nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[26:0]),
      (nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_0[26:0]),
      {and_1181_cse , and_1183_cse , and_1185_cse , and_1152_cse , and_1154_cse ,
      and_1190_cse , and_1191_cse});
  assign nl_Silu_for_11_else_else_acc_rg_1_nl = conv_s2u_29_30(Tanh_for_1_else_else_mul_1_cmp_z[53:25])
      + conv_s2u_27_30(Silu_for_else_else_mux1h_3_nl);
  assign Silu_for_11_else_else_acc_rg_1_nl = nl_Silu_for_11_else_else_acc_rg_1_nl[29:0];
  assign z_out_4_29_1 = readslicef_30_29_1(Silu_for_11_else_else_acc_rg_1_nl);

  function automatic  MUX1HOT_s_1_14_2;
    input  input_13;
    input  input_12;
    input  input_11;
    input  input_10;
    input  input_9;
    input  input_8;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [13:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    result = result | (input_9 & sel[9]);
    result = result | (input_10 & sel[10]);
    result = result | (input_11 & sel[11]);
    result = result | (input_12 & sel[12]);
    result = result | (input_13 & sel[13]);
    MUX1HOT_s_1_14_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_1_2;
    input  input_0;
    input  sel;
    reg  result;
  begin
    result = input_0 & sel;
    MUX1HOT_s_1_1_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_3_2;
    input  input_2;
    input  input_1;
    input  input_0;
    input [2:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_4_2;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [3:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_6_2;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [5:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    MUX1HOT_s_1_6_2 = result;
  end
  endfunction


  function automatic [25:0] MUX1HOT_v_26_13_2;
    input [25:0] input_12;
    input [25:0] input_11;
    input [25:0] input_10;
    input [25:0] input_9;
    input [25:0] input_8;
    input [25:0] input_7;
    input [25:0] input_6;
    input [25:0] input_5;
    input [25:0] input_4;
    input [25:0] input_3;
    input [25:0] input_2;
    input [25:0] input_1;
    input [25:0] input_0;
    input [12:0] sel;
    reg [25:0] result;
  begin
    result = input_0 & {26{sel[0]}};
    result = result | (input_1 & {26{sel[1]}});
    result = result | (input_2 & {26{sel[2]}});
    result = result | (input_3 & {26{sel[3]}});
    result = result | (input_4 & {26{sel[4]}});
    result = result | (input_5 & {26{sel[5]}});
    result = result | (input_6 & {26{sel[6]}});
    result = result | (input_7 & {26{sel[7]}});
    result = result | (input_8 & {26{sel[8]}});
    result = result | (input_9 & {26{sel[9]}});
    result = result | (input_10 & {26{sel[10]}});
    result = result | (input_11 & {26{sel[11]}});
    result = result | (input_12 & {26{sel[12]}});
    MUX1HOT_v_26_13_2 = result;
  end
  endfunction


  function automatic [25:0] MUX1HOT_v_26_3_2;
    input [25:0] input_2;
    input [25:0] input_1;
    input [25:0] input_0;
    input [2:0] sel;
    reg [25:0] result;
  begin
    result = input_0 & {26{sel[0]}};
    result = result | (input_1 & {26{sel[1]}});
    result = result | (input_2 & {26{sel[2]}});
    MUX1HOT_v_26_3_2 = result;
  end
  endfunction


  function automatic [25:0] MUX1HOT_v_26_5_2;
    input [25:0] input_4;
    input [25:0] input_3;
    input [25:0] input_2;
    input [25:0] input_1;
    input [25:0] input_0;
    input [4:0] sel;
    reg [25:0] result;
  begin
    result = input_0 & {26{sel[0]}};
    result = result | (input_1 & {26{sel[1]}});
    result = result | (input_2 & {26{sel[2]}});
    result = result | (input_3 & {26{sel[3]}});
    result = result | (input_4 & {26{sel[4]}});
    MUX1HOT_v_26_5_2 = result;
  end
  endfunction


  function automatic [25:0] MUX1HOT_v_26_6_2;
    input [25:0] input_5;
    input [25:0] input_4;
    input [25:0] input_3;
    input [25:0] input_2;
    input [25:0] input_1;
    input [25:0] input_0;
    input [5:0] sel;
    reg [25:0] result;
  begin
    result = input_0 & {26{sel[0]}};
    result = result | (input_1 & {26{sel[1]}});
    result = result | (input_2 & {26{sel[2]}});
    result = result | (input_3 & {26{sel[3]}});
    result = result | (input_4 & {26{sel[4]}});
    result = result | (input_5 & {26{sel[5]}});
    MUX1HOT_v_26_6_2 = result;
  end
  endfunction


  function automatic [25:0] MUX1HOT_v_26_7_2;
    input [25:0] input_6;
    input [25:0] input_5;
    input [25:0] input_4;
    input [25:0] input_3;
    input [25:0] input_2;
    input [25:0] input_1;
    input [25:0] input_0;
    input [6:0] sel;
    reg [25:0] result;
  begin
    result = input_0 & {26{sel[0]}};
    result = result | (input_1 & {26{sel[1]}});
    result = result | (input_2 & {26{sel[2]}});
    result = result | (input_3 & {26{sel[3]}});
    result = result | (input_4 & {26{sel[4]}});
    result = result | (input_5 & {26{sel[5]}});
    result = result | (input_6 & {26{sel[6]}});
    MUX1HOT_v_26_7_2 = result;
  end
  endfunction


  function automatic [25:0] MUX1HOT_v_26_8_2;
    input [25:0] input_7;
    input [25:0] input_6;
    input [25:0] input_5;
    input [25:0] input_4;
    input [25:0] input_3;
    input [25:0] input_2;
    input [25:0] input_1;
    input [25:0] input_0;
    input [7:0] sel;
    reg [25:0] result;
  begin
    result = input_0 & {26{sel[0]}};
    result = result | (input_1 & {26{sel[1]}});
    result = result | (input_2 & {26{sel[2]}});
    result = result | (input_3 & {26{sel[3]}});
    result = result | (input_4 & {26{sel[4]}});
    result = result | (input_5 & {26{sel[5]}});
    result = result | (input_6 & {26{sel[6]}});
    result = result | (input_7 & {26{sel[7]}});
    MUX1HOT_v_26_8_2 = result;
  end
  endfunction


  function automatic [26:0] MUX1HOT_v_27_10_2;
    input [26:0] input_9;
    input [26:0] input_8;
    input [26:0] input_7;
    input [26:0] input_6;
    input [26:0] input_5;
    input [26:0] input_4;
    input [26:0] input_3;
    input [26:0] input_2;
    input [26:0] input_1;
    input [26:0] input_0;
    input [9:0] sel;
    reg [26:0] result;
  begin
    result = input_0 & {27{sel[0]}};
    result = result | (input_1 & {27{sel[1]}});
    result = result | (input_2 & {27{sel[2]}});
    result = result | (input_3 & {27{sel[3]}});
    result = result | (input_4 & {27{sel[4]}});
    result = result | (input_5 & {27{sel[5]}});
    result = result | (input_6 & {27{sel[6]}});
    result = result | (input_7 & {27{sel[7]}});
    result = result | (input_8 & {27{sel[8]}});
    result = result | (input_9 & {27{sel[9]}});
    MUX1HOT_v_27_10_2 = result;
  end
  endfunction


  function automatic [26:0] MUX1HOT_v_27_7_2;
    input [26:0] input_6;
    input [26:0] input_5;
    input [26:0] input_4;
    input [26:0] input_3;
    input [26:0] input_2;
    input [26:0] input_1;
    input [26:0] input_0;
    input [6:0] sel;
    reg [26:0] result;
  begin
    result = input_0 & {27{sel[0]}};
    result = result | (input_1 & {27{sel[1]}});
    result = result | (input_2 & {27{sel[2]}});
    result = result | (input_3 & {27{sel[3]}});
    result = result | (input_4 & {27{sel[4]}});
    result = result | (input_5 & {27{sel[5]}});
    result = result | (input_6 & {27{sel[6]}});
    MUX1HOT_v_27_7_2 = result;
  end
  endfunction


  function automatic [26:0] MUX1HOT_v_27_8_2;
    input [26:0] input_7;
    input [26:0] input_6;
    input [26:0] input_5;
    input [26:0] input_4;
    input [26:0] input_3;
    input [26:0] input_2;
    input [26:0] input_1;
    input [26:0] input_0;
    input [7:0] sel;
    reg [26:0] result;
  begin
    result = input_0 & {27{sel[0]}};
    result = result | (input_1 & {27{sel[1]}});
    result = result | (input_2 & {27{sel[2]}});
    result = result | (input_3 & {27{sel[3]}});
    result = result | (input_4 & {27{sel[4]}});
    result = result | (input_5 & {27{sel[5]}});
    result = result | (input_6 & {27{sel[6]}});
    result = result | (input_7 & {27{sel[7]}});
    MUX1HOT_v_27_8_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_4_2;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [3:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    result = result | (input_3 & {2{sel[3]}});
    MUX1HOT_v_2_4_2 = result;
  end
  endfunction


  function automatic [30:0] MUX1HOT_v_31_3_2;
    input [30:0] input_2;
    input [30:0] input_1;
    input [30:0] input_0;
    input [2:0] sel;
    reg [30:0] result;
  begin
    result = input_0 & {31{sel[0]}};
    result = result | (input_1 & {31{sel[1]}});
    result = result | (input_2 & {31{sel[2]}});
    MUX1HOT_v_31_3_2 = result;
  end
  endfunction


  function automatic [30:0] MUX1HOT_v_31_4_2;
    input [30:0] input_3;
    input [30:0] input_2;
    input [30:0] input_1;
    input [30:0] input_0;
    input [3:0] sel;
    reg [30:0] result;
  begin
    result = input_0 & {31{sel[0]}};
    result = result | (input_1 & {31{sel[1]}});
    result = result | (input_2 & {31{sel[2]}});
    result = result | (input_3 & {31{sel[3]}});
    MUX1HOT_v_31_4_2 = result;
  end
  endfunction


  function automatic [30:0] MUX1HOT_v_31_5_2;
    input [30:0] input_4;
    input [30:0] input_3;
    input [30:0] input_2;
    input [30:0] input_1;
    input [30:0] input_0;
    input [4:0] sel;
    reg [30:0] result;
  begin
    result = input_0 & {31{sel[0]}};
    result = result | (input_1 & {31{sel[1]}});
    result = result | (input_2 & {31{sel[2]}});
    result = result | (input_3 & {31{sel[3]}});
    result = result | (input_4 & {31{sel[4]}});
    MUX1HOT_v_31_5_2 = result;
  end
  endfunction


  function automatic [30:0] MUX1HOT_v_31_8_2;
    input [30:0] input_7;
    input [30:0] input_6;
    input [30:0] input_5;
    input [30:0] input_4;
    input [30:0] input_3;
    input [30:0] input_2;
    input [30:0] input_1;
    input [30:0] input_0;
    input [7:0] sel;
    reg [30:0] result;
  begin
    result = input_0 & {31{sel[0]}};
    result = result | (input_1 & {31{sel[1]}});
    result = result | (input_2 & {31{sel[2]}});
    result = result | (input_3 & {31{sel[3]}});
    result = result | (input_4 & {31{sel[4]}});
    result = result | (input_5 & {31{sel[5]}});
    result = result | (input_6 & {31{sel[6]}});
    result = result | (input_7 & {31{sel[7]}});
    MUX1HOT_v_31_8_2 = result;
  end
  endfunction


  function automatic [45:0] MUX1HOT_v_46_4_2;
    input [45:0] input_3;
    input [45:0] input_2;
    input [45:0] input_1;
    input [45:0] input_0;
    input [3:0] sel;
    reg [45:0] result;
  begin
    result = input_0 & {46{sel[0]}};
    result = result | (input_1 & {46{sel[1]}});
    result = result | (input_2 & {46{sel[2]}});
    result = result | (input_3 & {46{sel[3]}});
    MUX1HOT_v_46_4_2 = result;
  end
  endfunction


  function automatic [48:0] MUX1HOT_v_49_3_2;
    input [48:0] input_2;
    input [48:0] input_1;
    input [48:0] input_0;
    input [2:0] sel;
    reg [48:0] result;
  begin
    result = input_0 & {49{sel[0]}};
    result = result | (input_1 & {49{sel[1]}});
    result = result | (input_2 & {49{sel[2]}});
    MUX1HOT_v_49_3_2 = result;
  end
  endfunction


  function automatic [48:0] MUX1HOT_v_49_5_2;
    input [48:0] input_4;
    input [48:0] input_3;
    input [48:0] input_2;
    input [48:0] input_1;
    input [48:0] input_0;
    input [4:0] sel;
    reg [48:0] result;
  begin
    result = input_0 & {49{sel[0]}};
    result = result | (input_1 & {49{sel[1]}});
    result = result | (input_2 & {49{sel[2]}});
    result = result | (input_3 & {49{sel[3]}});
    result = result | (input_4 & {49{sel[4]}});
    MUX1HOT_v_49_5_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_3_2;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [2:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    MUX1HOT_v_5_3_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_4_2;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [3:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    result = result | (input_3 & {5{sel[3]}});
    MUX1HOT_v_5_4_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_4_2;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [3:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | (input_1 & {6{sel[1]}});
    result = result | (input_2 & {6{sel[2]}});
    result = result | (input_3 & {6{sel[3]}});
    MUX1HOT_v_6_4_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_4_2;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [3:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    result = result | (input_3 & {8{sel[3]}});
    MUX1HOT_v_8_4_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_4_2;
    input  input_0;
    input  input_1;
    input  input_2;
    input  input_3;
    input [1:0] sel;
    reg  result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      2'b10 : begin
        result = input_2;
      end
      default : begin
        result = input_3;
      end
    endcase
    MUX_s_1_4_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_64_2;
    input  input_0;
    input  input_1;
    input  input_2;
    input  input_3;
    input  input_4;
    input  input_5;
    input  input_6;
    input  input_7;
    input  input_8;
    input  input_9;
    input  input_10;
    input  input_11;
    input  input_12;
    input  input_13;
    input  input_14;
    input  input_15;
    input  input_16;
    input  input_17;
    input  input_18;
    input  input_19;
    input  input_20;
    input  input_21;
    input  input_22;
    input  input_23;
    input  input_24;
    input  input_25;
    input  input_26;
    input  input_27;
    input  input_28;
    input  input_29;
    input  input_30;
    input  input_31;
    input  input_32;
    input  input_33;
    input  input_34;
    input  input_35;
    input  input_36;
    input  input_37;
    input  input_38;
    input  input_39;
    input  input_40;
    input  input_41;
    input  input_42;
    input  input_43;
    input  input_44;
    input  input_45;
    input  input_46;
    input  input_47;
    input  input_48;
    input  input_49;
    input  input_50;
    input  input_51;
    input  input_52;
    input  input_53;
    input  input_54;
    input  input_55;
    input  input_56;
    input  input_57;
    input  input_58;
    input  input_59;
    input  input_60;
    input  input_61;
    input  input_62;
    input  input_63;
    input [5:0] sel;
    reg  result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      6'b110111 : begin
        result = input_55;
      end
      6'b111000 : begin
        result = input_56;
      end
      6'b111001 : begin
        result = input_57;
      end
      6'b111010 : begin
        result = input_58;
      end
      6'b111011 : begin
        result = input_59;
      end
      6'b111100 : begin
        result = input_60;
      end
      6'b111101 : begin
        result = input_61;
      end
      6'b111110 : begin
        result = input_62;
      end
      default : begin
        result = input_63;
      end
    endcase
    MUX_s_1_64_2 = result;
  end
  endfunction


  function automatic [25:0] MUX_v_26_2_2;
    input [25:0] input_0;
    input [25:0] input_1;
    input  sel;
    reg [25:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_26_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input  sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_32_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [1:0] input_2;
    input [1:0] input_3;
    input [1:0] input_4;
    input [1:0] input_5;
    input [1:0] input_6;
    input [1:0] input_7;
    input [1:0] input_8;
    input [1:0] input_9;
    input [1:0] input_10;
    input [1:0] input_11;
    input [1:0] input_12;
    input [1:0] input_13;
    input [1:0] input_14;
    input [1:0] input_15;
    input [1:0] input_16;
    input [1:0] input_17;
    input [1:0] input_18;
    input [1:0] input_19;
    input [1:0] input_20;
    input [1:0] input_21;
    input [1:0] input_22;
    input [1:0] input_23;
    input [1:0] input_24;
    input [1:0] input_25;
    input [1:0] input_26;
    input [1:0] input_27;
    input [1:0] input_28;
    input [1:0] input_29;
    input [1:0] input_30;
    input [1:0] input_31;
    input [4:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      5'b00000 : begin
        result = input_0;
      end
      5'b00001 : begin
        result = input_1;
      end
      5'b00010 : begin
        result = input_2;
      end
      5'b00011 : begin
        result = input_3;
      end
      5'b00100 : begin
        result = input_4;
      end
      5'b00101 : begin
        result = input_5;
      end
      5'b00110 : begin
        result = input_6;
      end
      5'b00111 : begin
        result = input_7;
      end
      5'b01000 : begin
        result = input_8;
      end
      5'b01001 : begin
        result = input_9;
      end
      5'b01010 : begin
        result = input_10;
      end
      5'b01011 : begin
        result = input_11;
      end
      5'b01100 : begin
        result = input_12;
      end
      5'b01101 : begin
        result = input_13;
      end
      5'b01110 : begin
        result = input_14;
      end
      5'b01111 : begin
        result = input_15;
      end
      5'b10000 : begin
        result = input_16;
      end
      5'b10001 : begin
        result = input_17;
      end
      5'b10010 : begin
        result = input_18;
      end
      5'b10011 : begin
        result = input_19;
      end
      5'b10100 : begin
        result = input_20;
      end
      5'b10101 : begin
        result = input_21;
      end
      5'b10110 : begin
        result = input_22;
      end
      5'b10111 : begin
        result = input_23;
      end
      5'b11000 : begin
        result = input_24;
      end
      5'b11001 : begin
        result = input_25;
      end
      5'b11010 : begin
        result = input_26;
      end
      5'b11011 : begin
        result = input_27;
      end
      5'b11100 : begin
        result = input_28;
      end
      5'b11101 : begin
        result = input_29;
      end
      5'b11110 : begin
        result = input_30;
      end
      default : begin
        result = input_31;
      end
    endcase
    MUX_v_2_32_2 = result;
  end
  endfunction


  function automatic [30:0] MUX_v_31_2_2;
    input [30:0] input_0;
    input [30:0] input_1;
    input  sel;
    reg [30:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_31_2_2 = result;
  end
  endfunction


  function automatic [30:0] MUX_v_31_4_2;
    input [30:0] input_0;
    input [30:0] input_1;
    input [30:0] input_2;
    input [30:0] input_3;
    input [1:0] sel;
    reg [30:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      2'b10 : begin
        result = input_2;
      end
      default : begin
        result = input_3;
      end
    endcase
    MUX_v_31_4_2 = result;
  end
  endfunction


  function automatic [30:0] MUX_v_31_64_2;
    input [30:0] input_0;
    input [30:0] input_1;
    input [30:0] input_2;
    input [30:0] input_3;
    input [30:0] input_4;
    input [30:0] input_5;
    input [30:0] input_6;
    input [30:0] input_7;
    input [30:0] input_8;
    input [30:0] input_9;
    input [30:0] input_10;
    input [30:0] input_11;
    input [30:0] input_12;
    input [30:0] input_13;
    input [30:0] input_14;
    input [30:0] input_15;
    input [30:0] input_16;
    input [30:0] input_17;
    input [30:0] input_18;
    input [30:0] input_19;
    input [30:0] input_20;
    input [30:0] input_21;
    input [30:0] input_22;
    input [30:0] input_23;
    input [30:0] input_24;
    input [30:0] input_25;
    input [30:0] input_26;
    input [30:0] input_27;
    input [30:0] input_28;
    input [30:0] input_29;
    input [30:0] input_30;
    input [30:0] input_31;
    input [30:0] input_32;
    input [30:0] input_33;
    input [30:0] input_34;
    input [30:0] input_35;
    input [30:0] input_36;
    input [30:0] input_37;
    input [30:0] input_38;
    input [30:0] input_39;
    input [30:0] input_40;
    input [30:0] input_41;
    input [30:0] input_42;
    input [30:0] input_43;
    input [30:0] input_44;
    input [30:0] input_45;
    input [30:0] input_46;
    input [30:0] input_47;
    input [30:0] input_48;
    input [30:0] input_49;
    input [30:0] input_50;
    input [30:0] input_51;
    input [30:0] input_52;
    input [30:0] input_53;
    input [30:0] input_54;
    input [30:0] input_55;
    input [30:0] input_56;
    input [30:0] input_57;
    input [30:0] input_58;
    input [30:0] input_59;
    input [30:0] input_60;
    input [30:0] input_61;
    input [30:0] input_62;
    input [30:0] input_63;
    input [5:0] sel;
    reg [30:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      6'b110111 : begin
        result = input_55;
      end
      6'b111000 : begin
        result = input_56;
      end
      6'b111001 : begin
        result = input_57;
      end
      6'b111010 : begin
        result = input_58;
      end
      6'b111011 : begin
        result = input_59;
      end
      6'b111100 : begin
        result = input_60;
      end
      6'b111101 : begin
        result = input_61;
      end
      6'b111110 : begin
        result = input_62;
      end
      default : begin
        result = input_63;
      end
    endcase
    MUX_v_31_64_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_16_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [31:0] input_3;
    input [31:0] input_4;
    input [31:0] input_5;
    input [31:0] input_6;
    input [31:0] input_7;
    input [31:0] input_8;
    input [31:0] input_9;
    input [31:0] input_10;
    input [31:0] input_11;
    input [31:0] input_12;
    input [31:0] input_13;
    input [31:0] input_14;
    input [31:0] input_15;
    input [3:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      4'b0000 : begin
        result = input_0;
      end
      4'b0001 : begin
        result = input_1;
      end
      4'b0010 : begin
        result = input_2;
      end
      4'b0011 : begin
        result = input_3;
      end
      4'b0100 : begin
        result = input_4;
      end
      4'b0101 : begin
        result = input_5;
      end
      4'b0110 : begin
        result = input_6;
      end
      4'b0111 : begin
        result = input_7;
      end
      4'b1000 : begin
        result = input_8;
      end
      4'b1001 : begin
        result = input_9;
      end
      4'b1010 : begin
        result = input_10;
      end
      4'b1011 : begin
        result = input_11;
      end
      4'b1100 : begin
        result = input_12;
      end
      4'b1101 : begin
        result = input_13;
      end
      4'b1110 : begin
        result = input_14;
      end
      default : begin
        result = input_15;
      end
    endcase
    MUX_v_32_16_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input  sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_32_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [31:0] input_3;
    input [31:0] input_4;
    input [31:0] input_5;
    input [31:0] input_6;
    input [31:0] input_7;
    input [31:0] input_8;
    input [31:0] input_9;
    input [31:0] input_10;
    input [31:0] input_11;
    input [31:0] input_12;
    input [31:0] input_13;
    input [31:0] input_14;
    input [31:0] input_15;
    input [31:0] input_16;
    input [31:0] input_17;
    input [31:0] input_18;
    input [31:0] input_19;
    input [31:0] input_20;
    input [31:0] input_21;
    input [31:0] input_22;
    input [31:0] input_23;
    input [31:0] input_24;
    input [31:0] input_25;
    input [31:0] input_26;
    input [31:0] input_27;
    input [31:0] input_28;
    input [31:0] input_29;
    input [31:0] input_30;
    input [31:0] input_31;
    input [4:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      5'b00000 : begin
        result = input_0;
      end
      5'b00001 : begin
        result = input_1;
      end
      5'b00010 : begin
        result = input_2;
      end
      5'b00011 : begin
        result = input_3;
      end
      5'b00100 : begin
        result = input_4;
      end
      5'b00101 : begin
        result = input_5;
      end
      5'b00110 : begin
        result = input_6;
      end
      5'b00111 : begin
        result = input_7;
      end
      5'b01000 : begin
        result = input_8;
      end
      5'b01001 : begin
        result = input_9;
      end
      5'b01010 : begin
        result = input_10;
      end
      5'b01011 : begin
        result = input_11;
      end
      5'b01100 : begin
        result = input_12;
      end
      5'b01101 : begin
        result = input_13;
      end
      5'b01110 : begin
        result = input_14;
      end
      5'b01111 : begin
        result = input_15;
      end
      5'b10000 : begin
        result = input_16;
      end
      5'b10001 : begin
        result = input_17;
      end
      5'b10010 : begin
        result = input_18;
      end
      5'b10011 : begin
        result = input_19;
      end
      5'b10100 : begin
        result = input_20;
      end
      5'b10101 : begin
        result = input_21;
      end
      5'b10110 : begin
        result = input_22;
      end
      5'b10111 : begin
        result = input_23;
      end
      5'b11000 : begin
        result = input_24;
      end
      5'b11001 : begin
        result = input_25;
      end
      5'b11010 : begin
        result = input_26;
      end
      5'b11011 : begin
        result = input_27;
      end
      5'b11100 : begin
        result = input_28;
      end
      5'b11101 : begin
        result = input_29;
      end
      5'b11110 : begin
        result = input_30;
      end
      default : begin
        result = input_31;
      end
    endcase
    MUX_v_32_32_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input  sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [48:0] MUX_v_49_2_2;
    input [48:0] input_0;
    input [48:0] input_1;
    input  sel;
    reg [48:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_49_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input  sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input  sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input  sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input  sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_32_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [7:0] input_2;
    input [7:0] input_3;
    input [7:0] input_4;
    input [7:0] input_5;
    input [7:0] input_6;
    input [7:0] input_7;
    input [7:0] input_8;
    input [7:0] input_9;
    input [7:0] input_10;
    input [7:0] input_11;
    input [7:0] input_12;
    input [7:0] input_13;
    input [7:0] input_14;
    input [7:0] input_15;
    input [7:0] input_16;
    input [7:0] input_17;
    input [7:0] input_18;
    input [7:0] input_19;
    input [7:0] input_20;
    input [7:0] input_21;
    input [7:0] input_22;
    input [7:0] input_23;
    input [7:0] input_24;
    input [7:0] input_25;
    input [7:0] input_26;
    input [7:0] input_27;
    input [7:0] input_28;
    input [7:0] input_29;
    input [7:0] input_30;
    input [7:0] input_31;
    input [4:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      5'b00000 : begin
        result = input_0;
      end
      5'b00001 : begin
        result = input_1;
      end
      5'b00010 : begin
        result = input_2;
      end
      5'b00011 : begin
        result = input_3;
      end
      5'b00100 : begin
        result = input_4;
      end
      5'b00101 : begin
        result = input_5;
      end
      5'b00110 : begin
        result = input_6;
      end
      5'b00111 : begin
        result = input_7;
      end
      5'b01000 : begin
        result = input_8;
      end
      5'b01001 : begin
        result = input_9;
      end
      5'b01010 : begin
        result = input_10;
      end
      5'b01011 : begin
        result = input_11;
      end
      5'b01100 : begin
        result = input_12;
      end
      5'b01101 : begin
        result = input_13;
      end
      5'b01110 : begin
        result = input_14;
      end
      5'b01111 : begin
        result = input_15;
      end
      5'b10000 : begin
        result = input_16;
      end
      5'b10001 : begin
        result = input_17;
      end
      5'b10010 : begin
        result = input_18;
      end
      5'b10011 : begin
        result = input_19;
      end
      5'b10100 : begin
        result = input_20;
      end
      5'b10101 : begin
        result = input_21;
      end
      5'b10110 : begin
        result = input_22;
      end
      5'b10111 : begin
        result = input_23;
      end
      5'b11000 : begin
        result = input_24;
      end
      5'b11001 : begin
        result = input_25;
      end
      5'b11010 : begin
        result = input_26;
      end
      5'b11011 : begin
        result = input_27;
      end
      5'b11100 : begin
        result = input_28;
      end
      5'b11101 : begin
        result = input_29;
      end
      5'b11110 : begin
        result = input_30;
      end
      default : begin
        result = input_31;
      end
    endcase
    MUX_v_8_32_2 = result;
  end
  endfunction


  function automatic [27:0] readslicef_29_28_1;
    input [28:0] vector;
    reg [28:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_29_28_1 = tmp[27:0];
  end
  endfunction


  function automatic [28:0] readslicef_30_29_1;
    input [29:0] vector;
    reg [29:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_30_29_1 = tmp[28:0];
  end
  endfunction


  function automatic [1:0] signext_2_1;
    input  vector;
  begin
    signext_2_1= {{1{vector}}, vector};
  end
  endfunction


  function automatic [31:0] signext_32_1;
    input  vector;
  begin
    signext_32_1= {{31{vector}}, vector};
  end
  endfunction


  function automatic [48:0] signext_49_47;
    input [46:0] vector;
  begin
    signext_49_47= {{2{vector[46]}}, vector};
  end
  endfunction


  function automatic [4:0] signext_5_1;
    input  vector;
  begin
    signext_5_1= {{4{vector}}, vector};
  end
  endfunction


  function automatic [28:0] conv_s2s_26_29 ;
    input [25:0]  vector ;
  begin
    conv_s2s_26_29 = {{3{vector[25]}}, vector};
  end
  endfunction


  function automatic [30:0] conv_s2s_26_31 ;
    input [25:0]  vector ;
  begin
    conv_s2s_26_31 = {{5{vector[25]}}, vector};
  end
  endfunction


  function automatic [29:0] conv_s2s_27_30 ;
    input [26:0]  vector ;
  begin
    conv_s2s_27_30 = {{3{vector[26]}}, vector};
  end
  endfunction


  function automatic [28:0] conv_s2s_28_29 ;
    input [27:0]  vector ;
  begin
    conv_s2s_28_29 = {vector[27], vector};
  end
  endfunction


  function automatic [29:0] conv_s2s_29_30 ;
    input [28:0]  vector ;
  begin
    conv_s2s_29_30 = {vector[28], vector};
  end
  endfunction


  function automatic [30:0] conv_s2s_30_31 ;
    input [29:0]  vector ;
  begin
    conv_s2s_30_31 = {vector[29], vector};
  end
  endfunction


  function automatic [28:0] conv_s2u_26_29 ;
    input [25:0]  vector ;
  begin
    conv_s2u_26_29 = {{3{vector[25]}}, vector};
  end
  endfunction


  function automatic [29:0] conv_s2u_27_30 ;
    input [26:0]  vector ;
  begin
    conv_s2u_27_30 = {{3{vector[26]}}, vector};
  end
  endfunction


  function automatic [28:0] conv_s2u_28_29 ;
    input [27:0]  vector ;
  begin
    conv_s2u_28_29 = {vector[27], vector};
  end
  endfunction


  function automatic [29:0] conv_s2u_29_30 ;
    input [28:0]  vector ;
  begin
    conv_s2u_29_30 = {vector[28], vector};
  end
  endfunction


  function automatic [4:0] conv_u2s_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2s_4_5 =  {1'b0, vector};
  end
  endfunction


  function automatic [6:0] conv_u2s_6_7 ;
    input [5:0]  vector ;
  begin
    conv_u2s_6_7 =  {1'b0, vector};
  end
  endfunction


  function automatic [8:0] conv_u2s_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2s_8_9 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit
// ------------------------------------------------------------------


module ActUnit (
  clk, rst, start_vld, start_rdy, start_dat, act_port_vld, act_port_rdy, act_port_dat,
      rva_in_vld, rva_in_rdy, rva_in_dat, rva_out_vld, rva_out_rdy, rva_out_dat,
      output_port_vld, output_port_rdy, output_port_dat, done_vld, done_rdy, done_dat
);
  input clk;
  input rst;
  input start_vld;
  output start_rdy;
  input start_dat;
  input act_port_vld;
  output act_port_rdy;
  input [511:0] act_port_dat;
  input rva_in_vld;
  output rva_in_rdy;
  input [600:0] rva_in_dat;
  output rva_out_vld;
  input rva_out_rdy;
  output [511:0] rva_out_dat;
  output output_port_vld;
  input output_port_rdy;
  output [521:0] output_port_dat;
  output done_vld;
  input done_rdy;
  output done_dat;



  // Interconnect Declarations for Component Instantiations 
  ActUnit_ActUnit_ActUnitRun ActUnit_ActUnitRun_inst (
      .clk(clk),
      .rst(rst),
      .start_vld(start_vld),
      .start_rdy(start_rdy),
      .start_dat(start_dat),
      .act_port_vld(act_port_vld),
      .act_port_rdy(act_port_rdy),
      .act_port_dat(act_port_dat),
      .rva_in_vld(rva_in_vld),
      .rva_in_rdy(rva_in_rdy),
      .rva_in_dat(rva_in_dat),
      .rva_out_vld(rva_out_vld),
      .rva_out_rdy(rva_out_rdy),
      .rva_out_dat(rva_out_dat),
      .output_port_vld(output_port_vld),
      .output_port_rdy(output_port_rdy),
      .output_port_dat(output_port_dat),
      .done_vld(done_vld),
      .done_rdy(done_rdy),
      .done_dat(done_dat)
    );
endmodule



