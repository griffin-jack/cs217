
//------> ./ActUnit_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ActUnit_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ./ActUnit_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ActUnit_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./ActUnit_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   code@iron-06
//  Generated date: Mon Jan 26 19:49:32 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_core
// ------------------------------------------------------------------


module ActUnit_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_core
    (
  this_vld, this_rdy, this_dat, data_data_rsc_z, data_addr_rsc_z, data_rw_rsc_z,
      return_rsc_z, ccs_ccore_start_rsc_dat, ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  reg this_rdy;
  input [600:0] this_dat;
  output [511:0] data_data_rsc_z;
  output [23:0] data_addr_rsc_z;
  output data_rw_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations
  wire [511:0] nl_data_data_rsci_d;
  assign nl_data_data_rsci_d = this_dat[511:0];
  wire [23:0] nl_data_addr_rsci_d;
  assign nl_data_addr_rsci_d = this_dat[535:512];
  wire  nl_data_rw_rsci_d;
  assign nl_data_rw_rsci_d = this_dat[600];
  ActUnit_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd1),
  .width(32'sd512)) data_data_rsci (
      .d(nl_data_data_rsci_d[511:0]),
      .z(data_data_rsc_z)
    );
  ActUnit_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd2),
  .width(32'sd24)) data_addr_rsci (
      .d(nl_data_addr_rsci_d[23:0]),
      .z(data_addr_rsc_z)
    );
  ActUnit_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd4),
  .width(32'sd1)) data_rw_rsci (
      .d(nl_data_rw_rsci_d),
      .z(data_rw_rsc_z)
    );
  ActUnit_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd6),
  .width(32'sd1)) return_rsci (
      .d(this_vld),
      .z(return_rsc_z)
    );
  ActUnit_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1
      #(.rscid(32'sd58),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_rdy <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB
// ------------------------------------------------------------------


module ActUnit_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB
    (
  this_vld, this_rdy, this_dat, data_data_rsc_z, data_addr_rsc_z, data_rw_rsc_z,
      return_rsc_z, ccs_ccore_start_rsc_dat, ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  input [600:0] this_dat;
  output [511:0] data_data_rsc_z;
  output [23:0] data_addr_rsc_z;
  output data_rw_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  ActUnit_Connections_InBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Writecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_core
      Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .data_data_rsc_z(data_data_rsc_z),
      .data_addr_rsc_z(data_addr_rsc_z),
      .data_rw_rsc_z(data_rw_rsc_z),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./ActUnit_Connections_InBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ActUnit_Connections_InBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ./ActUnit_Connections_InBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ActUnit_Connections_InBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./ActUnit_Connections_InBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_PopNB.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   code@iron-06
//  Generated date: Mon Jan 26 19:49:30 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_spec_ActVectorType_Connections_SYN_PORT_PopNB_core
// ------------------------------------------------------------------


module ActUnit_Connections_InBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_spec_ActVectorType_Connections_SYN_PORT_PopNB_core
    (
  this_vld, this_rdy, this_dat, data_data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  reg this_rdy;
  input [511:0] this_dat;
  output [511:0] data_data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations
  ActUnit_Connections_InBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd7),
  .width(32'sd512)) data_data_rsci (
      .d(this_dat),
      .z(data_data_rsc_z)
    );
  ActUnit_Connections_InBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd9),
  .width(32'sd1)) return_rsci (
      .d(this_vld),
      .z(return_rsc_z)
    );
  ActUnit_Connections_InBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1
      #(.rscid(32'sd57),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_rdy <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_spec_ActVectorType_Connections_SYN_PORT_PopNB
// ------------------------------------------------------------------


module ActUnit_Connections_InBlocking_spec_ActVectorType_Connections_SYN_PORT_PopNB (
  this_vld, this_rdy, this_dat, data_data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  input [511:0] this_dat;
  output [511:0] data_data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  ActUnit_Connections_InBlockingless_spec_ActVectorTypecomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_spec_ActVectorType_Connections_SYN_PORT_PopNB_core
      Connections_InBlocking_spec_ActVectorType_Connections_SYN_PORT_PopNB_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .data_data_rsc_z(data_data_rsc_z),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./ActUnit_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ActUnit_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./ActUnit_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module ActUnit_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./ActUnit_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   code@iron-06
//  Generated date: Mon Jan 26 19:49:27 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module ActUnit_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push_core
    (
  this_vld, this_rdy, this_dat, m_data_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  reg this_vld;
  input this_rdy;
  output [511:0] this_dat;
  reg [511:0] this_dat;
  input [511:0] m_data_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire [511:0] m_data_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  wire and_dcpl;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_4_cse;
  wire this_vld_mx0c1;


  // Interconnect Declarations for Component Instantiations
  wire  nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  ActUnit_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd11),
  .width(32'sd512)) m_data_rsci (
      .dat(m_data_rsc_dat),
      .idat(m_data_rsci_idat)
    );
  ActUnit_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd56),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  ActUnit_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1
      #(.rscid(32'sd61)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld)
    );
  assign or_4_cse = ccs_ccore_start_rsci_idat | and_dcpl;
  assign and_dcpl = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_rdy);
  assign this_vld_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_vld <= 1'b0;
    end
    else if ( or_4_cse | this_vld_mx0c1 ) begin
      this_vld <= ~ this_vld_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_dat <= 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~(and_dcpl | (~ ccs_ccore_start_rsci_idat)) ) begin
      this_dat <= m_data_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_4_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module ActUnit_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push
    (
  this_vld, this_rdy, this_dat, m_data_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  input this_rdy;
  output [511:0] this_dat;
  input [511:0] m_data_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  ActUnit_Connections_OutBlockingless_RVSinkless_spec_Axi_rvaCfggreater_Readcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push_core
      Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .m_data_rsc_dat(m_data_rsc_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./ActUnit_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ActUnit_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ./ActUnit_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ActUnit_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./ActUnit_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   code@iron-06
//  Generated date: Mon Jan 26 19:49:25 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_core
// ------------------------------------------------------------------


module ActUnit_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_core
    (
  this_vld, this_rdy, this_dat, data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  reg this_rdy;
  input this_dat;
  output data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations
  ActUnit_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd12),
  .width(32'sd1)) data_rsci (
      .d(this_dat),
      .z(data_rsc_z)
    );
  ActUnit_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_mgc_out_dreg_v2
      #(.rscid(32'sd14),
  .width(32'sd1)) return_rsci (
      .d(this_vld),
      .z(return_rsc_z)
    );
  ActUnit_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_ccs_in_v1
      #(.rscid(32'sd55),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_rdy <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_bool_Connections_SYN_PORT_PopNB
// ------------------------------------------------------------------


module ActUnit_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB (
  this_vld, this_rdy, this_dat, data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  input this_dat;
  output data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  ActUnit_Connections_InBlockingless_boolcomma_Connections_SYN_PORTgreater_PopNB_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_core
      Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_core_inst (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .data_rsc_z(data_rsc_z),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./ActUnit_Connections_OutBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ActUnit_Connections_OutBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./ActUnit_Connections_OutBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module ActUnit_Connections_OutBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./ActUnit_Connections_OutBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_Push.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   code@iron-06
//  Generated date: Mon Jan 26 19:49:23 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_spec_StreamType_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module ActUnit_Connections_OutBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_spec_StreamType_Connections_SYN_PORT_Push_core
    (
  this_vld, this_rdy, this_dat, m_data_data_rsc_dat, m_logical_addr_rsc_dat, ccs_ccore_start_rsc_dat,
      ccs_ccore_done_sync_vld, ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  reg this_vld;
  input this_rdy;
  output [521:0] this_dat;
  input [511:0] m_data_data_rsc_dat;
  input [7:0] m_logical_addr_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire [511:0] m_data_data_rsci_idat;
  wire [7:0] m_logical_addr_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  reg [7:0] m_logical_addr_buf_lpi_1_dfm;
  reg [511:0] m_data_data_buf_lpi_1_dfm;
  wire and_dcpl;
  wire or_dcpl_2;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_4_cse;
  wire this_vld_mx0c1;


  // Interconnect Declarations for Component Instantiations
  wire  nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  ActUnit_Connections_OutBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd15),
  .width(32'sd512)) m_data_data_rsci (
      .dat(m_data_data_rsc_dat),
      .idat(m_data_data_rsci_idat)
    );
  ActUnit_Connections_OutBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd17),
  .width(32'sd8)) m_logical_addr_rsci (
      .dat(m_logical_addr_rsc_dat),
      .idat(m_logical_addr_rsci_idat)
    );
  ActUnit_Connections_OutBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd54),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  ActUnit_Connections_OutBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1
      #(.rscid(32'sd60)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld)
    );
  assign this_dat = {m_logical_addr_buf_lpi_1_dfm , 2'b00 , m_data_data_buf_lpi_1_dfm};
  assign or_4_cse = ccs_ccore_start_rsci_idat | and_dcpl;
  assign and_dcpl = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_rdy);
  assign or_dcpl_2 = and_dcpl | (~ ccs_ccore_start_rsci_idat);
  assign this_vld_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_vld <= 1'b0;
    end
    else if ( or_4_cse | this_vld_mx0c1 ) begin
      this_vld <= ~ this_vld_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      m_logical_addr_buf_lpi_1_dfm <= 8'b00000000;
    end
    else if ( ~ or_dcpl_2 ) begin
      m_logical_addr_buf_lpi_1_dfm <= m_logical_addr_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      m_data_data_buf_lpi_1_dfm <= 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ or_dcpl_2 ) begin
      m_data_data_buf_lpi_1_dfm <= m_data_data_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_4_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_spec_StreamType_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module ActUnit_Connections_OutBlocking_spec_StreamType_Connections_SYN_PORT_Push (
  this_vld, this_rdy, this_dat, m_data_data_rsc_dat, m_logical_addr_rsc_dat, ccs_ccore_start_rsc_dat,
      ccs_ccore_done_sync_vld, ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  input this_rdy;
  output [521:0] this_dat;
  input [511:0] m_data_data_rsc_dat;
  input [7:0] m_logical_addr_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  ActUnit_Connections_OutBlockingless_spec_StreamTypecomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_spec_StreamType_Connections_SYN_PORT_Push_core
      Connections_OutBlocking_spec_StreamType_Connections_SYN_PORT_Push_core_inst
      (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .m_data_data_rsc_dat(m_data_data_rsc_dat),
      .m_logical_addr_rsc_dat(m_logical_addr_rsc_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./ActUnit_Connections_OutBlockingless_boolcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ActUnit_Connections_OutBlockingless_boolcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./ActUnit_Connections_OutBlockingless_boolcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module ActUnit_Connections_OutBlockingless_boolcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./ActUnit_Connections_OutBlockingless_boolcomma_Connections_SYN_PORTgreater_Push.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   code@iron-06
//  Generated date: Mon Jan 26 19:49:20 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlockingless_boolcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_bool_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module ActUnit_Connections_OutBlockingless_boolcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_bool_Connections_SYN_PORT_Push_core
    (
  this_vld, this_rdy, this_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  reg this_vld;
  input this_rdy;
  output this_dat;
  reg this_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_4_cse;
  wire this_vld_mx0c1;


  // Interconnect Declarations for Component Instantiations
  wire  nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  ActUnit_Connections_OutBlockingless_boolcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd53),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  ActUnit_Connections_OutBlockingless_boolcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1
      #(.rscid(32'sd59)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld)
    );
  assign or_4_cse = ccs_ccore_start_rsci_idat | (io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & (~ this_rdy));
  assign this_vld_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_vld <= 1'b0;
    end
    else if ( or_4_cse | this_vld_mx0c1 ) begin
      this_vld <= ~ this_vld_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_dat <= 1'b0;
    end
    else if ( (~((~ io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1) | this_rdy)) | ccs_ccore_start_rsci_idat
        ) begin
      this_dat <= 1'b1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_4_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_bool_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module ActUnit_Connections_OutBlocking_bool_Connections_SYN_PORT_Push (
  this_vld, this_rdy, this_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  input this_rdy;
  output this_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  ActUnit_Connections_OutBlockingless_boolcomma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_bool_Connections_SYN_PORT_Push_core
      Connections_OutBlocking_bool_Connections_SYN_PORT_Push_core_inst (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./ActUnit_mgc_mul_pipe_beh.v 
//
// File:      $Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_mul_pipe_beh.v
//
// BASELINE:  Catapult-C version 2006b.63
// MODIFIED:  2007-04-03, tnagler
//
// Note: this file uses Verilog2001 features;
//       please enable Verilog2001 in the flow!

module ActUnit_mgc_mul_pipe (a, b, clk, en, a_rst, s_rst, z);

    // Parameters:
    parameter integer width_a = 32'd4;  // input a bit width
    parameter         signd_a =  1'b1;  // input a type (1=signed, 0=unsigned)
    parameter integer width_b = 32'd4;  // input b bit width
    parameter         signd_b =  1'b1;  // input b type (1=signed, 0=unsigned)
    parameter integer width_z = 32'd8;  // result bit width (= width_a + width_b)
    parameter      clock_edge =  1'b0;  // clock polarity (1=posedge, 0=negedge)
    parameter   enable_active =  1'b0;  // enable polarity (1=posedge, 0=negedge)
    parameter    a_rst_active =  1'b1;  // unused
    parameter    s_rst_active =  1'b1;  // unused
    parameter integer  stages = 32'd2;  // number of output registers + 1 (careful!)
    parameter integer n_inreg = 32'd0;  // number of input registers

    localparam integer width_ab = width_a + width_b;  // multiplier result width
    localparam integer n_inreg_min = (n_inreg > 1) ? (n_inreg-1) : 0; // for Synopsys DC

    // I/O ports:
    input  [width_a-1:0] a;      // input A
    input  [width_b-1:0] b;      // input B
    input                clk;    // clock
    input                en;     // enable
    input                a_rst;  // spyglass disable SYNTH_5121,W240
    input                s_rst;  // spyglass disable SYNTH_5121,W240
    output [width_z-1:0] z;      // output


    // Input registers:

    wire [width_a-1:0] a_f;
    wire [width_b-1:0] b_f;

    integer i;

    generate
    if (clock_edge == 1'b0)
    begin: NEG_EDGE1
        case (n_inreg)
        32'd0: begin: B1
            assign a_f = a,
                   b_f = b;
        end
        default: begin: B2
            reg [width_a-1:0] a_reg [n_inreg_min:0];
            reg [width_b-1:0] b_reg [n_inreg_min:0];
            always @(negedge clk)
            if (en == enable_active)
            begin: B21
                a_reg[0] <= a;
                b_reg[0] <= b;
                for (i = 0; i < n_inreg_min; i = i + 1)
                begin: B3
                    a_reg[i+1] <= a_reg[i]; //spyglass disable FlopEConst
                    b_reg[i+1] <= b_reg[i]; //spyglass disable FlopEConst
                end
            end
            assign a_f = a_reg[n_inreg_min],
                   b_f = b_reg[n_inreg_min];
        end
        endcase
    end
    else
    begin: POS_EDGE1
        case (n_inreg)
        32'd0: begin: B1
            assign a_f = a,
                   b_f = b;
        end
        default: begin: B2
            reg [width_a-1:0] a_reg [n_inreg_min:0];
            reg [width_b-1:0] b_reg [n_inreg_min:0];
            always @(posedge clk)
            if (en == enable_active)
            begin: B21
                a_reg[0] <= a; //spyglass disable FlopEConst
                b_reg[0] <= b; //spyglass disable FlopEConst
                for (i = 0; i < n_inreg_min; i = i + 1)
                begin: B3
                    a_reg[i+1] <= a_reg[i]; //spyglass disable FlopEConst
                    b_reg[i+1] <= b_reg[i]; //spyglass disable FlopEConst
                end
            end
            assign a_f = a_reg[n_inreg_min],
                   b_f = b_reg[n_inreg_min];
        end
        endcase
    end
    endgenerate


    // Output:
    wire [width_z-1:0]  xz;

    function signed [width_z-1:0] conv_signed;
      input signed [width_ab-1:0] res;
      conv_signed = res[width_z-1:0];
    endfunction

    generate
      wire signed [width_ab-1:0] res;
      if ( (signd_a == 1'b1) && (signd_b == 1'b1) )
      begin: SIGNED_AB
              assign res = $signed(a_f) * $signed(b_f);
              assign xz = conv_signed(res);
      end
      else if ( (signd_a == 1'b1) && (signd_b == 1'b0) )
      begin: SIGNED_A
              assign res = $signed(a_f) * $signed({1'b0, b_f});
              assign xz = conv_signed(res);
      end
      else if ( (signd_a == 1'b0) && (signd_b == 1'b1) )
      begin: SIGNED_B
              assign res = $signed({1'b0,a_f}) * $signed(b_f);
              assign xz = conv_signed(res);
      end
      else
      begin: UNSIGNED_AB
              assign res = a_f * b_f;
	      assign xz = res[width_z-1:0];
      end
    endgenerate


    // Output registers:

    reg  [width_z-1:0] reg_array[stages-2:0];
    wire [width_z-1:0] z;

    generate
    if (clock_edge == 1'b0)
    begin: NEG_EDGE2
        always @(negedge clk)
        if (en == enable_active)
            for (i = stages-2; i >= 0; i = i-1)
                if (i == 0)
                    reg_array[i] <= xz; //spyglass disable FlopEConst
                else
                    reg_array[i] <= reg_array[i-1]; //spyglass disable FlopEConst
    end
    else
    begin: POS_EDGE2
        always @(posedge clk)
        if (en == enable_active)
            for (i = stages-2; i >= 0; i = i-1)
                if (i == 0)
                    reg_array[i] <= xz; //spyglass disable FlopEConst
                else
                    reg_array[i] <= reg_array[i-1]; //spyglass disable FlopEConst
    end
    endgenerate

    assign z = reg_array[stages-2];
endmodule

//------> ./ActUnit.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
// 
//  Generated by:   code@iron-06
//  Generated date: Thu Jan 29 12:20:14 2026
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_ActUnitRun_fsm
//  FSM Module
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_ActUnitRun_fsm (
  clk, rst, ActUnitRun_wen, fsm_output, while_C_0_tr0, ActUnit_RunInst_case_2_for_C_0_tr0,
      while_C_3_tr0, ActUnit_PushOutput_if_for_C_0_tr0, while_C_5_tr0, ActUnit_RunLoad_if_else_for_C_0_tr0
);
  input clk;
  input rst;
  input ActUnitRun_wen;
  output [3:0] fsm_output;
  reg [3:0] fsm_output;
  input while_C_0_tr0;
  input ActUnit_RunInst_case_2_for_C_0_tr0;
  input while_C_3_tr0;
  input ActUnit_PushOutput_if_for_C_0_tr0;
  input while_C_5_tr0;
  input ActUnit_RunLoad_if_else_for_C_0_tr0;


  // FSM State Type Declaration for ActUnit_ActUnit_ActUnitRun_ActUnitRun_fsm_1
  parameter
    ActUnitRun_rlp_C_0 = 4'd0,
    while_C_0 = 4'd1,
    ActUnit_RunInst_case_2_for_C_0 = 4'd2,
    while_C_1 = 4'd3,
    while_C_2 = 4'd4,
    while_C_3 = 4'd5,
    ActUnit_PushOutput_if_for_C_0 = 4'd6,
    while_C_4 = 4'd7,
    while_C_5 = 4'd8,
    ActUnit_RunLoad_if_else_for_C_0 = 4'd9,
    while_C_6 = 4'd10,
    while_C_7 = 4'd11;

  reg [3:0] state_var;
  reg [3:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : ActUnit_ActUnit_ActUnitRun_ActUnitRun_fsm_1
    case (state_var)
      while_C_0 : begin
        fsm_output = 4'b0001;
        if ( while_C_0_tr0 ) begin
          state_var_NS = while_C_1;
        end
        else begin
          state_var_NS = ActUnit_RunInst_case_2_for_C_0;
        end
      end
      ActUnit_RunInst_case_2_for_C_0 : begin
        fsm_output = 4'b0010;
        if ( ActUnit_RunInst_case_2_for_C_0_tr0 ) begin
          state_var_NS = while_C_1;
        end
        else begin
          state_var_NS = ActUnit_RunInst_case_2_for_C_0;
        end
      end
      while_C_1 : begin
        fsm_output = 4'b0011;
        state_var_NS = while_C_2;
      end
      while_C_2 : begin
        fsm_output = 4'b0100;
        state_var_NS = while_C_3;
      end
      while_C_3 : begin
        fsm_output = 4'b0101;
        if ( while_C_3_tr0 ) begin
          state_var_NS = while_C_4;
        end
        else begin
          state_var_NS = ActUnit_PushOutput_if_for_C_0;
        end
      end
      ActUnit_PushOutput_if_for_C_0 : begin
        fsm_output = 4'b0110;
        if ( ActUnit_PushOutput_if_for_C_0_tr0 ) begin
          state_var_NS = while_C_4;
        end
        else begin
          state_var_NS = ActUnit_PushOutput_if_for_C_0;
        end
      end
      while_C_4 : begin
        fsm_output = 4'b0111;
        state_var_NS = while_C_5;
      end
      while_C_5 : begin
        fsm_output = 4'b1000;
        if ( while_C_5_tr0 ) begin
          state_var_NS = while_C_6;
        end
        else begin
          state_var_NS = ActUnit_RunLoad_if_else_for_C_0;
        end
      end
      ActUnit_RunLoad_if_else_for_C_0 : begin
        fsm_output = 4'b1001;
        if ( ActUnit_RunLoad_if_else_for_C_0_tr0 ) begin
          state_var_NS = while_C_6;
        end
        else begin
          state_var_NS = ActUnit_RunLoad_if_else_for_C_0;
        end
      end
      while_C_6 : begin
        fsm_output = 4'b1010;
        state_var_NS = while_C_7;
      end
      while_C_7 : begin
        fsm_output = 4'b1011;
        state_var_NS = while_C_0;
      end
      // ActUnitRun_rlp_C_0
      default : begin
        fsm_output = 4'b0000;
        state_var_NS = while_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      state_var <= ActUnitRun_rlp_C_0;
    end
    else if ( ActUnitRun_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_staller
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_staller (
  clk, rst, ActUnitRun_wen, ActUnitRun_wten, rva_out_Push_mioi_wen_comp, output_port_Push_mioi_wen_comp,
      done_Push_mioi_wen_comp
);
  input clk;
  input rst;
  output ActUnitRun_wen;
  output ActUnitRun_wten;
  input rva_out_Push_mioi_wen_comp;
  input output_port_Push_mioi_wen_comp;
  input done_Push_mioi_wen_comp;


  // Interconnect Declarations
  reg ActUnitRun_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign ActUnitRun_wen = rva_out_Push_mioi_wen_comp & output_port_Push_mioi_wen_comp
      & done_Push_mioi_wen_comp;
  assign ActUnitRun_wten = ActUnitRun_wten_reg;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnitRun_wten_reg <= 1'b0;
    end
    else begin
      ActUnitRun_wten_reg <= ~ ActUnitRun_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_wait_dp
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_wait_dp (
  ActUnitRun_wen, Gelu_for_1_else_else_else_if_mul_cmp_cgo, Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg,
      Gelu_for_1_else_else_else_if_mul_cmp_en, Gelu_for_1_else_else_else_if_mul_cmp_cgo_1,
      Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_1, Gelu_for_1_else_else_else_if_mul_cmp_1_en,
      Gelu_for_1_else_else_else_if_mul_cmp_cgo_2, Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_2,
      Gelu_for_1_else_else_else_if_mul_cmp_2_en, Gelu_for_1_else_else_else_if_mul_cmp_cgo_3,
      Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_3, Gelu_for_1_else_else_else_if_mul_cmp_3_en,
      Gelu_for_1_else_else_else_if_mul_cmp_cgo_4, Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_4,
      Gelu_for_1_else_else_else_if_mul_cmp_4_en, Gelu_for_1_else_else_else_if_mul_cmp_cgo_5,
      Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_5, Gelu_for_1_else_else_else_if_mul_cmp_5_en,
      Gelu_for_1_else_else_else_if_mul_cmp_cgo_6, Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_6,
      Gelu_for_1_else_else_else_if_mul_cmp_6_en, Gelu_for_1_else_else_else_if_mul_cmp_cgo_7,
      Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_7, Gelu_for_1_else_else_else_if_mul_cmp_7_en,
      Gelu_for_1_else_else_else_if_mul_cmp_cgo_8, Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_8,
      Gelu_for_1_else_else_else_if_mul_cmp_8_en, Gelu_for_1_else_else_else_if_mul_cmp_cgo_9,
      Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_9, Gelu_for_1_else_else_else_if_mul_cmp_9_en,
      Gelu_for_1_else_else_else_if_mul_cmp_cgo_10, Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_10,
      Gelu_for_1_else_else_else_if_mul_cmp_10_en, Gelu_for_1_else_else_else_if_mul_cmp_cgo_11,
      Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_11, Gelu_for_1_else_else_else_if_mul_cmp_11_en,
      Gelu_for_1_else_else_else_if_mul_cmp_cgo_12, Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_12,
      Gelu_for_1_else_else_else_if_mul_cmp_12_en, Gelu_for_1_else_else_else_if_mul_cmp_cgo_13,
      Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_13, Gelu_for_1_else_else_else_if_mul_cmp_13_en,
      Gelu_for_1_else_else_else_if_mul_cmp_cgo_14, Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_14,
      Gelu_for_1_else_else_else_if_mul_cmp_14_en, Gelu_for_1_else_else_else_if_mul_cmp_cgo_15,
      Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_15, Gelu_for_1_else_else_else_if_mul_cmp_15_en,
      Gelu_for_1_else_else_if_mul_cmp_cgo, Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg,
      Gelu_for_1_else_else_if_mul_cmp_en, Gelu_for_1_else_else_if_mul_cmp_cgo_1,
      Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_1, Gelu_for_1_else_else_if_mul_cmp_1_en,
      Gelu_for_1_else_else_if_mul_cmp_cgo_2, Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_2,
      Gelu_for_1_else_else_if_mul_cmp_2_en, Gelu_for_1_else_else_if_mul_cmp_cgo_3,
      Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_3, Gelu_for_1_else_else_if_mul_cmp_3_en,
      Gelu_for_1_else_else_if_mul_cmp_cgo_4, Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_4,
      Gelu_for_1_else_else_if_mul_cmp_4_en, Gelu_for_1_else_else_if_mul_cmp_cgo_5,
      Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_5, Gelu_for_1_else_else_if_mul_cmp_5_en,
      Gelu_for_1_else_else_if_mul_cmp_cgo_6, Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_6,
      Gelu_for_1_else_else_if_mul_cmp_6_en, Gelu_for_1_else_else_if_mul_cmp_cgo_7,
      Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_7, Gelu_for_1_else_else_if_mul_cmp_7_en,
      Gelu_for_1_else_else_if_mul_cmp_cgo_8, Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_8,
      Gelu_for_1_else_else_if_mul_cmp_8_en, Gelu_for_1_else_else_if_mul_cmp_cgo_9,
      Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_9, Gelu_for_1_else_else_if_mul_cmp_9_en,
      Gelu_for_1_else_else_if_mul_cmp_cgo_10, Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_10,
      Gelu_for_1_else_else_if_mul_cmp_10_en, Gelu_for_1_else_else_if_mul_cmp_cgo_11,
      Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_11, Gelu_for_1_else_else_if_mul_cmp_11_en,
      Gelu_for_1_else_else_if_mul_cmp_cgo_12, Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_12,
      Gelu_for_1_else_else_if_mul_cmp_12_en, Gelu_for_1_else_else_if_mul_cmp_cgo_13,
      Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_13, Gelu_for_1_else_else_if_mul_cmp_13_en,
      Gelu_for_1_else_else_if_mul_cmp_cgo_14, Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_14,
      Gelu_for_1_else_else_if_mul_cmp_14_en, Gelu_for_1_else_else_if_mul_cmp_cgo_15,
      Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_15, Gelu_for_1_else_else_if_mul_cmp_15_en,
      Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo, Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_unreg,
      Silu_for_1_else_if_Silu_for_else_if_mul_cmp_en, Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_1,
      Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_unreg_1, Silu_for_1_else_if_Silu_for_else_if_mul_cmp_1_en,
      Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_2, Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_unreg_2,
      Silu_for_1_else_if_Silu_for_else_if_mul_cmp_2_en, Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_3,
      Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_unreg_3, Silu_for_1_else_if_Silu_for_else_if_mul_cmp_3_en,
      Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_4, Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_unreg_4,
      Silu_for_1_else_if_Silu_for_else_if_mul_cmp_4_en, Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_5,
      Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_unreg_5, Silu_for_1_else_if_Silu_for_else_if_mul_cmp_5_en,
      Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_6, Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_unreg_6,
      Silu_for_1_else_if_Silu_for_else_if_mul_cmp_6_en, Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_7,
      Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_unreg_7, Silu_for_1_else_if_Silu_for_else_if_mul_cmp_7_en
);
  input ActUnitRun_wen;
  input Gelu_for_1_else_else_else_if_mul_cmp_cgo;
  input Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg;
  output Gelu_for_1_else_else_else_if_mul_cmp_en;
  input Gelu_for_1_else_else_else_if_mul_cmp_cgo_1;
  input Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_1;
  output Gelu_for_1_else_else_else_if_mul_cmp_1_en;
  input Gelu_for_1_else_else_else_if_mul_cmp_cgo_2;
  input Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_2;
  output Gelu_for_1_else_else_else_if_mul_cmp_2_en;
  input Gelu_for_1_else_else_else_if_mul_cmp_cgo_3;
  input Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_3;
  output Gelu_for_1_else_else_else_if_mul_cmp_3_en;
  input Gelu_for_1_else_else_else_if_mul_cmp_cgo_4;
  input Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_4;
  output Gelu_for_1_else_else_else_if_mul_cmp_4_en;
  input Gelu_for_1_else_else_else_if_mul_cmp_cgo_5;
  input Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_5;
  output Gelu_for_1_else_else_else_if_mul_cmp_5_en;
  input Gelu_for_1_else_else_else_if_mul_cmp_cgo_6;
  input Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_6;
  output Gelu_for_1_else_else_else_if_mul_cmp_6_en;
  input Gelu_for_1_else_else_else_if_mul_cmp_cgo_7;
  input Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_7;
  output Gelu_for_1_else_else_else_if_mul_cmp_7_en;
  input Gelu_for_1_else_else_else_if_mul_cmp_cgo_8;
  input Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_8;
  output Gelu_for_1_else_else_else_if_mul_cmp_8_en;
  input Gelu_for_1_else_else_else_if_mul_cmp_cgo_9;
  input Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_9;
  output Gelu_for_1_else_else_else_if_mul_cmp_9_en;
  input Gelu_for_1_else_else_else_if_mul_cmp_cgo_10;
  input Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_10;
  output Gelu_for_1_else_else_else_if_mul_cmp_10_en;
  input Gelu_for_1_else_else_else_if_mul_cmp_cgo_11;
  input Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_11;
  output Gelu_for_1_else_else_else_if_mul_cmp_11_en;
  input Gelu_for_1_else_else_else_if_mul_cmp_cgo_12;
  input Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_12;
  output Gelu_for_1_else_else_else_if_mul_cmp_12_en;
  input Gelu_for_1_else_else_else_if_mul_cmp_cgo_13;
  input Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_13;
  output Gelu_for_1_else_else_else_if_mul_cmp_13_en;
  input Gelu_for_1_else_else_else_if_mul_cmp_cgo_14;
  input Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_14;
  output Gelu_for_1_else_else_else_if_mul_cmp_14_en;
  input Gelu_for_1_else_else_else_if_mul_cmp_cgo_15;
  input Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_15;
  output Gelu_for_1_else_else_else_if_mul_cmp_15_en;
  input Gelu_for_1_else_else_if_mul_cmp_cgo;
  input Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg;
  output Gelu_for_1_else_else_if_mul_cmp_en;
  input Gelu_for_1_else_else_if_mul_cmp_cgo_1;
  input Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_1;
  output Gelu_for_1_else_else_if_mul_cmp_1_en;
  input Gelu_for_1_else_else_if_mul_cmp_cgo_2;
  input Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_2;
  output Gelu_for_1_else_else_if_mul_cmp_2_en;
  input Gelu_for_1_else_else_if_mul_cmp_cgo_3;
  input Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_3;
  output Gelu_for_1_else_else_if_mul_cmp_3_en;
  input Gelu_for_1_else_else_if_mul_cmp_cgo_4;
  input Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_4;
  output Gelu_for_1_else_else_if_mul_cmp_4_en;
  input Gelu_for_1_else_else_if_mul_cmp_cgo_5;
  input Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_5;
  output Gelu_for_1_else_else_if_mul_cmp_5_en;
  input Gelu_for_1_else_else_if_mul_cmp_cgo_6;
  input Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_6;
  output Gelu_for_1_else_else_if_mul_cmp_6_en;
  input Gelu_for_1_else_else_if_mul_cmp_cgo_7;
  input Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_7;
  output Gelu_for_1_else_else_if_mul_cmp_7_en;
  input Gelu_for_1_else_else_if_mul_cmp_cgo_8;
  input Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_8;
  output Gelu_for_1_else_else_if_mul_cmp_8_en;
  input Gelu_for_1_else_else_if_mul_cmp_cgo_9;
  input Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_9;
  output Gelu_for_1_else_else_if_mul_cmp_9_en;
  input Gelu_for_1_else_else_if_mul_cmp_cgo_10;
  input Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_10;
  output Gelu_for_1_else_else_if_mul_cmp_10_en;
  input Gelu_for_1_else_else_if_mul_cmp_cgo_11;
  input Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_11;
  output Gelu_for_1_else_else_if_mul_cmp_11_en;
  input Gelu_for_1_else_else_if_mul_cmp_cgo_12;
  input Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_12;
  output Gelu_for_1_else_else_if_mul_cmp_12_en;
  input Gelu_for_1_else_else_if_mul_cmp_cgo_13;
  input Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_13;
  output Gelu_for_1_else_else_if_mul_cmp_13_en;
  input Gelu_for_1_else_else_if_mul_cmp_cgo_14;
  input Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_14;
  output Gelu_for_1_else_else_if_mul_cmp_14_en;
  input Gelu_for_1_else_else_if_mul_cmp_cgo_15;
  input Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_15;
  output Gelu_for_1_else_else_if_mul_cmp_15_en;
  input Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo;
  input Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_unreg;
  output Silu_for_1_else_if_Silu_for_else_if_mul_cmp_en;
  input Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_1;
  input Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_unreg_1;
  output Silu_for_1_else_if_Silu_for_else_if_mul_cmp_1_en;
  input Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_2;
  input Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_unreg_2;
  output Silu_for_1_else_if_Silu_for_else_if_mul_cmp_2_en;
  input Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_3;
  input Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_unreg_3;
  output Silu_for_1_else_if_Silu_for_else_if_mul_cmp_3_en;
  input Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_4;
  input Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_unreg_4;
  output Silu_for_1_else_if_Silu_for_else_if_mul_cmp_4_en;
  input Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_5;
  input Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_unreg_5;
  output Silu_for_1_else_if_Silu_for_else_if_mul_cmp_5_en;
  input Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_6;
  input Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_unreg_6;
  output Silu_for_1_else_if_Silu_for_else_if_mul_cmp_6_en;
  input Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_7;
  input Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_unreg_7;
  output Silu_for_1_else_if_Silu_for_else_if_mul_cmp_7_en;



  // Interconnect Declarations for Component Instantiations 
  assign Gelu_for_1_else_else_else_if_mul_cmp_en = ActUnitRun_wen & (Gelu_for_1_else_else_else_if_mul_cmp_cgo
      | Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg);
  assign Gelu_for_1_else_else_else_if_mul_cmp_1_en = ActUnitRun_wen & (Gelu_for_1_else_else_else_if_mul_cmp_cgo_1
      | Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_1);
  assign Gelu_for_1_else_else_else_if_mul_cmp_2_en = ActUnitRun_wen & (Gelu_for_1_else_else_else_if_mul_cmp_cgo_2
      | Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_2);
  assign Gelu_for_1_else_else_else_if_mul_cmp_3_en = ActUnitRun_wen & (Gelu_for_1_else_else_else_if_mul_cmp_cgo_3
      | Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_3);
  assign Gelu_for_1_else_else_else_if_mul_cmp_4_en = ActUnitRun_wen & (Gelu_for_1_else_else_else_if_mul_cmp_cgo_4
      | Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_4);
  assign Gelu_for_1_else_else_else_if_mul_cmp_5_en = ActUnitRun_wen & (Gelu_for_1_else_else_else_if_mul_cmp_cgo_5
      | Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_5);
  assign Gelu_for_1_else_else_else_if_mul_cmp_6_en = ActUnitRun_wen & (Gelu_for_1_else_else_else_if_mul_cmp_cgo_6
      | Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_6);
  assign Gelu_for_1_else_else_else_if_mul_cmp_7_en = ActUnitRun_wen & (Gelu_for_1_else_else_else_if_mul_cmp_cgo_7
      | Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_7);
  assign Gelu_for_1_else_else_else_if_mul_cmp_8_en = ActUnitRun_wen & (Gelu_for_1_else_else_else_if_mul_cmp_cgo_8
      | Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_8);
  assign Gelu_for_1_else_else_else_if_mul_cmp_9_en = ActUnitRun_wen & (Gelu_for_1_else_else_else_if_mul_cmp_cgo_9
      | Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_9);
  assign Gelu_for_1_else_else_else_if_mul_cmp_10_en = ActUnitRun_wen & (Gelu_for_1_else_else_else_if_mul_cmp_cgo_10
      | Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_10);
  assign Gelu_for_1_else_else_else_if_mul_cmp_11_en = ActUnitRun_wen & (Gelu_for_1_else_else_else_if_mul_cmp_cgo_11
      | Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_11);
  assign Gelu_for_1_else_else_else_if_mul_cmp_12_en = ActUnitRun_wen & (Gelu_for_1_else_else_else_if_mul_cmp_cgo_12
      | Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_12);
  assign Gelu_for_1_else_else_else_if_mul_cmp_13_en = ActUnitRun_wen & (Gelu_for_1_else_else_else_if_mul_cmp_cgo_13
      | Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_13);
  assign Gelu_for_1_else_else_else_if_mul_cmp_14_en = ActUnitRun_wen & (Gelu_for_1_else_else_else_if_mul_cmp_cgo_14
      | Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_14);
  assign Gelu_for_1_else_else_else_if_mul_cmp_15_en = ActUnitRun_wen & (Gelu_for_1_else_else_else_if_mul_cmp_cgo_15
      | Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_15);
  assign Gelu_for_1_else_else_if_mul_cmp_en = ActUnitRun_wen & (Gelu_for_1_else_else_if_mul_cmp_cgo
      | Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg);
  assign Gelu_for_1_else_else_if_mul_cmp_1_en = ActUnitRun_wen & (Gelu_for_1_else_else_if_mul_cmp_cgo_1
      | Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_1);
  assign Gelu_for_1_else_else_if_mul_cmp_2_en = ActUnitRun_wen & (Gelu_for_1_else_else_if_mul_cmp_cgo_2
      | Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_2);
  assign Gelu_for_1_else_else_if_mul_cmp_3_en = ActUnitRun_wen & (Gelu_for_1_else_else_if_mul_cmp_cgo_3
      | Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_3);
  assign Gelu_for_1_else_else_if_mul_cmp_4_en = ActUnitRun_wen & (Gelu_for_1_else_else_if_mul_cmp_cgo_4
      | Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_4);
  assign Gelu_for_1_else_else_if_mul_cmp_5_en = ActUnitRun_wen & (Gelu_for_1_else_else_if_mul_cmp_cgo_5
      | Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_5);
  assign Gelu_for_1_else_else_if_mul_cmp_6_en = ActUnitRun_wen & (Gelu_for_1_else_else_if_mul_cmp_cgo_6
      | Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_6);
  assign Gelu_for_1_else_else_if_mul_cmp_7_en = ActUnitRun_wen & (Gelu_for_1_else_else_if_mul_cmp_cgo_7
      | Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_7);
  assign Gelu_for_1_else_else_if_mul_cmp_8_en = ActUnitRun_wen & (Gelu_for_1_else_else_if_mul_cmp_cgo_8
      | Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_8);
  assign Gelu_for_1_else_else_if_mul_cmp_9_en = ActUnitRun_wen & (Gelu_for_1_else_else_if_mul_cmp_cgo_9
      | Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_9);
  assign Gelu_for_1_else_else_if_mul_cmp_10_en = ActUnitRun_wen & (Gelu_for_1_else_else_if_mul_cmp_cgo_10
      | Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_10);
  assign Gelu_for_1_else_else_if_mul_cmp_11_en = ActUnitRun_wen & (Gelu_for_1_else_else_if_mul_cmp_cgo_11
      | Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_11);
  assign Gelu_for_1_else_else_if_mul_cmp_12_en = ActUnitRun_wen & (Gelu_for_1_else_else_if_mul_cmp_cgo_12
      | Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_12);
  assign Gelu_for_1_else_else_if_mul_cmp_13_en = ActUnitRun_wen & (Gelu_for_1_else_else_if_mul_cmp_cgo_13
      | Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_13);
  assign Gelu_for_1_else_else_if_mul_cmp_14_en = ActUnitRun_wen & (Gelu_for_1_else_else_if_mul_cmp_cgo_14
      | Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_14);
  assign Gelu_for_1_else_else_if_mul_cmp_15_en = ActUnitRun_wen & (Gelu_for_1_else_else_if_mul_cmp_cgo_15
      | Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_15);
  assign Silu_for_1_else_if_Silu_for_else_if_mul_cmp_en = ActUnitRun_wen & (Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo
      | Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_unreg);
  assign Silu_for_1_else_if_Silu_for_else_if_mul_cmp_1_en = ActUnitRun_wen & (Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_1
      | Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_unreg_1);
  assign Silu_for_1_else_if_Silu_for_else_if_mul_cmp_2_en = ActUnitRun_wen & (Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_2
      | Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_unreg_2);
  assign Silu_for_1_else_if_Silu_for_else_if_mul_cmp_3_en = ActUnitRun_wen & (Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_3
      | Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_unreg_3);
  assign Silu_for_1_else_if_Silu_for_else_if_mul_cmp_4_en = ActUnitRun_wen & (Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_4
      | Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_unreg_4);
  assign Silu_for_1_else_if_Silu_for_else_if_mul_cmp_5_en = ActUnitRun_wen & (Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_5
      | Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_unreg_5);
  assign Silu_for_1_else_if_Silu_for_else_if_mul_cmp_6_en = ActUnitRun_wen & (Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_6
      | Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_unreg_6);
  assign Silu_for_1_else_if_Silu_for_else_if_mul_cmp_7_en = ActUnitRun_wen & (Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_7
      | Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_unreg_7);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_done_Push_mioi_done_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_done_Push_mioi_done_Push_mio_wait_ctrl (
  ActUnitRun_wten, done_Push_mioi_iswt0, done_Push_mioi_biwt, done_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct,
      done_Push_mioi_ccs_ccore_done_sync_vld, done_Push_mioi_iswt0_pff
);
  input ActUnitRun_wten;
  input done_Push_mioi_iswt0;
  output done_Push_mioi_biwt;
  output done_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct;
  input done_Push_mioi_ccs_ccore_done_sync_vld;
  input done_Push_mioi_iswt0_pff;



  // Interconnect Declarations for Component Instantiations 
  assign done_Push_mioi_biwt = done_Push_mioi_iswt0 & done_Push_mioi_ccs_ccore_done_sync_vld;
  assign done_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct = (~ ActUnitRun_wten)
      & done_Push_mioi_iswt0_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_output_port_Push_mioi_output_port_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_output_port_Push_mioi_output_port_Push_mio_wait_ctrl
    (
  ActUnitRun_wten, output_port_Push_mioi_iswt0, output_port_Push_mioi_biwt, output_port_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct,
      output_port_Push_mioi_ccs_ccore_done_sync_vld, output_port_Push_mioi_iswt0_pff
);
  input ActUnitRun_wten;
  input output_port_Push_mioi_iswt0;
  output output_port_Push_mioi_biwt;
  output output_port_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct;
  input output_port_Push_mioi_ccs_ccore_done_sync_vld;
  input output_port_Push_mioi_iswt0_pff;



  // Interconnect Declarations for Component Instantiations 
  assign output_port_Push_mioi_biwt = output_port_Push_mioi_iswt0 & output_port_Push_mioi_ccs_ccore_done_sync_vld;
  assign output_port_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct = (~ ActUnitRun_wten)
      & output_port_Push_mioi_iswt0_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_start_PopNB_mioi_start_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_start_PopNB_mioi_start_PopNB_mio_wait_dp (
  clk, rst, start_PopNB_mioi_data_rsc_z_mxwt, start_PopNB_mioi_return_rsc_z_mxwt,
      start_PopNB_mioi_biwt, start_PopNB_mioi_bdwt, start_PopNB_mioi_data_rsc_z,
      start_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output start_PopNB_mioi_data_rsc_z_mxwt;
  output start_PopNB_mioi_return_rsc_z_mxwt;
  input start_PopNB_mioi_biwt;
  input start_PopNB_mioi_bdwt;
  input start_PopNB_mioi_data_rsc_z;
  input start_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg start_PopNB_mioi_bcwt;
  reg start_PopNB_mioi_data_rsc_z_bfwt;
  reg start_PopNB_mioi_return_rsc_z_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign start_PopNB_mioi_data_rsc_z_mxwt = MUX_s_1_2_2(start_PopNB_mioi_data_rsc_z,
      start_PopNB_mioi_data_rsc_z_bfwt, start_PopNB_mioi_bcwt);
  assign start_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(start_PopNB_mioi_return_rsc_z,
      start_PopNB_mioi_return_rsc_z_bfwt, start_PopNB_mioi_bcwt);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      start_PopNB_mioi_bcwt <= 1'b0;
    end
    else begin
      start_PopNB_mioi_bcwt <= ~((~(start_PopNB_mioi_bcwt | start_PopNB_mioi_biwt))
          | start_PopNB_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      start_PopNB_mioi_data_rsc_z_bfwt <= 1'b0;
      start_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else if ( start_PopNB_mioi_biwt ) begin
      start_PopNB_mioi_data_rsc_z_bfwt <= start_PopNB_mioi_data_rsc_z;
      start_PopNB_mioi_return_rsc_z_bfwt <= start_PopNB_mioi_return_rsc_z;
    end
  end

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_start_PopNB_mioi_start_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_start_PopNB_mioi_start_PopNB_mio_wait_ctrl (
  ActUnitRun_wen, ActUnitRun_wten, start_PopNB_mioi_oswt, start_PopNB_mioi_biwt,
      start_PopNB_mioi_bdwt, start_PopNB_mioi_biwt_pff, start_PopNB_mioi_oswt_pff
);
  input ActUnitRun_wen;
  input ActUnitRun_wten;
  input start_PopNB_mioi_oswt;
  output start_PopNB_mioi_biwt;
  output start_PopNB_mioi_bdwt;
  output start_PopNB_mioi_biwt_pff;
  input start_PopNB_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign start_PopNB_mioi_bdwt = start_PopNB_mioi_oswt & ActUnitRun_wen;
  assign start_PopNB_mioi_biwt = (~ ActUnitRun_wten) & start_PopNB_mioi_oswt;
  assign start_PopNB_mioi_biwt_pff = ActUnitRun_wen & start_PopNB_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl (
  ActUnitRun_wten, rva_out_Push_mioi_iswt0, rva_out_Push_mioi_biwt, rva_out_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct,
      rva_out_Push_mioi_ccs_ccore_done_sync_vld, rva_out_Push_mioi_iswt0_pff
);
  input ActUnitRun_wten;
  input rva_out_Push_mioi_iswt0;
  output rva_out_Push_mioi_biwt;
  output rva_out_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct;
  input rva_out_Push_mioi_ccs_ccore_done_sync_vld;
  input rva_out_Push_mioi_iswt0_pff;



  // Interconnect Declarations for Component Instantiations 
  assign rva_out_Push_mioi_biwt = rva_out_Push_mioi_iswt0 & rva_out_Push_mioi_ccs_ccore_done_sync_vld;
  assign rva_out_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct = (~ ActUnitRun_wten)
      & rva_out_Push_mioi_iswt0_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_act_port_PopNB_mioi_act_port_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_act_port_PopNB_mioi_act_port_PopNB_mio_wait_dp
    (
  clk, rst, act_port_PopNB_mioi_data_data_rsc_z_mxwt, act_port_PopNB_mioi_return_rsc_z_mxwt,
      act_port_PopNB_mioi_biwt, act_port_PopNB_mioi_bdwt, act_port_PopNB_mioi_data_data_rsc_z,
      act_port_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output [511:0] act_port_PopNB_mioi_data_data_rsc_z_mxwt;
  output act_port_PopNB_mioi_return_rsc_z_mxwt;
  input act_port_PopNB_mioi_biwt;
  input act_port_PopNB_mioi_bdwt;
  input [511:0] act_port_PopNB_mioi_data_data_rsc_z;
  input act_port_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg act_port_PopNB_mioi_bcwt;
  reg [511:0] act_port_PopNB_mioi_data_data_rsc_z_bfwt;
  reg act_port_PopNB_mioi_return_rsc_z_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign act_port_PopNB_mioi_data_data_rsc_z_mxwt = MUX_v_512_2_2(act_port_PopNB_mioi_data_data_rsc_z,
      act_port_PopNB_mioi_data_data_rsc_z_bfwt, act_port_PopNB_mioi_bcwt);
  assign act_port_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(act_port_PopNB_mioi_return_rsc_z,
      act_port_PopNB_mioi_return_rsc_z_bfwt, act_port_PopNB_mioi_bcwt);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_PopNB_mioi_bcwt <= 1'b0;
    end
    else begin
      act_port_PopNB_mioi_bcwt <= ~((~(act_port_PopNB_mioi_bcwt | act_port_PopNB_mioi_biwt))
          | act_port_PopNB_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_PopNB_mioi_data_data_rsc_z_bfwt <= 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      act_port_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else if ( act_port_PopNB_mioi_biwt ) begin
      act_port_PopNB_mioi_data_data_rsc_z_bfwt <= act_port_PopNB_mioi_data_data_rsc_z;
      act_port_PopNB_mioi_return_rsc_z_bfwt <= act_port_PopNB_mioi_return_rsc_z;
    end
  end

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [511:0] MUX_v_512_2_2;
    input [511:0] input_0;
    input [511:0] input_1;
    input  sel;
    reg [511:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_512_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_act_port_PopNB_mioi_act_port_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_act_port_PopNB_mioi_act_port_PopNB_mio_wait_ctrl
    (
  ActUnitRun_wen, ActUnitRun_wten, act_port_PopNB_mioi_oswt, act_port_PopNB_mioi_biwt,
      act_port_PopNB_mioi_bdwt, act_port_PopNB_mioi_biwt_pff, act_port_PopNB_mioi_oswt_pff
);
  input ActUnitRun_wen;
  input ActUnitRun_wten;
  input act_port_PopNB_mioi_oswt;
  output act_port_PopNB_mioi_biwt;
  output act_port_PopNB_mioi_bdwt;
  output act_port_PopNB_mioi_biwt_pff;
  input act_port_PopNB_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign act_port_PopNB_mioi_bdwt = act_port_PopNB_mioi_oswt & ActUnitRun_wen;
  assign act_port_PopNB_mioi_biwt = (~ ActUnitRun_wten) & act_port_PopNB_mioi_oswt;
  assign act_port_PopNB_mioi_biwt_pff = ActUnitRun_wen & act_port_PopNB_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp (
  clk, rst, rva_in_PopNB_mioi_data_data_rsc_z_mxwt, rva_in_PopNB_mioi_data_addr_rsc_z_mxwt,
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt, rva_in_PopNB_mioi_return_rsc_z_mxwt,
      rva_in_PopNB_mioi_biwt, rva_in_PopNB_mioi_bdwt, rva_in_PopNB_mioi_data_data_rsc_z,
      rva_in_PopNB_mioi_data_addr_rsc_z, rva_in_PopNB_mioi_data_rw_rsc_z, rva_in_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output [511:0] rva_in_PopNB_mioi_data_data_rsc_z_mxwt;
  output [11:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt;
  output rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  output rva_in_PopNB_mioi_return_rsc_z_mxwt;
  input rva_in_PopNB_mioi_biwt;
  input rva_in_PopNB_mioi_bdwt;
  input [511:0] rva_in_PopNB_mioi_data_data_rsc_z;
  input [23:0] rva_in_PopNB_mioi_data_addr_rsc_z;
  input rva_in_PopNB_mioi_data_rw_rsc_z;
  input rva_in_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg rva_in_PopNB_mioi_bcwt;
  reg [511:0] rva_in_PopNB_mioi_data_data_rsc_z_bfwt;
  reg rva_in_PopNB_mioi_data_rw_rsc_z_bfwt;
  reg rva_in_PopNB_mioi_return_rsc_z_bfwt;
  reg [3:0] rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_23_20;
  reg [7:0] rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_11_4;

  wire[3:0] ActUnit_DecodeAxi_if_mux_3_nl;
  wire[7:0] ActUnit_DecodeAxi_if_mux_9_nl;

  // Interconnect Declarations for Component Instantiations 
  assign rva_in_PopNB_mioi_data_data_rsc_z_mxwt = MUX_v_512_2_2(rva_in_PopNB_mioi_data_data_rsc_z,
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt, rva_in_PopNB_mioi_bcwt);
  assign rva_in_PopNB_mioi_data_rw_rsc_z_mxwt = MUX_s_1_2_2(rva_in_PopNB_mioi_data_rw_rsc_z,
      rva_in_PopNB_mioi_data_rw_rsc_z_bfwt, rva_in_PopNB_mioi_bcwt);
  assign rva_in_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(rva_in_PopNB_mioi_return_rsc_z,
      rva_in_PopNB_mioi_return_rsc_z_bfwt, rva_in_PopNB_mioi_bcwt);
  assign ActUnit_DecodeAxi_if_mux_3_nl = MUX_v_4_2_2((rva_in_PopNB_mioi_data_addr_rsc_z[23:20]),
      rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_23_20, rva_in_PopNB_mioi_bcwt);
  assign ActUnit_DecodeAxi_if_mux_9_nl = MUX_v_8_2_2((rva_in_PopNB_mioi_data_addr_rsc_z[11:4]),
      rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_11_4, rva_in_PopNB_mioi_bcwt);
  assign rva_in_PopNB_mioi_data_addr_rsc_z_mxwt = {ActUnit_DecodeAxi_if_mux_3_nl
      , ActUnit_DecodeAxi_if_mux_9_nl};
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_PopNB_mioi_bcwt <= 1'b0;
    end
    else begin
      rva_in_PopNB_mioi_bcwt <= ~((~(rva_in_PopNB_mioi_bcwt | rva_in_PopNB_mioi_biwt))
          | rva_in_PopNB_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt <= 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_23_20 <= 4'b0000;
      rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_11_4 <= 8'b00000000;
      rva_in_PopNB_mioi_data_rw_rsc_z_bfwt <= 1'b0;
      rva_in_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else if ( rva_in_PopNB_mioi_biwt ) begin
      rva_in_PopNB_mioi_data_data_rsc_z_bfwt <= rva_in_PopNB_mioi_data_data_rsc_z;
      rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_23_20 <= rva_in_PopNB_mioi_data_addr_rsc_z[23:20];
      rva_in_PopNB_mioi_data_addr_rsc_z_bfwt_11_4 <= rva_in_PopNB_mioi_data_addr_rsc_z[11:4];
      rva_in_PopNB_mioi_data_rw_rsc_z_bfwt <= rva_in_PopNB_mioi_data_rw_rsc_z;
      rva_in_PopNB_mioi_return_rsc_z_bfwt <= rva_in_PopNB_mioi_return_rsc_z;
    end
  end

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input  sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [511:0] MUX_v_512_2_2;
    input [511:0] input_0;
    input [511:0] input_1;
    input  sel;
    reg [511:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_512_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl (
  ActUnitRun_wen, ActUnitRun_wten, rva_in_PopNB_mioi_oswt, rva_in_PopNB_mioi_biwt,
      rva_in_PopNB_mioi_bdwt, rva_in_PopNB_mioi_biwt_pff, rva_in_PopNB_mioi_oswt_pff
);
  input ActUnitRun_wen;
  input ActUnitRun_wten;
  input rva_in_PopNB_mioi_oswt;
  output rva_in_PopNB_mioi_biwt;
  output rva_in_PopNB_mioi_bdwt;
  output rva_in_PopNB_mioi_biwt_pff;
  input rva_in_PopNB_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign rva_in_PopNB_mioi_bdwt = rva_in_PopNB_mioi_oswt & ActUnitRun_wen;
  assign rva_in_PopNB_mioi_biwt = (~ ActUnitRun_wten) & rva_in_PopNB_mioi_oswt;
  assign rva_in_PopNB_mioi_biwt_pff = ActUnitRun_wen & rva_in_PopNB_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_done_Push_mioi
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_done_Push_mioi (
  clk, rst, done_vld, done_rdy, done_dat, ActUnitRun_wten, done_Push_mioi_oswt, done_Push_mioi_wen_comp,
      done_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output done_vld;
  input done_rdy;
  output done_dat;
  input ActUnitRun_wten;
  input done_Push_mioi_oswt;
  output done_Push_mioi_wen_comp;
  input done_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire done_Push_mioi_biwt;
  wire done_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct;
  wire done_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  ActUnit_Connections_OutBlocking_bool_Connections_SYN_PORT_Push  done_Push_mioi
      (
      .this_vld(done_vld),
      .this_rdy(done_rdy),
      .this_dat(done_dat),
      .ccs_ccore_start_rsc_dat(done_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct),
      .ccs_ccore_done_sync_vld(done_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  ActUnit_ActUnit_ActUnitRun_done_Push_mioi_done_Push_mio_wait_ctrl ActUnit_ActUnitRun_done_Push_mioi_done_Push_mio_wait_ctrl_inst
      (
      .ActUnitRun_wten(ActUnitRun_wten),
      .done_Push_mioi_iswt0(done_Push_mioi_oswt),
      .done_Push_mioi_biwt(done_Push_mioi_biwt),
      .done_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct(done_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct),
      .done_Push_mioi_ccs_ccore_done_sync_vld(done_Push_mioi_ccs_ccore_done_sync_vld),
      .done_Push_mioi_iswt0_pff(done_Push_mioi_oswt_pff)
    );
  assign done_Push_mioi_wen_comp = (~ done_Push_mioi_oswt) | done_Push_mioi_biwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_output_port_Push_mioi
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_output_port_Push_mioi (
  clk, rst, output_port_vld, output_port_rdy, output_port_dat, ActUnitRun_wten, output_port_Push_mioi_oswt,
      output_port_Push_mioi_wen_comp, output_port_Push_mioi_m_data_data_rsc_dat_ActUnitRun,
      output_port_Push_mioi_m_logical_addr_rsc_dat_ActUnitRun, output_port_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output output_port_vld;
  input output_port_rdy;
  output [521:0] output_port_dat;
  input ActUnitRun_wten;
  input output_port_Push_mioi_oswt;
  output output_port_Push_mioi_wen_comp;
  input [511:0] output_port_Push_mioi_m_data_data_rsc_dat_ActUnitRun;
  input [7:0] output_port_Push_mioi_m_logical_addr_rsc_dat_ActUnitRun;
  input output_port_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire output_port_Push_mioi_biwt;
  wire output_port_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct;
  wire output_port_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  ActUnit_Connections_OutBlocking_spec_StreamType_Connections_SYN_PORT_Push  output_port_Push_mioi
      (
      .this_vld(output_port_vld),
      .this_rdy(output_port_rdy),
      .this_dat(output_port_dat),
      .m_data_data_rsc_dat(output_port_Push_mioi_m_data_data_rsc_dat_ActUnitRun),
      .m_logical_addr_rsc_dat(output_port_Push_mioi_m_logical_addr_rsc_dat_ActUnitRun),
      .ccs_ccore_start_rsc_dat(output_port_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct),
      .ccs_ccore_done_sync_vld(output_port_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  ActUnit_ActUnit_ActUnitRun_output_port_Push_mioi_output_port_Push_mio_wait_ctrl
      ActUnit_ActUnitRun_output_port_Push_mioi_output_port_Push_mio_wait_ctrl_inst
      (
      .ActUnitRun_wten(ActUnitRun_wten),
      .output_port_Push_mioi_iswt0(output_port_Push_mioi_oswt),
      .output_port_Push_mioi_biwt(output_port_Push_mioi_biwt),
      .output_port_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct(output_port_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct),
      .output_port_Push_mioi_ccs_ccore_done_sync_vld(output_port_Push_mioi_ccs_ccore_done_sync_vld),
      .output_port_Push_mioi_iswt0_pff(output_port_Push_mioi_oswt_pff)
    );
  assign output_port_Push_mioi_wen_comp = (~ output_port_Push_mioi_oswt) | output_port_Push_mioi_biwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_start_PopNB_mioi
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_start_PopNB_mioi (
  clk, rst, start_vld, start_rdy, start_dat, ActUnitRun_wen, ActUnitRun_wten, start_PopNB_mioi_oswt,
      start_PopNB_mioi_data_rsc_z_mxwt, start_PopNB_mioi_return_rsc_z_mxwt, start_PopNB_mioi_oswt_pff
);
  input clk;
  input rst;
  input start_vld;
  output start_rdy;
  input start_dat;
  input ActUnitRun_wen;
  input ActUnitRun_wten;
  input start_PopNB_mioi_oswt;
  output start_PopNB_mioi_data_rsc_z_mxwt;
  output start_PopNB_mioi_return_rsc_z_mxwt;
  input start_PopNB_mioi_oswt_pff;


  // Interconnect Declarations
  wire start_PopNB_mioi_biwt;
  wire start_PopNB_mioi_bdwt;
  wire start_PopNB_mioi_data_rsc_z;
  wire start_PopNB_mioi_return_rsc_z;
  wire start_PopNB_mioi_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  ActUnit_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB  start_PopNB_mioi
      (
      .this_vld(start_vld),
      .this_rdy(start_rdy),
      .this_dat(start_dat),
      .data_rsc_z(start_PopNB_mioi_data_rsc_z),
      .return_rsc_z(start_PopNB_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(start_PopNB_mioi_biwt_iff),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  ActUnit_ActUnit_ActUnitRun_start_PopNB_mioi_start_PopNB_mio_wait_ctrl ActUnit_ActUnitRun_start_PopNB_mioi_start_PopNB_mio_wait_ctrl_inst
      (
      .ActUnitRun_wen(ActUnitRun_wen),
      .ActUnitRun_wten(ActUnitRun_wten),
      .start_PopNB_mioi_oswt(start_PopNB_mioi_oswt),
      .start_PopNB_mioi_biwt(start_PopNB_mioi_biwt),
      .start_PopNB_mioi_bdwt(start_PopNB_mioi_bdwt),
      .start_PopNB_mioi_biwt_pff(start_PopNB_mioi_biwt_iff),
      .start_PopNB_mioi_oswt_pff(start_PopNB_mioi_oswt_pff)
    );
  ActUnit_ActUnit_ActUnitRun_start_PopNB_mioi_start_PopNB_mio_wait_dp ActUnit_ActUnitRun_start_PopNB_mioi_start_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .start_PopNB_mioi_data_rsc_z_mxwt(start_PopNB_mioi_data_rsc_z_mxwt),
      .start_PopNB_mioi_return_rsc_z_mxwt(start_PopNB_mioi_return_rsc_z_mxwt),
      .start_PopNB_mioi_biwt(start_PopNB_mioi_biwt),
      .start_PopNB_mioi_bdwt(start_PopNB_mioi_bdwt),
      .start_PopNB_mioi_data_rsc_z(start_PopNB_mioi_data_rsc_z),
      .start_PopNB_mioi_return_rsc_z(start_PopNB_mioi_return_rsc_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_rva_out_Push_mioi
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_rva_out_Push_mioi (
  clk, rst, rva_out_vld, rva_out_rdy, rva_out_dat, ActUnitRun_wten, rva_out_Push_mioi_oswt,
      rva_out_Push_mioi_wen_comp, rva_out_Push_mioi_m_data_rsc_dat_ActUnitRun, rva_out_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output rva_out_vld;
  input rva_out_rdy;
  output [511:0] rva_out_dat;
  input ActUnitRun_wten;
  input rva_out_Push_mioi_oswt;
  output rva_out_Push_mioi_wen_comp;
  input [511:0] rva_out_Push_mioi_m_data_rsc_dat_ActUnitRun;
  input rva_out_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire rva_out_Push_mioi_biwt;
  wire rva_out_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct;
  wire rva_out_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  ActUnit_Connections_OutBlocking_RVSink_spec_Axi_rvaCfg_Read_Connections_SYN_PORT_Push
      rva_out_Push_mioi (
      .this_vld(rva_out_vld),
      .this_rdy(rva_out_rdy),
      .this_dat(rva_out_dat),
      .m_data_rsc_dat(rva_out_Push_mioi_m_data_rsc_dat_ActUnitRun),
      .ccs_ccore_start_rsc_dat(rva_out_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct),
      .ccs_ccore_done_sync_vld(rva_out_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  ActUnit_ActUnit_ActUnitRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl ActUnit_ActUnitRun_rva_out_Push_mioi_rva_out_Push_mio_wait_ctrl_inst
      (
      .ActUnitRun_wten(ActUnitRun_wten),
      .rva_out_Push_mioi_iswt0(rva_out_Push_mioi_oswt),
      .rva_out_Push_mioi_biwt(rva_out_Push_mioi_biwt),
      .rva_out_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct(rva_out_Push_mioi_ccs_ccore_start_rsc_dat_ActUnitRun_sct),
      .rva_out_Push_mioi_ccs_ccore_done_sync_vld(rva_out_Push_mioi_ccs_ccore_done_sync_vld),
      .rva_out_Push_mioi_iswt0_pff(rva_out_Push_mioi_oswt_pff)
    );
  assign rva_out_Push_mioi_wen_comp = (~ rva_out_Push_mioi_oswt) | rva_out_Push_mioi_biwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_act_port_PopNB_mioi
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_act_port_PopNB_mioi (
  clk, rst, act_port_vld, act_port_rdy, act_port_dat, ActUnitRun_wen, ActUnitRun_wten,
      act_port_PopNB_mioi_oswt, act_port_PopNB_mioi_data_data_rsc_z_mxwt, act_port_PopNB_mioi_return_rsc_z_mxwt,
      act_port_PopNB_mioi_oswt_pff
);
  input clk;
  input rst;
  input act_port_vld;
  output act_port_rdy;
  input [511:0] act_port_dat;
  input ActUnitRun_wen;
  input ActUnitRun_wten;
  input act_port_PopNB_mioi_oswt;
  output [511:0] act_port_PopNB_mioi_data_data_rsc_z_mxwt;
  output act_port_PopNB_mioi_return_rsc_z_mxwt;
  input act_port_PopNB_mioi_oswt_pff;


  // Interconnect Declarations
  wire act_port_PopNB_mioi_biwt;
  wire act_port_PopNB_mioi_bdwt;
  wire [511:0] act_port_PopNB_mioi_data_data_rsc_z;
  wire act_port_PopNB_mioi_return_rsc_z;
  wire act_port_PopNB_mioi_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  ActUnit_Connections_InBlocking_spec_ActVectorType_Connections_SYN_PORT_PopNB  act_port_PopNB_mioi
      (
      .this_vld(act_port_vld),
      .this_rdy(act_port_rdy),
      .this_dat(act_port_dat),
      .data_data_rsc_z(act_port_PopNB_mioi_data_data_rsc_z),
      .return_rsc_z(act_port_PopNB_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(act_port_PopNB_mioi_biwt_iff),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  ActUnit_ActUnit_ActUnitRun_act_port_PopNB_mioi_act_port_PopNB_mio_wait_ctrl ActUnit_ActUnitRun_act_port_PopNB_mioi_act_port_PopNB_mio_wait_ctrl_inst
      (
      .ActUnitRun_wen(ActUnitRun_wen),
      .ActUnitRun_wten(ActUnitRun_wten),
      .act_port_PopNB_mioi_oswt(act_port_PopNB_mioi_oswt),
      .act_port_PopNB_mioi_biwt(act_port_PopNB_mioi_biwt),
      .act_port_PopNB_mioi_bdwt(act_port_PopNB_mioi_bdwt),
      .act_port_PopNB_mioi_biwt_pff(act_port_PopNB_mioi_biwt_iff),
      .act_port_PopNB_mioi_oswt_pff(act_port_PopNB_mioi_oswt_pff)
    );
  ActUnit_ActUnit_ActUnitRun_act_port_PopNB_mioi_act_port_PopNB_mio_wait_dp ActUnit_ActUnitRun_act_port_PopNB_mioi_act_port_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .act_port_PopNB_mioi_data_data_rsc_z_mxwt(act_port_PopNB_mioi_data_data_rsc_z_mxwt),
      .act_port_PopNB_mioi_return_rsc_z_mxwt(act_port_PopNB_mioi_return_rsc_z_mxwt),
      .act_port_PopNB_mioi_biwt(act_port_PopNB_mioi_biwt),
      .act_port_PopNB_mioi_bdwt(act_port_PopNB_mioi_bdwt),
      .act_port_PopNB_mioi_data_data_rsc_z(act_port_PopNB_mioi_data_data_rsc_z),
      .act_port_PopNB_mioi_return_rsc_z(act_port_PopNB_mioi_return_rsc_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun_rva_in_PopNB_mioi
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun_rva_in_PopNB_mioi (
  clk, rst, rva_in_vld, rva_in_rdy, rva_in_dat, ActUnitRun_wen, ActUnitRun_wten,
      rva_in_PopNB_mioi_oswt, rva_in_PopNB_mioi_data_data_rsc_z_mxwt, rva_in_PopNB_mioi_data_addr_rsc_z_mxwt,
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt, rva_in_PopNB_mioi_return_rsc_z_mxwt,
      rva_in_PopNB_mioi_oswt_pff
);
  input clk;
  input rst;
  input rva_in_vld;
  output rva_in_rdy;
  input [600:0] rva_in_dat;
  input ActUnitRun_wen;
  input ActUnitRun_wten;
  input rva_in_PopNB_mioi_oswt;
  output [511:0] rva_in_PopNB_mioi_data_data_rsc_z_mxwt;
  output [11:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt;
  output rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  output rva_in_PopNB_mioi_return_rsc_z_mxwt;
  input rva_in_PopNB_mioi_oswt_pff;


  // Interconnect Declarations
  wire rva_in_PopNB_mioi_biwt;
  wire rva_in_PopNB_mioi_bdwt;
  wire [511:0] rva_in_PopNB_mioi_data_data_rsc_z;
  wire [23:0] rva_in_PopNB_mioi_data_addr_rsc_z;
  wire rva_in_PopNB_mioi_data_rw_rsc_z;
  wire rva_in_PopNB_mioi_return_rsc_z;
  wire [11:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt_pconst;
  wire rva_in_PopNB_mioi_biwt_iff;


  // Interconnect Declarations for Component Instantiations 
  ActUnit_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB
      rva_in_PopNB_mioi (
      .this_vld(rva_in_vld),
      .this_rdy(rva_in_rdy),
      .this_dat(rva_in_dat),
      .data_data_rsc_z(rva_in_PopNB_mioi_data_data_rsc_z),
      .data_addr_rsc_z(rva_in_PopNB_mioi_data_addr_rsc_z),
      .data_rw_rsc_z(rva_in_PopNB_mioi_data_rw_rsc_z),
      .return_rsc_z(rva_in_PopNB_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(rva_in_PopNB_mioi_biwt_iff),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  ActUnit_ActUnit_ActUnitRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl ActUnit_ActUnitRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_ctrl_inst
      (
      .ActUnitRun_wen(ActUnitRun_wen),
      .ActUnitRun_wten(ActUnitRun_wten),
      .rva_in_PopNB_mioi_oswt(rva_in_PopNB_mioi_oswt),
      .rva_in_PopNB_mioi_biwt(rva_in_PopNB_mioi_biwt),
      .rva_in_PopNB_mioi_bdwt(rva_in_PopNB_mioi_bdwt),
      .rva_in_PopNB_mioi_biwt_pff(rva_in_PopNB_mioi_biwt_iff),
      .rva_in_PopNB_mioi_oswt_pff(rva_in_PopNB_mioi_oswt_pff)
    );
  ActUnit_ActUnit_ActUnitRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp ActUnit_ActUnitRun_rva_in_PopNB_mioi_rva_in_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_in_PopNB_mioi_data_data_rsc_z_mxwt(rva_in_PopNB_mioi_data_data_rsc_z_mxwt),
      .rva_in_PopNB_mioi_data_addr_rsc_z_mxwt(rva_in_PopNB_mioi_data_addr_rsc_z_mxwt_pconst),
      .rva_in_PopNB_mioi_data_rw_rsc_z_mxwt(rva_in_PopNB_mioi_data_rw_rsc_z_mxwt),
      .rva_in_PopNB_mioi_return_rsc_z_mxwt(rva_in_PopNB_mioi_return_rsc_z_mxwt),
      .rva_in_PopNB_mioi_biwt(rva_in_PopNB_mioi_biwt),
      .rva_in_PopNB_mioi_bdwt(rva_in_PopNB_mioi_bdwt),
      .rva_in_PopNB_mioi_data_data_rsc_z(rva_in_PopNB_mioi_data_data_rsc_z),
      .rva_in_PopNB_mioi_data_addr_rsc_z(rva_in_PopNB_mioi_data_addr_rsc_z),
      .rva_in_PopNB_mioi_data_rw_rsc_z(rva_in_PopNB_mioi_data_rw_rsc_z),
      .rva_in_PopNB_mioi_return_rsc_z(rva_in_PopNB_mioi_return_rsc_z)
    );
  assign rva_in_PopNB_mioi_data_addr_rsc_z_mxwt = rva_in_PopNB_mioi_data_addr_rsc_z_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit_ActUnit_ActUnitRun
// ------------------------------------------------------------------


module ActUnit_ActUnit_ActUnitRun (
  clk, rst, start_vld, start_rdy, start_dat, act_port_vld, act_port_rdy, act_port_dat,
      rva_in_vld, rva_in_rdy, rva_in_dat, rva_out_vld, rva_out_rdy, rva_out_dat,
      output_port_vld, output_port_rdy, output_port_dat, done_vld, done_rdy, done_dat
);
  input clk;
  input rst;
  input start_vld;
  output start_rdy;
  input start_dat;
  input act_port_vld;
  output act_port_rdy;
  input [511:0] act_port_dat;
  input rva_in_vld;
  output rva_in_rdy;
  input [600:0] rva_in_dat;
  output rva_out_vld;
  input rva_out_rdy;
  output [511:0] rva_out_dat;
  output output_port_vld;
  input output_port_rdy;
  output [521:0] output_port_dat;
  output done_vld;
  input done_rdy;
  output done_dat;


  // Interconnect Declarations
  wire ActUnitRun_wen;
  wire ActUnitRun_wten;
  wire [511:0] rva_in_PopNB_mioi_data_data_rsc_z_mxwt;
  wire [11:0] rva_in_PopNB_mioi_data_addr_rsc_z_mxwt;
  wire rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  wire rva_in_PopNB_mioi_return_rsc_z_mxwt;
  wire [511:0] act_port_PopNB_mioi_data_data_rsc_z_mxwt;
  wire act_port_PopNB_mioi_return_rsc_z_mxwt;
  wire rva_out_Push_mioi_wen_comp;
  wire start_PopNB_mioi_data_rsc_z_mxwt;
  wire start_PopNB_mioi_return_rsc_z_mxwt;
  wire output_port_Push_mioi_wen_comp;
  wire done_Push_mioi_wen_comp;
  wire Gelu_for_1_else_else_else_if_mul_cmp_en;
  wire [50:0] Gelu_for_1_else_else_else_if_mul_cmp_z;
  wire Gelu_for_1_else_else_else_if_mul_cmp_1_en;
  wire [50:0] Gelu_for_1_else_else_else_if_mul_cmp_1_z;
  wire Gelu_for_1_else_else_else_if_mul_cmp_2_en;
  wire [50:0] Gelu_for_1_else_else_else_if_mul_cmp_2_z;
  wire Gelu_for_1_else_else_else_if_mul_cmp_3_en;
  wire [50:0] Gelu_for_1_else_else_else_if_mul_cmp_3_z;
  wire Gelu_for_1_else_else_else_if_mul_cmp_4_en;
  wire [50:0] Gelu_for_1_else_else_else_if_mul_cmp_4_z;
  wire Gelu_for_1_else_else_else_if_mul_cmp_5_en;
  wire [50:0] Gelu_for_1_else_else_else_if_mul_cmp_5_z;
  wire Gelu_for_1_else_else_else_if_mul_cmp_6_en;
  wire [50:0] Gelu_for_1_else_else_else_if_mul_cmp_6_z;
  wire Gelu_for_1_else_else_else_if_mul_cmp_7_en;
  wire [50:0] Gelu_for_1_else_else_else_if_mul_cmp_7_z;
  wire Gelu_for_1_else_else_else_if_mul_cmp_8_en;
  wire [50:0] Gelu_for_1_else_else_else_if_mul_cmp_8_z;
  wire Gelu_for_1_else_else_else_if_mul_cmp_9_en;
  wire [50:0] Gelu_for_1_else_else_else_if_mul_cmp_9_z;
  wire Gelu_for_1_else_else_else_if_mul_cmp_10_en;
  wire [50:0] Gelu_for_1_else_else_else_if_mul_cmp_10_z;
  wire Gelu_for_1_else_else_else_if_mul_cmp_11_en;
  wire [50:0] Gelu_for_1_else_else_else_if_mul_cmp_11_z;
  wire Gelu_for_1_else_else_else_if_mul_cmp_12_en;
  wire [50:0] Gelu_for_1_else_else_else_if_mul_cmp_12_z;
  wire Gelu_for_1_else_else_else_if_mul_cmp_13_en;
  wire [50:0] Gelu_for_1_else_else_else_if_mul_cmp_13_z;
  wire Gelu_for_1_else_else_else_if_mul_cmp_14_en;
  wire [50:0] Gelu_for_1_else_else_else_if_mul_cmp_14_z;
  wire Gelu_for_1_else_else_else_if_mul_cmp_15_en;
  wire [50:0] Gelu_for_1_else_else_else_if_mul_cmp_15_z;
  wire Gelu_for_1_else_else_if_mul_cmp_en;
  wire [46:0] Gelu_for_1_else_else_if_mul_cmp_z;
  wire Gelu_for_1_else_else_if_mul_cmp_1_en;
  wire [46:0] Gelu_for_1_else_else_if_mul_cmp_1_z;
  wire Gelu_for_1_else_else_if_mul_cmp_2_en;
  wire [46:0] Gelu_for_1_else_else_if_mul_cmp_2_z;
  wire Gelu_for_1_else_else_if_mul_cmp_3_en;
  wire [46:0] Gelu_for_1_else_else_if_mul_cmp_3_z;
  wire Gelu_for_1_else_else_if_mul_cmp_4_en;
  wire [46:0] Gelu_for_1_else_else_if_mul_cmp_4_z;
  wire Gelu_for_1_else_else_if_mul_cmp_5_en;
  wire [46:0] Gelu_for_1_else_else_if_mul_cmp_5_z;
  wire Gelu_for_1_else_else_if_mul_cmp_6_en;
  wire [46:0] Gelu_for_1_else_else_if_mul_cmp_6_z;
  wire Gelu_for_1_else_else_if_mul_cmp_7_en;
  wire [46:0] Gelu_for_1_else_else_if_mul_cmp_7_z;
  wire Gelu_for_1_else_else_if_mul_cmp_8_en;
  wire [46:0] Gelu_for_1_else_else_if_mul_cmp_8_z;
  wire Gelu_for_1_else_else_if_mul_cmp_9_en;
  wire [46:0] Gelu_for_1_else_else_if_mul_cmp_9_z;
  wire Gelu_for_1_else_else_if_mul_cmp_10_en;
  wire [46:0] Gelu_for_1_else_else_if_mul_cmp_10_z;
  wire Gelu_for_1_else_else_if_mul_cmp_11_en;
  wire [46:0] Gelu_for_1_else_else_if_mul_cmp_11_z;
  wire Gelu_for_1_else_else_if_mul_cmp_12_en;
  wire [46:0] Gelu_for_1_else_else_if_mul_cmp_12_z;
  wire Gelu_for_1_else_else_if_mul_cmp_13_en;
  wire [46:0] Gelu_for_1_else_else_if_mul_cmp_13_z;
  wire Gelu_for_1_else_else_if_mul_cmp_14_en;
  wire [46:0] Gelu_for_1_else_else_if_mul_cmp_14_z;
  wire Gelu_for_1_else_else_if_mul_cmp_15_en;
  wire [46:0] Gelu_for_1_else_else_if_mul_cmp_15_z;
  wire Silu_for_1_else_if_Silu_for_else_if_mul_cmp_en;
  wire [47:0] Silu_for_1_else_if_Silu_for_else_if_mul_cmp_z;
  wire Silu_for_1_else_if_Silu_for_else_if_mul_cmp_1_en;
  wire [47:0] Silu_for_1_else_if_Silu_for_else_if_mul_cmp_1_z;
  wire Silu_for_1_else_if_Silu_for_else_if_mul_cmp_2_en;
  wire [47:0] Silu_for_1_else_if_Silu_for_else_if_mul_cmp_2_z;
  wire Silu_for_1_else_if_Silu_for_else_if_mul_cmp_3_en;
  wire [47:0] Silu_for_1_else_if_Silu_for_else_if_mul_cmp_3_z;
  wire Silu_for_1_else_if_Silu_for_else_if_mul_cmp_4_en;
  wire [47:0] Silu_for_1_else_if_Silu_for_else_if_mul_cmp_4_z;
  wire Silu_for_1_else_if_Silu_for_else_if_mul_cmp_5_en;
  wire [47:0] Silu_for_1_else_if_Silu_for_else_if_mul_cmp_5_z;
  wire Silu_for_1_else_if_Silu_for_else_if_mul_cmp_6_en;
  wire [47:0] Silu_for_1_else_if_Silu_for_else_if_mul_cmp_6_z;
  wire Silu_for_1_else_if_Silu_for_else_if_mul_cmp_7_en;
  wire [47:0] Silu_for_1_else_if_Silu_for_else_if_mul_cmp_7_z;
  wire [3:0] fsm_output;
  wire act_config_InstIncr_if_act_config_InstIncr_if_if_nor_tmp;
  wire act_config_InstIncr_if_equal_1_tmp;
  wire [6:0] operator_6_false_acc_tmp;
  wire [7:0] nl_operator_6_false_acc_tmp;
  wire Silu_for_else_and_19_tmp;
  wire Gelu_for_else_and_31_tmp;
  wire Gelu_for_else_and_29_tmp;
  wire Gelu_for_else_and_27_tmp;
  wire Gelu_for_else_and_25_tmp;
  wire Gelu_for_else_and_23_tmp;
  wire Gelu_for_else_and_21_tmp;
  wire Gelu_for_else_and_19_tmp;
  wire Gelu_for_else_and_17_tmp;
  wire Gelu_for_else_and_15_tmp;
  wire Gelu_for_else_and_13_tmp;
  wire Gelu_for_else_and_11_tmp;
  wire Gelu_for_else_and_9_tmp;
  wire Gelu_for_else_and_7_tmp;
  wire Gelu_for_else_and_5_tmp;
  wire Gelu_for_else_and_3_tmp;
  wire Gelu_for_else_and_1_tmp;
  wire Silu_for_else_and_15_tmp;
  wire Silu_for_else_and_13_tmp;
  wire Silu_for_else_and_11_tmp;
  wire Silu_for_else_and_9_tmp;
  wire Silu_for_else_and_7_tmp;
  wire Silu_for_else_and_5_tmp;
  wire Silu_for_else_and_3_tmp;
  wire Silu_for_else_and_1_tmp;
  wire ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_2_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_3_less_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_3_less_1_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_3_less_2_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_3_less_3_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_3_less_4_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_3_less_5_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_3_less_6_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_3_less_7_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_3_less_8_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_3_less_9_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_3_less_10_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_3_less_11_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_3_less_12_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_3_less_13_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_3_less_14_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_3_less_15_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_7_less_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_6_less_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_7_less_1_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_6_less_1_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_7_less_2_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_6_less_2_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_7_less_3_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_6_less_3_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_7_less_4_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_6_less_4_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_7_less_5_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_6_less_5_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_7_less_6_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_6_less_6_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_7_less_7_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_6_less_7_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_7_less_8_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_6_less_8_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_7_less_9_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_6_less_9_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_7_less_10_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_6_less_10_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_7_less_11_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_6_less_11_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_7_less_12_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_6_less_12_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_7_less_13_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_6_less_13_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_7_less_14_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_6_less_14_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_7_less_15_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_6_less_15_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_less_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_less_1_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_less_2_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_less_3_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_less_4_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_less_5_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_less_6_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_less_7_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_1_less_8_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_less_8_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_1_less_9_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_less_9_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_1_less_10_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_less_10_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_1_less_11_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_less_11_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_1_less_12_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_less_12_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_1_less_13_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_less_13_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_1_less_14_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_less_14_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_1_less_15_tmp;
  wire operator_32_8_true_AC_TRN_AC_WRAP_less_15_tmp;
  wire Gelu_for_if_less_tmp;
  wire Gelu_for_if_less_1_tmp;
  wire Gelu_for_if_less_2_tmp;
  wire Gelu_for_if_less_3_tmp;
  wire Gelu_for_if_less_4_tmp;
  wire Gelu_for_if_less_5_tmp;
  wire Gelu_for_if_less_6_tmp;
  wire Gelu_for_if_less_7_tmp;
  wire Gelu_for_else_if_less_8_tmp;
  wire Gelu_for_if_less_8_tmp;
  wire Gelu_for_else_if_less_9_tmp;
  wire Gelu_for_if_less_9_tmp;
  wire Gelu_for_else_if_less_10_tmp;
  wire Gelu_for_if_less_10_tmp;
  wire Gelu_for_else_if_less_11_tmp;
  wire Gelu_for_if_less_11_tmp;
  wire Gelu_for_else_if_less_12_tmp;
  wire Gelu_for_if_less_12_tmp;
  wire Gelu_for_else_if_less_13_tmp;
  wire Gelu_for_if_less_13_tmp;
  wire Gelu_for_else_if_less_14_tmp;
  wire Gelu_for_if_less_14_tmp;
  wire Gelu_for_else_if_less_15_tmp;
  wire Gelu_for_if_less_15_tmp;
  wire [7:0] act_config_in_InstFetch_mux_tmp;
  wire [4:0] while_mux_55_tmp;
  wire while_and_1_tmp;
  wire and_dcpl_7;
  wire and_dcpl_9;
  wire and_dcpl_40;
  wire and_dcpl_43;
  wire or_tmp;
  wire or_dcpl_28;
  wire and_dcpl_78;
  wire and_dcpl_83;
  wire and_dcpl_84;
  wire and_dcpl_86;
  wire and_dcpl_117;
  wire and_dcpl_331;
  wire and_dcpl_332;
  wire and_dcpl_333;
  wire or_tmp_146;
  wire not_tmp_237;
  wire and_dcpl_337;
  wire or_tmp_158;
  wire mux_tmp_108;
  wire and_dcpl_469;
  wire or_tmp_397;
  wire or_dcpl_450;
  wire and_dcpl_846;
  wire and_dcpl_847;
  wire and_dcpl_848;
  wire and_dcpl_849;
  wire and_dcpl_852;
  wire and_dcpl_855;
  wire or_dcpl_457;
  wire and_dcpl_856;
  wire or_tmp_409;
  wire mux_tmp_315;
  wire mux_tmp_317;
  wire mux_tmp_318;
  wire nand_tmp_23;
  wire mux_tmp_325;
  wire mux_tmp_327;
  wire mux_tmp_328;
  wire nand_tmp_25;
  wire mux_tmp_335;
  wire mux_tmp_337;
  wire mux_tmp_338;
  wire nand_tmp_27;
  wire mux_tmp_345;
  wire mux_tmp_347;
  wire mux_tmp_348;
  wire nand_tmp_29;
  wire mux_tmp_355;
  wire mux_tmp_357;
  wire mux_tmp_358;
  wire nand_tmp_31;
  wire mux_tmp_365;
  wire mux_tmp_367;
  wire mux_tmp_368;
  wire nand_tmp_33;
  wire mux_tmp_375;
  wire mux_tmp_377;
  wire mux_tmp_378;
  wire nand_tmp_35;
  wire mux_tmp_385;
  wire mux_tmp_387;
  wire mux_tmp_388;
  wire nand_tmp_37;
  wire and_dcpl_867;
  wire not_tmp_445;
  wire and_dcpl_872;
  wire and_dcpl_953;
  wire and_dcpl_1048;
  wire and_dcpl_1051;
  wire and_dcpl_1056;
  wire and_dcpl_1061;
  wire and_dcpl_1062;
  wire and_dcpl_1063;
  wire and_dcpl_1072;
  wire and_dcpl_1077;
  wire and_dcpl_1081;
  wire and_dcpl_1082;
  wire and_dcpl_1083;
  wire and_dcpl_1085;
  wire or_dcpl_462;
  wire or_dcpl_464;
  wire or_dcpl_465;
  wire and_dcpl_1088;
  wire or_dcpl_466;
  wire or_dcpl_468;
  wire or_dcpl_469;
  wire and_dcpl_1090;
  wire or_dcpl_475;
  wire or_dcpl_485;
  wire or_dcpl_487;
  wire or_tmp_484;
  wire mux_tmp_413;
  wire and_dcpl_1093;
  wire and_dcpl_1094;
  wire and_dcpl_1096;
  wire or_tmp_485;
  wire not_tmp_495;
  wire or_dcpl_492;
  wire or_dcpl_493;
  wire or_dcpl_494;
  wire or_dcpl_496;
  wire or_dcpl_498;
  wire or_dcpl_500;
  wire or_dcpl_501;
  wire or_dcpl_504;
  wire or_dcpl_505;
  wire or_dcpl_508;
  wire or_dcpl_509;
  wire or_dcpl_512;
  wire or_dcpl_513;
  wire or_dcpl_516;
  wire or_dcpl_519;
  wire or_dcpl_522;
  wire or_dcpl_525;
  wire or_dcpl_526;
  wire or_dcpl_529;
  wire or_dcpl_532;
  wire or_dcpl_535;
  wire or_dcpl_538;
  wire or_dcpl_539;
  wire or_dcpl_542;
  wire or_dcpl_545;
  wire or_dcpl_548;
  wire or_dcpl_552;
  wire not_tmp_503;
  wire or_dcpl_586;
  wire and_dcpl_1104;
  wire and_dcpl_1106;
  wire and_dcpl_1109;
  wire and_dcpl_1112;
  wire or_dcpl_593;
  wire or_dcpl_595;
  wire or_dcpl_596;
  wire or_dcpl_616;
  wire or_dcpl_622;
  wire or_dcpl_623;
  wire and_dcpl_1116;
  wire and_dcpl_1118;
  wire or_dcpl_717;
  wire and_dcpl_1143;
  wire and_dcpl_1144;
  wire and_dcpl_1174;
  wire and_dcpl_1228;
  wire and_dcpl_1233;
  wire and_dcpl_1235;
  wire and_dcpl_1236;
  wire or_dcpl_815;
  wire or_dcpl_817;
  wire or_dcpl_822;
  wire or_dcpl_823;
  wire and_dcpl_1240;
  wire or_dcpl_824;
  wire or_dcpl_825;
  wire or_dcpl_826;
  wire or_dcpl_827;
  wire or_dcpl_828;
  wire or_dcpl_829;
  wire or_dcpl_830;
  wire or_dcpl_831;
  wire or_dcpl_833;
  wire or_dcpl_835;
  wire or_dcpl_836;
  wire or_dcpl_837;
  wire or_dcpl_838;
  wire or_dcpl_839;
  wire or_dcpl_840;
  wire or_dcpl_841;
  wire or_dcpl_842;
  wire or_dcpl_843;
  wire and_dcpl_1244;
  wire and_dcpl_1246;
  wire and_dcpl_1257;
  wire and_dcpl_1262;
  wire mux_tmp_433;
  wire or_dcpl_846;
  wire or_dcpl_847;
  wire or_dcpl_848;
  wire or_dcpl_849;
  wire or_dcpl_850;
  wire or_dcpl_851;
  wire or_dcpl_852;
  wire or_dcpl_853;
  wire or_dcpl_854;
  wire or_dcpl_855;
  wire or_dcpl_856;
  wire or_dcpl_857;
  wire or_dcpl_858;
  wire or_dcpl_859;
  wire or_dcpl_860;
  wire or_dcpl_861;
  wire or_dcpl_862;
  wire or_dcpl_863;
  wire or_dcpl_864;
  wire or_dcpl_865;
  wire or_dcpl_866;
  wire or_dcpl_867;
  wire or_dcpl_868;
  wire or_dcpl_869;
  wire or_dcpl_870;
  wire or_dcpl_871;
  wire or_dcpl_872;
  wire or_dcpl_873;
  wire or_dcpl_874;
  wire or_dcpl_875;
  wire or_tmp_490;
  wire and_dcpl_1264;
  wire and_dcpl_1265;
  wire and_dcpl_1266;
  wire and_dcpl_1267;
  wire and_dcpl_1270;
  wire and_dcpl_1271;
  wire and_dcpl_1272;
  wire and_dcpl_1274;
  wire and_dcpl_1275;
  wire or_dcpl_877;
  wire or_dcpl_878;
  wire and_dcpl_1277;
  wire and_dcpl_1278;
  wire and_dcpl_1280;
  wire and_dcpl_1281;
  wire and_dcpl_1282;
  wire and_dcpl_1284;
  wire and_dcpl_1285;
  wire and_dcpl_1287;
  wire and_dcpl_1288;
  wire and_dcpl_1289;
  wire and_dcpl_1291;
  wire and_dcpl_1292;
  wire and_dcpl_1294;
  wire and_dcpl_1295;
  wire and_dcpl_1297;
  wire and_dcpl_1299;
  wire and_dcpl_1300;
  wire or_dcpl_887;
  wire and_dcpl_1302;
  wire and_dcpl_1304;
  wire and_dcpl_1306;
  wire and_dcpl_1308;
  wire and_dcpl_1310;
  wire and_dcpl_1312;
  wire and_dcpl_1314;
  wire and_dcpl_1316;
  wire and_dcpl_1317;
  wire and_dcpl_1318;
  wire or_dcpl_896;
  wire or_dcpl_897;
  wire and_dcpl_1320;
  wire and_dcpl_1322;
  wire and_dcpl_1324;
  wire and_dcpl_1326;
  wire and_dcpl_1328;
  wire and_dcpl_1330;
  wire and_dcpl_1332;
  wire and_dcpl_1334;
  wire and_dcpl_1335;
  wire and_dcpl_1336;
  wire or_dcpl_906;
  wire and_dcpl_1338;
  wire and_dcpl_1340;
  wire and_dcpl_1342;
  wire and_dcpl_1344;
  wire and_dcpl_1346;
  wire and_dcpl_1348;
  wire and_dcpl_1350;
  wire and_dcpl_1352;
  wire and_dcpl_1353;
  wire or_dcpl_915;
  wire or_dcpl_916;
  wire and_dcpl_1355;
  wire and_dcpl_1357;
  wire and_dcpl_1359;
  wire and_dcpl_1361;
  wire and_dcpl_1363;
  wire and_dcpl_1365;
  wire and_dcpl_1367;
  wire and_dcpl_1369;
  wire and_dcpl_1370;
  wire or_dcpl_925;
  wire and_dcpl_1372;
  wire and_dcpl_1374;
  wire and_dcpl_1376;
  wire and_dcpl_1378;
  wire and_dcpl_1380;
  wire and_dcpl_1382;
  wire and_dcpl_1384;
  wire and_dcpl_1386;
  wire not_tmp_620;
  wire and_dcpl_1388;
  wire and_dcpl_1390;
  wire and_dcpl_1391;
  wire and_dcpl_1393;
  wire and_dcpl_1395;
  wire and_dcpl_1396;
  wire and_dcpl_1402;
  wire not_tmp_640;
  wire or_dcpl_934;
  wire or_dcpl_936;
  wire or_dcpl_945;
  wire or_dcpl_946;
  wire or_dcpl_955;
  wire or_dcpl_956;
  wire or_dcpl_965;
  wire or_dcpl_974;
  wire or_dcpl_975;
  wire or_dcpl_984;
  wire or_dcpl_985;
  wire or_dcpl_994;
  wire or_dcpl_1003;
  wire act_config_InstIncr_act_config_InstIncr_if_and_svs_1;
  wire [8:0] operator_8_false_acc_sdt_sva_1;
  wire [9:0] nl_operator_8_false_acc_sdt_sva_1;
  reg ActUnit_PushOutput_if_for_and_stg_2_7_sva;
  reg Gelu_for_and_2_cse_sva;
  reg ActUnit_RunInst_switch_lp_equal_tmp_8;
  reg is_start_sva;
  reg ActUnit_RunInst_switch_lp_equal_tmp_7;
  reg ActUnit_RunInst_switch_lp_equal_tmp_6;
  reg ActUnit_RunInst_switch_lp_equal_tmp_5;
  reg ActUnit_RunInst_switch_lp_equal_tmp_4;
  reg ActUnit_CheckStart_start_reg_sva;
  reg ActUnit_RunInst_switch_lp_equal_tmp_2;
  reg while_nor_48_itm;
  reg ActUnit_RunInst_switch_lp_and_32_tmp;
  reg while_nor_32_itm;
  reg ActUnit_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva;
  reg while_nor_16_itm;
  reg ActUnit_RunInst_switch_lp_and_tmp;
  reg while_nor_itm;
  reg Gelu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs;
  reg Gelu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs;
  wire Silu_for_else_and_31_m1c_mx1;
  reg Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs;
  reg Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  reg Gelu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs;
  reg Gelu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs;
  wire Silu_for_else_and_29_m1c_mx1;
  reg Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs;
  reg Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  reg Gelu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs;
  reg Gelu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs;
  wire Silu_for_else_and_27_m1c_mx1;
  reg Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs;
  reg Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  reg Gelu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs;
  reg Gelu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs;
  wire Silu_for_else_and_25_m1c_mx1;
  reg Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs;
  reg Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  reg Gelu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs;
  reg Gelu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs;
  wire Silu_for_else_and_23_m1c_mx1;
  reg Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs;
  reg Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  reg Gelu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs;
  reg Gelu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs;
  wire Silu_for_else_and_21_m1c_mx1;
  reg Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs;
  reg Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  reg Gelu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs;
  reg Gelu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs;
  wire Silu_for_else_and_19_m1c_mx1;
  reg Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs;
  reg Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  reg Gelu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs;
  reg Gelu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs;
  wire Silu_for_else_and_17_m1c_mx1;
  reg Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs;
  reg Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  wire Gelu_for_else_and_31_m1c_mx1;
  reg Gelu_for_16_else_slc_32_svs;
  wire Gelu_for_else_and_29_m1c_mx1;
  reg Gelu_for_15_else_slc_32_svs;
  wire Gelu_for_else_and_27_m1c_mx1;
  reg Gelu_for_14_else_slc_32_svs;
  wire Gelu_for_else_and_25_m1c_mx1;
  reg Gelu_for_13_else_slc_32_svs;
  wire Gelu_for_else_and_23_m1c_mx1;
  reg Gelu_for_12_else_slc_32_svs;
  wire Gelu_for_else_and_21_m1c_mx1;
  reg Gelu_for_11_else_slc_32_svs;
  wire Gelu_for_else_and_19_m1c_mx1;
  reg Gelu_for_10_else_slc_32_svs;
  wire Gelu_for_else_and_17_m1c_mx1;
  reg Gelu_for_9_else_slc_32_svs;
  reg Gelu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs;
  reg Gelu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs;
  wire Gelu_for_else_and_15_m1c_mx1;
  reg Gelu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs;
  reg Gelu_for_8_else_slc_32_svs;
  reg Gelu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs;
  reg Gelu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs;
  wire Gelu_for_else_and_13_m1c_mx1;
  reg Gelu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs;
  reg Gelu_for_7_else_slc_32_svs;
  reg Gelu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs;
  reg Gelu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs;
  wire Gelu_for_else_and_11_m1c_mx1;
  reg Gelu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs;
  reg Gelu_for_6_else_slc_32_svs;
  reg Gelu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs;
  reg Gelu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs;
  wire Gelu_for_else_and_9_m1c_mx1;
  reg Gelu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs;
  reg Gelu_for_5_else_slc_32_svs;
  reg Gelu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs;
  reg Gelu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs;
  wire Gelu_for_else_and_7_m1c_mx1;
  reg Gelu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs;
  reg Gelu_for_4_else_slc_32_svs;
  reg Gelu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs;
  reg Gelu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs;
  wire Gelu_for_else_and_5_m1c_mx1;
  reg Gelu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs;
  reg Gelu_for_3_else_slc_32_svs;
  reg Gelu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs;
  reg Gelu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs;
  wire Gelu_for_else_and_3_m1c_mx1;
  reg Gelu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs;
  reg Gelu_for_2_else_slc_32_svs;
  reg Gelu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs;
  reg Gelu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs;
  wire Gelu_for_else_and_1_m1c_mx1;
  reg Gelu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs;
  reg Gelu_for_1_else_slc_32_svs;
  wire Silu_for_else_and_15_m1c_mx1;
  reg Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs;
  reg Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  wire Silu_for_else_and_13_m1c_mx1;
  reg Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs;
  reg Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  wire Silu_for_else_and_11_m1c_mx1;
  reg Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs;
  reg Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  wire Silu_for_else_and_9_m1c_mx1;
  reg Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs;
  reg Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  wire Silu_for_else_and_7_m1c_mx1;
  reg Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs;
  reg Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  wire Silu_for_else_and_5_m1c_mx1;
  reg Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs;
  reg Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  wire Silu_for_else_and_3_m1c_mx1;
  reg Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs;
  reg Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  wire Silu_for_else_and_1_m1c_mx1;
  reg Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs;
  reg Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  wire act_config_ActConfigRead_unequal_tmp_1;
  wire ActUnit_DecodeAxi_if_or_7_tmp_1;
  wire while_and_88_tmp_1;
  wire ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_mx1;
  wire ActUnit_DecodeAxi_rva_in_reg_rw_sva_mx1;
  wire act_config_ActConfigRead_else_unequal_tmp_1;
  wire ActUnit_DecodeAxiRead_unequal_tmp_1;
  wire Tanh_for_nor_cse_sva_mx0w0;
  wire ActUnit_RunInst_switch_lp_nor_tmp_mx0;
  wire Tanh_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
  wire Tanh_for_15_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
  wire Tanh_for_14_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
  wire Tanh_for_13_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
  wire Tanh_for_12_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
  wire Tanh_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
  wire Tanh_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
  wire Tanh_for_9_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
  wire Tanh_for_8_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
  wire Tanh_for_7_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
  wire Tanh_for_6_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
  wire Tanh_for_5_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
  wire Tanh_for_4_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
  wire Tanh_for_3_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
  wire Tanh_for_2_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
  wire Tanh_for_1_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
  reg act_config_is_zero_first_sva_dfm_4;
  reg w_load_lpi_1_dfm_1;
  reg is_incr_lpi_1_dfm_1;
  reg act_config_is_valid_sva;
  reg [7:0] act_config_inst_regs_16_sva_dfm_6;
  reg [7:0] act_config_inst_regs_17_sva_dfm_6;
  reg [7:0] act_config_inst_regs_18_sva_dfm_6;
  reg [7:0] act_config_inst_regs_19_sva_dfm_6;
  reg [7:0] act_config_inst_regs_20_sva_dfm_6;
  reg [7:0] act_config_inst_regs_21_sva_dfm_6;
  reg [7:0] act_config_inst_regs_22_sva_dfm_6;
  reg [7:0] act_config_inst_regs_23_sva_dfm_6;
  reg [7:0] act_config_inst_regs_24_sva_dfm_6;
  reg [7:0] act_config_inst_regs_25_sva_dfm_6;
  reg [7:0] act_config_inst_regs_26_sva_dfm_6;
  reg [7:0] act_config_inst_regs_27_sva_dfm_6;
  reg [7:0] act_config_inst_regs_28_sva_dfm_6;
  reg [7:0] act_config_inst_regs_29_sva_dfm_6;
  reg [7:0] act_config_inst_regs_30_sva_dfm_6;
  reg [7:0] act_config_inst_regs_31_sva_dfm_6;
  reg [4:0] act_config_inst_counter_sva_dfm_3;
  wire [7:0] ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_23_4_mx1_tmp_7_0;
  reg Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  reg [5:0] act_config_in_InstFetch_return_sva_7_2;
  reg Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  reg Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  reg Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  reg Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  reg Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  reg Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  reg Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  reg Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  reg act_config_is_zero_first_sva;
  reg Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  reg Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  reg Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  reg Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  reg Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  reg Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  reg Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  reg Gelu_for_1_slc_32_1_svs;
  reg Gelu_for_2_slc_32_1_svs;
  reg Gelu_for_3_slc_32_1_svs;
  reg Gelu_for_4_slc_32_1_svs;
  reg Gelu_for_5_slc_32_1_svs;
  reg Gelu_for_6_slc_32_1_svs;
  reg Gelu_for_7_slc_32_1_svs;
  reg Gelu_for_8_slc_32_1_svs;
  reg Gelu_for_9_slc_32_1_svs;
  reg Gelu_for_10_slc_32_1_svs;
  reg Gelu_for_11_slc_32_1_svs;
  reg Gelu_for_12_slc_32_1_svs;
  reg Gelu_for_13_slc_32_1_svs;
  reg Gelu_for_14_slc_32_1_svs;
  reg Gelu_for_15_slc_32_1_svs;
  reg Gelu_for_16_slc_32_1_svs;
  reg ActUnit_RunInst_switch_lp_equal_tmp_3;
  reg [3:0] ActUnit_PushOutput_if_for_i_4_0_sva_3_0;
  reg w_axi_rsp_lpi_1_dfm_1;
  reg act_read_req_valid_lpi_1_dfm_6;
  reg [1:0] nvhls_get_slc_2U_NVUINT8_return_3_sva;
  reg while_asn_262_itm;
  reg act_write_req_valid_lpi_1_dfm_5;
  wire ActUnit_RunInst_switch_lp_equal_tmp_1_mx0w0;
  wire ActUnit_RunInst_switch_lp_equal_tmp_2_mx0w0;
  wire ActUnit_RunInst_switch_lp_equal_tmp_3_mx0w0;
  wire ActUnit_RunInst_switch_lp_equal_tmp_4_mx0w0;
  wire ActUnit_RunInst_switch_lp_equal_tmp_5_mx0w0;
  wire ActUnit_RunInst_switch_lp_equal_tmp_6_mx0w0;
  wire ActUnit_RunInst_switch_lp_equal_tmp_7_mx0w0;
  wire ActUnit_RunInst_switch_lp_equal_tmp_8_mx0w0;
  wire [1:0] nvhls_get_slc_2U_NVUINT8_return_3_sva_1;
  reg [7:0] act_config_inst_regs_0_sva_dfm_5;
  reg [7:0] act_config_inst_regs_1_sva_dfm_5;
  reg [7:0] act_config_inst_regs_2_sva_dfm_5;
  reg [7:0] act_config_inst_regs_3_sva_dfm_5;
  reg [7:0] act_config_inst_regs_4_sva_dfm_5;
  reg [7:0] act_config_inst_regs_5_sva_dfm_5;
  reg [7:0] act_config_inst_regs_6_sva_dfm_5;
  reg [7:0] act_config_inst_regs_7_sva_dfm_5;
  reg [7:0] act_config_inst_regs_8_sva_dfm_5;
  reg [7:0] act_config_inst_regs_9_sva_dfm_5;
  reg [7:0] act_config_inst_regs_10_sva_dfm_5;
  reg [7:0] act_config_inst_regs_11_sva_dfm_5;
  reg [7:0] act_config_inst_regs_12_sva_dfm_5;
  reg [7:0] act_config_inst_regs_13_sva_dfm_5;
  reg [7:0] act_config_inst_regs_14_sva_dfm_5;
  reg [7:0] act_config_inst_regs_15_sva_dfm_5;
  reg [7:0] reg_ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_23_4_ftd_12;
  reg [2:0] reg_Silu_for_16_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd;
  reg [21:0] reg_Silu_for_16_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1;
  reg [2:0] reg_Silu_for_15_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd;
  reg [21:0] reg_Silu_for_15_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1;
  reg [2:0] reg_Silu_for_14_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd;
  reg [21:0] reg_Silu_for_14_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1;
  reg [2:0] reg_Silu_for_13_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd;
  reg [21:0] reg_Silu_for_13_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1;
  wire Silu_for_else_else_else_if_and_3_ssc;
  reg [2:0] reg_Silu_for_12_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd;
  reg [21:0] reg_Silu_for_12_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1;
  wire Silu_for_else_else_else_if_and_2_ssc;
  reg [2:0] reg_Silu_for_11_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd;
  reg [21:0] reg_Silu_for_11_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1;
  wire Silu_for_else_else_else_if_and_1_ssc;
  reg [2:0] reg_Silu_for_10_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd;
  reg [21:0] reg_Silu_for_10_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1;
  reg reg_act_regs_data_0_13_ftd;
  reg [4:0] reg_act_regs_data_0_13_ftd_1;
  reg [21:0] reg_act_regs_data_0_13_ftd_3;
  reg reg_act_regs_data_0_12_ftd;
  reg [4:0] reg_act_regs_data_0_12_ftd_1;
  reg [21:0] reg_act_regs_data_0_12_ftd_3;
  reg reg_act_regs_data_0_11_ftd;
  reg [4:0] reg_act_regs_data_0_11_ftd_1;
  reg [21:0] reg_act_regs_data_0_11_ftd_3;
  reg reg_act_regs_data_0_10_ftd;
  reg [4:0] reg_act_regs_data_0_10_ftd_1;
  reg [21:0] reg_act_regs_data_0_10_ftd_3;
  reg reg_act_regs_data_0_1_ftd;
  reg [4:0] reg_act_regs_data_0_1_ftd_1;
  reg [21:0] reg_act_regs_data_0_1_ftd_3;
  reg reg_act_regs_data_0_0_ftd;
  reg [4:0] reg_act_regs_data_0_0_ftd_1;
  reg [21:0] reg_act_regs_data_0_0_ftd_3;
  wire [7:0] operator_8_false_acc_sdt;
  wire [8:0] nl_operator_8_false_acc_sdt;
  wire act_config_output_counter_and_ssc;
  wire act_regs_data_and_ssc;
  wire rva_out_reg_data_and_ssc;
  wire act_mem_banks_write_if_for_if_mux_cse;
  wire act_mem_banks_write_if_for_if_mux_1_cse;
  wire act_mem_banks_read_for_mux_cse;
  wire act_mem_banks_read_for_mux_1_cse;
  reg reg_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_7_cse;
  reg reg_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_6_cse;
  reg reg_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_5_cse;
  reg reg_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_4_cse;
  reg reg_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_3_cse;
  reg reg_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_2_cse;
  reg reg_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_1_cse;
  reg reg_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_cse;
  reg reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_15_cse;
  reg reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_14_cse;
  reg reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_13_cse;
  reg reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_12_cse;
  reg reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_11_cse;
  reg reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_10_cse;
  reg reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_9_cse;
  reg reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_8_cse;
  reg reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_7_cse;
  reg reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_6_cse;
  reg reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_5_cse;
  reg reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_4_cse;
  reg reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_3_cse;
  reg reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_2_cse;
  reg reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_1_cse;
  reg reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_cse;
  reg reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_15_cse;
  reg reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_14_cse;
  reg reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_13_cse;
  reg reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_12_cse;
  reg reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_11_cse;
  reg reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_10_cse;
  reg reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_9_cse;
  reg reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_8_cse;
  reg reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_7_cse;
  reg reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_6_cse;
  reg reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_5_cse;
  reg reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_4_cse;
  reg reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_3_cse;
  reg reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_2_cse;
  reg reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_1_cse;
  reg reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_cse;
  reg reg_done_Push_mioi_iswt0_cse;
  reg reg_output_port_Push_mioi_iswt0_cse;
  reg reg_start_PopNB_mioi_iswt0_cse;
  reg reg_rva_out_Push_mioi_iswt0_cse;
  reg reg_act_port_PopNB_mioi_iswt0_cse;
  reg reg_rva_in_PopNB_mioi_iswt0_cse;
  wire act_config_num_inst_and_cse;
  wire act_mem_banks_bank_a_and_cse;
  wire act_mem_banks_bank_a_and_1_cse;
  wire act_mem_banks_bank_a_and_2_cse;
  wire act_mem_banks_bank_a_and_3_cse;
  wire act_mem_banks_bank_a_and_4_cse;
  wire act_mem_banks_bank_a_and_5_cse;
  wire act_mem_banks_bank_a_and_6_cse;
  wire act_mem_banks_bank_a_and_7_cse;
  wire act_mem_banks_bank_a_and_8_cse;
  wire act_mem_banks_bank_a_and_9_cse;
  wire act_mem_banks_bank_a_and_10_cse;
  wire act_mem_banks_bank_a_and_11_cse;
  wire act_mem_banks_bank_a_and_12_cse;
  wire act_mem_banks_bank_a_and_13_cse;
  wire act_mem_banks_bank_a_and_14_cse;
  wire act_mem_banks_bank_a_and_15_cse;
  wire act_mem_banks_bank_a_and_16_cse;
  wire act_mem_banks_bank_a_and_17_cse;
  wire act_mem_banks_bank_a_and_18_cse;
  wire act_mem_banks_bank_a_and_19_cse;
  wire act_mem_banks_bank_a_and_20_cse;
  wire act_mem_banks_bank_a_and_21_cse;
  wire act_mem_banks_bank_a_and_22_cse;
  wire act_mem_banks_bank_a_and_23_cse;
  wire act_mem_banks_bank_a_and_24_cse;
  wire act_mem_banks_bank_a_and_25_cse;
  wire act_mem_banks_bank_a_and_26_cse;
  wire act_mem_banks_bank_a_and_27_cse;
  wire act_mem_banks_bank_a_and_28_cse;
  wire act_mem_banks_bank_a_and_29_cse;
  wire act_mem_banks_bank_a_and_30_cse;
  wire act_mem_banks_bank_a_and_31_cse;
  wire act_config_inst_regs_and_4_cse;
  wire act_config_inst_regs_and_20_cse;
  wire act_mem_banks_read_read_data_and_cse;
  wire act_port_read_out_data_and_cse;
  wire rva_out_reg_data_and_15_cse;
  wire ActUnit_RunInst_switch_lp_and_802_cse;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_and_cse;
  wire act_regs_data_and_124_cse;
  wire act_regs_data_and_128_cse;
  wire act_regs_data_and_132_cse;
  wire act_regs_data_and_136_cse;
  wire act_regs_data_and_140_cse;
  wire act_regs_data_and_144_cse;
  wire act_regs_data_and_148_cse;
  wire act_regs_data_and_152_cse;
  wire act_regs_data_and_156_cse;
  wire act_regs_data_and_160_cse;
  wire act_regs_data_and_164_cse;
  wire act_regs_data_and_168_cse;
  wire act_regs_data_and_172_cse;
  wire act_regs_data_and_176_cse;
  wire act_regs_data_and_180_cse;
  wire act_regs_data_and_184_cse;
  wire act_regs_data_and_188_cse;
  wire act_regs_data_and_192_cse;
  wire act_regs_data_and_196_cse;
  wire act_regs_data_and_200_cse;
  wire act_regs_data_and_204_cse;
  wire act_regs_data_and_208_cse;
  wire act_regs_data_and_212_cse;
  wire act_regs_data_and_216_cse;
  wire act_regs_data_and_220_cse;
  wire act_regs_data_and_224_cse;
  wire act_regs_data_and_228_cse;
  wire act_regs_data_and_232_cse;
  wire act_regs_data_and_236_cse;
  wire act_regs_data_and_240_cse;
  wire act_regs_data_and_244_cse;
  wire act_regs_data_and_248_cse;
  wire act_regs_data_and_252_cse;
  wire act_regs_data_and_256_cse;
  wire act_regs_data_and_260_cse;
  wire act_regs_data_and_264_cse;
  wire act_regs_data_and_268_cse;
  wire act_regs_data_and_272_cse;
  wire act_regs_data_and_276_cse;
  wire act_regs_data_and_280_cse;
  wire act_regs_data_and_284_cse;
  wire act_regs_data_and_288_cse;
  wire act_regs_data_and_292_cse;
  wire act_regs_data_and_296_cse;
  wire act_regs_data_and_300_cse;
  wire act_regs_data_and_304_cse;
  wire act_regs_data_and_308_cse;
  wire act_regs_data_and_312_cse;
  wire act_regs_data_and_316_cse;
  wire act_config_output_counter_and_1_cse;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_and_22_cse;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_and_25_cse;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_and_28_cse;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_and_31_cse;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_and_33_cse;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_and_36_cse;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_and_38_cse;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_and_40_cse;
  wire and_1648_cse;
  wire nor_447_cse;
  wire or_1427_cse;
  wire nor_222_cse;
  wire nor_215_cse;
  reg ActUnit_RunInst_switch_lp_nor_tmp;
  wire Tanh_for_and_2_cse_sva_mx0w0;
  wire ActUnit_RunInst_switch_lp_and_48_tmp_1;
  wire Tanh_for_and_cse_sva_mx0w0;
  wire ActUnit_RunInst_switch_lp_and_32_tmp_mx0w1;
  wire Tanh_for_and_1_cse_sva_mx0w0;
  wire ActUnit_RunInst_switch_lp_and_16_tmp_mx0w1;
  wire ActUnit_RunInst_switch_lp_and_tmp_mx0w0;
  wire Tanh_for_and_85_m1c;
  reg [3:0] reg_act_config_output_counter_sva_dfm_3_ftd;
  wire act_write_data_data_and_ssc;
  wire ActUnit_RunInst_case_2_for_and_27_seb;
  wire while_and_282_cse;
  wire while_and_283_cse;
  reg reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_nor_cse;
  reg reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_2_cse;
  reg reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_1_cse;
  reg reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_cse;
  reg act_config_InstIncr_if_act_config_InstIncr_if_if_nor_mdf_sva;
  wire Tanh_for_or_cse;
  wire Tanh_for_and_87_cse;
  wire [2:0] mux_15_rmff;
  wire [2:0] mux_14_rmff;
  wire [2:0] mux_13_rmff;
  wire [2:0] mux_12_rmff;
  wire [2:0] mux_11_rmff;
  wire [2:0] mux_10_rmff;
  wire [2:0] mux_9_rmff;
  wire [2:0] mux_8_rmff;
  wire [2:0] mux_7_rmff;
  wire [2:0] mux_6_rmff;
  wire [2:0] mux_5_rmff;
  wire [2:0] mux_4_rmff;
  wire [2:0] mux_3_rmff;
  wire [2:0] mux_2_rmff;
  wire [2:0] mux_1_rmff;
  wire [2:0] mux_rmff;
  wire and_1088_rmff;
  wire and_1082_rmff;
  wire and_1076_rmff;
  wire and_1070_rmff;
  wire and_1064_rmff;
  wire and_1058_rmff;
  wire and_1052_rmff;
  wire and_1046_rmff;
  wire and_1040_rmff;
  wire and_1034_rmff;
  wire and_1028_rmff;
  wire and_1022_rmff;
  wire and_1016_rmff;
  wire and_1010_rmff;
  wire and_1004_rmff;
  wire and_998_rmff;
  wire and_990_rmff;
  wire and_985_rmff;
  wire and_980_rmff;
  wire and_975_rmff;
  wire and_970_rmff;
  wire and_965_rmff;
  wire and_960_rmff;
  wire and_955_rmff;
  wire and_950_rmff;
  wire and_945_rmff;
  wire and_940_rmff;
  wire and_935_rmff;
  wire and_930_rmff;
  wire and_925_rmff;
  wire and_920_rmff;
  wire and_915_rmff;
  wire and_906_rmff;
  wire and_905_rmff;
  wire and_904_rmff;
  wire and_903_rmff;
  wire and_902_rmff;
  wire and_901_rmff;
  wire and_900_rmff;
  wire and_899_rmff;
  wire and_1116_rmff;
  wire and_1113_rmff;
  wire and_1108_rmff;
  wire and_1106_rmff;
  wire and_1102_rmff;
  wire and_1097_rmff;
  reg [7:0] act_config_output_addr_base_sva;
  reg [31:0] rva_out_reg_data_511_480_sva_dfm_3;
  wire [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_511_480_mx1;
  reg [31:0] rva_out_reg_data_479_448_sva_dfm_3;
  wire [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_479_448_mx1;
  reg [31:0] rva_out_reg_data_447_416_sva_dfm_3;
  wire [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_447_416_mx1;
  reg [31:0] rva_out_reg_data_415_384_sva_dfm_3;
  wire [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_415_384_mx1;
  reg [31:0] rva_out_reg_data_383_352_sva_dfm_3;
  wire [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_383_352_mx1;
  reg [31:0] rva_out_reg_data_351_320_sva_dfm_3;
  wire [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_351_320_mx1;
  reg [31:0] rva_out_reg_data_319_288_sva_dfm_3;
  wire [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_319_288_mx1;
  reg [31:0] rva_out_reg_data_287_256_sva_dfm_3;
  wire [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_287_256_mx1;
  reg [31:0] rva_out_reg_data_255_224_sva_dfm_3;
  wire [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_255_224_mx1;
  reg [31:0] rva_out_reg_data_223_192_sva_dfm_3;
  wire [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_223_192_mx1;
  reg [31:0] rva_out_reg_data_191_160_sva_dfm_3;
  wire [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_191_160_mx1;
  reg [31:0] rva_out_reg_data_159_128_sva_dfm_3;
  wire [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_159_128_mx1;
  reg [7:0] rva_out_reg_data_127_120_sva_dfm_3;
  wire [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_127_96_mx1;
  reg [7:0] rva_out_reg_data_119_112_sva_dfm_3;
  reg [7:0] rva_out_reg_data_111_104_sva_dfm_3;
  reg [7:0] rva_out_reg_data_103_96_sva_dfm_3;
  reg [7:0] rva_out_reg_data_95_88_sva_dfm_3;
  wire [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_95_64_mx1;
  reg [7:0] rva_out_reg_data_87_80_sva_dfm_3;
  reg [7:0] rva_out_reg_data_79_72_sva_dfm_3;
  reg [7:0] rva_out_reg_data_63_56_sva_dfm_3;
  wire [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_63_32_mx1;
  reg [2:0] rva_out_reg_data_55_53_sva_dfm_3;
  reg [4:0] rva_out_reg_data_52_48_sva_dfm_3;
  reg [7:0] rva_out_reg_data_47_40_sva_dfm_3;
  reg [1:0] rva_out_reg_data_31_30_sva_dfm_3;
  wire [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_31_0_mx1;
  reg [7:0] rva_out_reg_data_23_16_sva_dfm_3;
  reg [6:0] rva_out_reg_data_15_9_sva_dfm_3;
  reg rva_out_reg_data_8_sva_dfm_3;
  reg [6:0] rva_out_reg_data_7_1_sva_dfm_3;
  reg rva_out_reg_data_0_sva_dfm_3;
  reg ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_31;
  wire ActUnit_PushOutput_if_for_and_27_seb_1;
  reg [4:0] ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_30_26;
  reg ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_1_31;
  reg [4:0] ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_1_30_26;
  reg [21:0] Silu_for_2_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0;
  reg ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_1_31;
  reg [4:0] ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_1_30_26;
  reg ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_1_31;
  reg [4:0] ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_1_30_26;
  reg ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_1_31;
  reg [4:0] ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_1_30_26;
  reg ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_1_31;
  reg [4:0] ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_1_30_26;
  reg ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_1_31;
  reg [4:0] ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_1_30_26;
  reg [21:0] Silu_for_y_8_sva_3_21_0;
  reg ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_1_31;
  reg [4:0] ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_1_30_26;
  reg [21:0] Silu_for_y_1_sva_3_21_0;
  reg ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_1_31;
  reg [4:0] ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_1_30_26;
  reg [21:0] Silu_for_9_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0;
  reg ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_1_31;
  reg [4:0] ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_1_30_26;
  reg [21:0] Silu_for_7_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0;
  reg ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_1_31;
  reg [4:0] ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_1_30_26;
  reg [21:0] Silu_for_6_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0;
  reg ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_1_31;
  reg [4:0] ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_1_30_26;
  reg [21:0] Silu_for_5_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0;
  reg ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_1_31;
  reg [4:0] ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_1_30_26;
  reg [21:0] Silu_for_4_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0;
  reg ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_1_31;
  reg [4:0] ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_1_30_26;
  reg [21:0] Silu_for_3_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0;
  reg ActUnit_PushOutput_if_output_port_reg_data_data_1_sva_1_31;
  reg [4:0] rva_out_reg_data_71_64_sva_dfm_6_4_0;
  reg ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_1_31;
  reg [4:0] ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_1_30_26;
  wire and_dcpl_1426;
  wire or_dcpl_1012;
  wire or_dcpl_1013;
  wire or_dcpl_1014;
  wire or_dcpl_1015;
  wire [31:0] ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1;
  wire [22:0] Silu_for_y_8_sva_1_22_0_1;
  wire [23:0] nl_Silu_for_y_8_sva_1_22_0_1;
  wire [22:0] Silu_for_y_7_sva_1_22_0_1;
  wire [23:0] nl_Silu_for_y_7_sva_1_22_0_1;
  wire [22:0] Silu_for_y_6_sva_1_22_0_1;
  wire [23:0] nl_Silu_for_y_6_sva_1_22_0_1;
  wire [22:0] Silu_for_y_5_sva_1_22_0_1;
  wire [23:0] nl_Silu_for_y_5_sva_1_22_0_1;
  wire [22:0] Silu_for_y_4_sva_1_22_0_1;
  wire [23:0] nl_Silu_for_y_4_sva_1_22_0_1;
  wire [22:0] Silu_for_y_3_sva_1_22_0_1;
  wire [23:0] nl_Silu_for_y_3_sva_1_22_0_1;
  wire [22:0] Silu_for_y_2_sva_1_22_0_1;
  wire [23:0] nl_Silu_for_y_2_sva_1_22_0_1;
  wire [22:0] Silu_for_y_1_sva_1_22_0_1;
  wire [23:0] nl_Silu_for_y_1_sva_1_22_0_1;
  reg [511:0] ActUnit_RunInst_case_3_act_port_reg_data_sva;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_291;
  wire act_config_ActConfigRead_else_else_not_21;
  reg [1:0] Silu_for_3_else_else_if_acc_itm;
  wire [2:0] nl_Silu_for_3_else_else_if_acc_itm;
  wire Silu_for_else_and_4_ssc_1;
  wire Silu_for_else_else_else_and_5_ssc_1;
  wire Silu_for_else_and_34_ssc_1;
  wire Silu_for_else_else_else_and_4_ssc_1;
  wire [4:0] ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_30_26_2;
  reg [4:0] act_regs_data_0_1_sva_dfm_2_30_26;
  reg [4:0] act_config_inst_counter_sva;
  reg [3:0] act_config_output_counter_sva_7_4;
  wire [21:0] ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_21_0_mx0w1;
  reg [21:0] act_regs_data_0_7_sva_dfm_2_21_0;
  reg [21:0] act_regs_data_0_14_sva_dfm_2_21_0;
  reg [21:0] act_regs_data_0_15_sva_dfm_2_21_0;
  reg [21:0] act_regs_data_0_2_sva_dfm_2_21_0;
  reg [21:0] act_regs_data_0_3_sva_dfm_2_21_0;
  reg [21:0] act_regs_data_0_4_sva_dfm_2_21_0;
  reg [21:0] act_regs_data_0_5_sva_dfm_2_21_0;
  reg [21:0] act_regs_data_0_8_sva_dfm_2_21_0;
  reg [21:0] act_regs_data_0_6_sva_dfm_2_21_0;
  wire or_1527_tmp;
  wire and_1720_cse;
  wire and_1751_cse;
  wire [5:0] act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_20_itm;
  wire [7:0] act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_21_itm;
  wire [7:0] act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_23_itm;
  wire nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  wire [4:0] nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
  wire [21:0] nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
  wire nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  wire [4:0] nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
  wire [21:0] nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
  wire nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  wire [4:0] nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
  wire [21:0] nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
  wire nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  wire [4:0] nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
  wire [21:0] nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
  wire nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  wire [4:0] nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
  wire [21:0] nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
  wire nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  wire [4:0] nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
  wire [21:0] nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
  wire nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  wire [4:0] nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
  wire [21:0] nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
  wire nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  wire [4:0] nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
  wire [21:0] nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
  wire nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  wire [4:0] nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
  wire [21:0] nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
  wire nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  wire [4:0] nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
  wire [21:0] nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
  wire nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  wire [4:0] nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
  wire [21:0] nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
  wire nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  wire [4:0] nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
  wire [21:0] nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
  wire nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  wire [4:0] nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
  wire [21:0] nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
  wire nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  wire [4:0] nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
  wire [21:0] nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
  wire nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  wire [4:0] nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
  wire [21:0] nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
  wire nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  wire [4:0] nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
  wire [21:0] nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
  wire [31:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_23_itm;
  wire mux_448_itm;
  wire mux_450_itm;
  wire not_tmp_646;
  wire [4:0] z_out;
  wire [5:0] nl_z_out;
  reg [5:0] act_config_num_inst_sva;
  reg [7:0] act_config_num_output_sva;
  reg [4:0] act_config_buffer_addr_base_sva;
  reg ActUnit_DecodeAxi_rva_in_reg_rw_sva;
  reg ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva;
  reg ActUnit_DecodeAxiWrite_else_unequal_tmp;
  reg ActUnit_DecodeAxiRead_else_unequal_tmp;
  reg [4:0] act_write_addrs_lpi_1_dfm_5;
  reg [31:0] act_mem_banks_bank_a_0_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_0_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_0_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_0_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_0_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_0_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_0_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_0_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_0_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_0_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_0_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_0_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_0_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_0_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_0_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_0_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_1_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_1_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_1_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_1_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_1_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_1_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_1_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_1_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_1_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_1_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_1_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_1_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_1_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_1_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_1_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_1_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_2_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_2_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_2_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_2_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_2_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_2_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_2_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_2_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_2_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_2_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_2_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_2_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_2_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_2_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_2_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_2_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_3_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_3_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_3_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_3_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_3_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_3_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_3_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_3_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_3_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_3_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_3_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_3_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_3_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_3_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_3_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_3_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_4_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_4_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_4_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_4_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_4_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_4_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_4_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_4_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_4_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_4_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_4_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_4_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_4_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_4_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_4_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_4_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_5_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_5_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_5_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_5_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_5_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_5_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_5_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_5_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_5_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_5_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_5_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_5_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_5_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_5_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_5_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_5_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_6_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_6_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_6_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_6_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_6_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_6_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_6_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_6_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_6_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_6_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_6_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_6_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_6_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_6_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_6_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_6_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_7_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_7_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_7_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_7_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_7_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_7_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_7_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_7_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_7_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_7_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_7_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_7_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_7_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_7_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_7_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_7_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_8_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_8_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_8_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_8_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_8_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_8_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_8_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_8_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_8_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_8_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_8_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_8_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_8_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_8_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_8_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_8_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_9_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_9_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_9_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_9_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_9_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_9_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_9_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_9_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_9_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_9_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_9_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_9_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_9_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_9_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_9_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_9_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_10_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_10_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_10_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_10_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_10_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_10_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_10_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_10_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_10_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_10_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_10_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_10_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_10_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_10_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_10_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_10_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_11_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_11_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_11_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_11_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_11_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_11_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_11_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_11_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_11_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_11_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_11_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_11_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_11_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_11_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_11_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_11_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_12_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_12_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_12_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_12_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_12_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_12_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_12_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_12_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_12_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_12_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_12_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_12_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_12_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_12_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_12_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_12_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_13_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_13_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_13_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_13_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_13_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_13_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_13_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_13_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_13_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_13_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_13_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_13_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_13_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_13_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_13_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_13_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_14_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_14_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_14_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_14_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_14_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_14_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_14_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_14_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_14_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_14_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_14_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_14_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_14_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_14_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_14_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_14_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_15_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_15_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_15_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_15_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_15_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_15_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_15_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_15_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_15_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_15_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_15_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_15_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_15_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_15_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_15_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_15_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_16_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_16_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_16_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_16_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_16_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_16_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_16_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_16_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_16_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_16_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_16_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_16_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_16_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_16_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_16_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_16_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_17_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_17_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_17_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_17_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_17_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_17_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_17_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_17_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_17_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_17_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_17_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_17_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_17_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_17_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_17_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_17_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_18_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_18_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_18_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_18_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_18_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_18_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_18_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_18_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_18_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_18_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_18_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_18_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_18_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_18_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_18_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_18_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_19_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_19_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_19_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_19_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_19_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_19_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_19_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_19_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_19_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_19_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_19_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_19_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_19_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_19_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_19_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_19_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_20_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_20_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_20_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_20_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_20_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_20_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_20_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_20_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_20_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_20_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_20_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_20_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_20_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_20_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_20_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_20_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_21_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_21_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_21_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_21_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_21_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_21_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_21_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_21_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_21_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_21_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_21_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_21_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_21_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_21_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_21_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_21_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_22_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_22_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_22_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_22_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_22_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_22_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_22_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_22_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_22_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_22_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_22_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_22_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_22_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_22_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_22_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_22_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_23_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_23_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_23_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_23_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_23_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_23_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_23_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_23_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_23_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_23_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_23_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_23_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_23_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_23_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_23_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_23_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_24_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_24_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_24_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_24_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_24_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_24_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_24_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_24_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_24_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_24_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_24_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_24_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_24_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_24_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_24_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_24_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_25_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_25_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_25_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_25_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_25_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_25_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_25_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_25_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_25_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_25_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_25_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_25_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_25_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_25_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_25_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_25_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_26_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_26_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_26_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_26_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_26_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_26_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_26_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_26_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_26_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_26_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_26_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_26_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_26_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_26_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_26_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_26_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_27_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_27_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_27_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_27_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_27_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_27_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_27_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_27_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_27_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_27_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_27_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_27_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_27_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_27_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_27_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_27_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_28_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_28_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_28_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_28_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_28_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_28_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_28_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_28_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_28_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_28_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_28_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_28_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_28_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_28_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_28_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_28_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_29_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_29_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_29_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_29_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_29_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_29_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_29_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_29_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_29_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_29_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_29_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_29_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_29_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_29_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_29_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_29_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_30_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_30_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_30_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_30_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_30_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_30_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_30_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_30_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_30_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_30_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_30_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_30_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_30_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_30_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_30_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_30_31_0_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_31_511_480_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_31_479_448_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_31_447_416_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_31_415_384_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_31_383_352_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_31_351_320_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_31_319_288_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_31_287_256_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_31_255_224_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_31_223_192_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_31_191_160_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_31_159_128_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_31_127_96_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_31_95_64_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_31_63_32_sva_dfm;
  reg [31:0] act_mem_banks_bank_a_31_31_0_sva_dfm;
  reg [31:0] act_port_read_out_data_0_0_sva_dfm;
  reg [31:0] act_port_read_out_data_0_1_sva_dfm;
  reg [31:0] act_port_read_out_data_0_2_sva_dfm;
  reg [31:0] act_port_read_out_data_0_3_sva_dfm;
  reg [31:0] act_port_read_out_data_0_4_sva_dfm;
  reg [31:0] act_port_read_out_data_0_5_sva_dfm;
  reg [31:0] act_port_read_out_data_0_6_sva_dfm;
  reg [31:0] act_port_read_out_data_0_7_sva_dfm;
  reg [31:0] act_port_read_out_data_0_8_sva_dfm;
  reg [31:0] act_port_read_out_data_0_9_sva_dfm;
  reg [31:0] act_port_read_out_data_0_10_sva_dfm;
  reg [31:0] act_port_read_out_data_0_11_sva_dfm;
  reg [31:0] act_port_read_out_data_0_12_sva_dfm;
  reg [31:0] act_port_read_out_data_0_13_sva_dfm;
  reg [31:0] act_port_read_out_data_0_14_sva_dfm;
  reg [31:0] act_port_read_out_data_0_15_sva_dfm;
  reg [1:0] nvhls_get_slc_2U_NVUINT8_return_2_sva;
  reg Silu_for_else_and_1_m1c;
  reg Silu_for_else_and_3_m1c;
  reg Silu_for_else_and_5_m1c;
  reg Silu_for_else_and_7_m1c;
  reg Silu_for_else_and_9_m1c;
  reg Silu_for_else_and_11_m1c;
  reg Silu_for_else_and_13_m1c;
  reg Silu_for_else_and_15_m1c;
  reg Silu_for_else_and_17_m1c;
  reg Silu_for_else_and_19_m1c;
  reg Silu_for_else_and_21_m1c;
  reg Silu_for_else_and_23_m1c;
  reg Silu_for_else_and_25_m1c;
  reg Silu_for_else_and_27_m1c;
  reg Silu_for_else_and_29_m1c;
  reg Silu_for_else_and_31_m1c;
  reg Gelu_for_else_and_1_m1c;
  reg Gelu_for_else_and_3_m1c;
  reg Gelu_for_else_and_5_m1c;
  reg Gelu_for_else_and_7_m1c;
  reg Gelu_for_else_and_9_m1c;
  reg Gelu_for_else_and_11_m1c;
  reg Gelu_for_else_and_13_m1c;
  reg Gelu_for_else_and_15_m1c;
  reg Gelu_for_else_and_17_m1c;
  reg Gelu_for_else_and_19_m1c;
  reg Gelu_for_else_and_21_m1c;
  reg Gelu_for_else_and_23_m1c;
  reg Gelu_for_else_and_25_m1c;
  reg Gelu_for_else_and_27_m1c;
  reg Gelu_for_else_and_29_m1c;
  reg Gelu_for_else_and_31_m1c;
  reg [1:0] Silu_for_1_else_else_if_acc_itm;
  wire [2:0] nl_Silu_for_1_else_else_if_acc_itm;
  reg [1:0] Silu_for_2_else_else_if_acc_itm;
  wire [2:0] nl_Silu_for_2_else_else_if_acc_itm;
  reg [1:0] Silu_for_4_else_else_if_acc_itm;
  wire [2:0] nl_Silu_for_4_else_else_if_acc_itm;
  reg [1:0] Silu_for_5_else_else_if_acc_itm;
  wire [2:0] nl_Silu_for_5_else_else_if_acc_itm;
  reg [1:0] Silu_for_6_else_else_if_acc_itm;
  wire [2:0] nl_Silu_for_6_else_else_if_acc_itm;
  reg [1:0] Silu_for_7_else_else_if_acc_itm;
  wire [2:0] nl_Silu_for_7_else_else_if_acc_itm;
  reg [1:0] Silu_for_8_else_else_if_acc_itm;
  wire [2:0] nl_Silu_for_8_else_else_if_acc_itm;
  reg [1:0] Silu_for_9_else_else_if_acc_itm;
  wire [2:0] nl_Silu_for_9_else_else_if_acc_itm;
  reg [1:0] Silu_for_10_else_else_if_acc_itm;
  wire [2:0] nl_Silu_for_10_else_else_if_acc_itm;
  reg [1:0] Silu_for_11_else_else_if_acc_itm;
  wire [2:0] nl_Silu_for_11_else_else_if_acc_itm;
  reg [1:0] Silu_for_12_else_else_if_acc_itm;
  wire [2:0] nl_Silu_for_12_else_else_if_acc_itm;
  reg [1:0] Silu_for_13_else_else_if_acc_itm;
  wire [2:0] nl_Silu_for_13_else_else_if_acc_itm;
  reg [1:0] Silu_for_14_else_else_if_acc_itm;
  wire [2:0] nl_Silu_for_14_else_else_if_acc_itm;
  reg [1:0] Silu_for_15_else_else_if_acc_itm;
  wire [2:0] nl_Silu_for_15_else_else_if_acc_itm;
  reg [1:0] Silu_for_16_else_else_if_acc_itm;
  wire [2:0] nl_Silu_for_16_else_else_if_acc_itm;
  reg [3:0] Gelu_for_1_else_if_acc_itm;
  reg [3:0] Gelu_for_2_else_if_acc_itm;
  reg [3:0] Gelu_for_3_else_if_acc_itm;
  reg [3:0] Gelu_for_4_else_if_acc_itm;
  reg [3:0] Gelu_for_5_else_if_acc_itm;
  reg [3:0] Gelu_for_6_else_if_acc_itm;
  reg [3:0] Gelu_for_7_else_if_acc_itm;
  reg [3:0] Gelu_for_8_else_if_acc_itm;
  reg [31:0] act_mem_banks_read_for_mux_itm;
  reg [31:0] act_mem_banks_read_for_mux_1_itm;
  reg [31:0] act_mem_banks_read_for_mux_2_itm;
  reg [31:0] act_mem_banks_read_for_mux_3_itm;
  reg [31:0] act_mem_banks_read_for_mux_4_itm;
  reg [31:0] act_mem_banks_read_for_mux_5_itm;
  reg [31:0] act_mem_banks_read_for_mux_6_itm;
  reg [31:0] act_mem_banks_read_for_mux_7_itm;
  reg [31:0] act_mem_banks_read_for_mux_8_itm;
  reg [31:0] act_mem_banks_read_for_mux_9_itm;
  reg [31:0] act_mem_banks_read_for_mux_10_itm;
  reg [31:0] act_mem_banks_read_for_mux_11_itm;
  reg [31:0] act_mem_banks_read_for_mux_12_itm;
  reg [31:0] act_mem_banks_read_for_mux_13_itm;
  reg [31:0] act_mem_banks_read_for_mux_14_itm;
  reg [31:0] act_mem_banks_read_for_mux_15_itm;
  reg while_else_1_mux_1_itm;
  reg Silu_for_y_1_lpi_1_dfm_4_31;
  reg [21:0] Silu_for_y_1_lpi_1_dfm_4_21_0;
  reg Silu_for_y_2_lpi_1_dfm_4_31;
  reg [21:0] Silu_for_y_2_lpi_1_dfm_4_21_0;
  reg Silu_for_y_3_lpi_1_dfm_4_31;
  reg [21:0] Silu_for_y_3_lpi_1_dfm_4_21_0;
  reg Silu_for_y_4_lpi_1_dfm_4_31;
  reg [21:0] Silu_for_y_4_lpi_1_dfm_4_21_0;
  reg Silu_for_y_5_lpi_1_dfm_4_31;
  reg [21:0] Silu_for_y_5_lpi_1_dfm_4_21_0;
  reg Silu_for_y_6_lpi_1_dfm_4_31;
  reg [21:0] Silu_for_y_6_lpi_1_dfm_4_21_0;
  reg Silu_for_y_7_lpi_1_dfm_4_31;
  reg [21:0] Silu_for_y_7_lpi_1_dfm_4_21_0;
  reg Silu_for_y_8_lpi_1_dfm_4_31;
  reg [21:0] Silu_for_y_8_lpi_1_dfm_4_21_0;
  reg act_regs_data_0_0_sva_dfm_2_31;
  reg [4:0] act_regs_data_0_0_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_0_0_sva_dfm_2_21_0;
  reg act_regs_data_0_1_sva_dfm_2_31;
  reg [21:0] act_regs_data_0_1_sva_dfm_2_21_0;
  reg act_regs_data_0_2_sva_dfm_2_31;
  reg [4:0] act_regs_data_0_2_sva_dfm_2_30_26;
  reg act_regs_data_0_3_sva_dfm_2_31;
  reg [4:0] act_regs_data_0_3_sva_dfm_2_30_26;
  reg act_regs_data_0_4_sva_dfm_2_31;
  reg [4:0] act_regs_data_0_4_sva_dfm_2_30_26;
  reg act_regs_data_0_5_sva_dfm_2_31;
  reg [4:0] act_regs_data_0_5_sva_dfm_2_30_26;
  reg act_regs_data_0_6_sva_dfm_2_31;
  reg [4:0] act_regs_data_0_6_sva_dfm_2_30_26;
  reg act_regs_data_0_7_sva_dfm_2_31;
  reg [4:0] act_regs_data_0_7_sva_dfm_2_30_26;
  reg act_regs_data_0_8_sva_dfm_2_31;
  reg [4:0] act_regs_data_0_8_sva_dfm_2_30_26;
  reg act_regs_data_0_9_sva_dfm_2_31;
  reg [4:0] act_regs_data_0_9_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_0_9_sva_dfm_2_21_0;
  reg act_regs_data_0_10_sva_dfm_2_31;
  reg [4:0] act_regs_data_0_10_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_0_10_sva_dfm_2_21_0;
  reg act_regs_data_0_11_sva_dfm_2_31;
  reg [4:0] act_regs_data_0_11_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_0_11_sva_dfm_2_21_0;
  reg act_regs_data_0_12_sva_dfm_2_31;
  reg [4:0] act_regs_data_0_12_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_0_12_sva_dfm_2_21_0;
  reg act_regs_data_0_13_sva_dfm_2_31;
  reg [4:0] act_regs_data_0_13_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_0_13_sva_dfm_2_21_0;
  reg act_regs_data_0_14_sva_dfm_2_31;
  reg [4:0] act_regs_data_0_14_sva_dfm_2_30_26;
  reg act_regs_data_0_15_sva_dfm_2_31;
  reg [4:0] act_regs_data_0_15_sva_dfm_2_30_26;
  reg act_regs_data_1_0_sva_dfm_2_31;
  reg [4:0] act_regs_data_1_0_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_1_0_sva_dfm_2_21_0;
  reg act_regs_data_1_1_sva_dfm_2_31;
  reg [4:0] act_regs_data_1_1_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_1_1_sva_dfm_2_21_0;
  reg act_regs_data_1_2_sva_dfm_2_31;
  reg [4:0] act_regs_data_1_2_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_1_2_sva_dfm_2_21_0;
  reg act_regs_data_1_3_sva_dfm_2_31;
  reg [4:0] act_regs_data_1_3_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_1_3_sva_dfm_2_21_0;
  reg act_regs_data_1_4_sva_dfm_2_31;
  reg [4:0] act_regs_data_1_4_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_1_4_sva_dfm_2_21_0;
  reg act_regs_data_1_5_sva_dfm_2_31;
  reg [4:0] act_regs_data_1_5_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_1_5_sva_dfm_2_21_0;
  reg act_regs_data_1_6_sva_dfm_2_31;
  reg [4:0] act_regs_data_1_6_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_1_6_sva_dfm_2_21_0;
  reg act_regs_data_1_7_sva_dfm_2_31;
  reg [4:0] act_regs_data_1_7_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_1_7_sva_dfm_2_21_0;
  reg act_regs_data_1_8_sva_dfm_2_31;
  reg [4:0] act_regs_data_1_8_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_1_8_sva_dfm_2_21_0;
  reg act_regs_data_1_9_sva_dfm_2_31;
  reg [4:0] act_regs_data_1_9_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_1_9_sva_dfm_2_21_0;
  reg act_regs_data_1_10_sva_dfm_2_31;
  reg [4:0] act_regs_data_1_10_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_1_10_sva_dfm_2_21_0;
  reg act_regs_data_1_11_sva_dfm_2_31;
  reg [4:0] act_regs_data_1_11_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_1_11_sva_dfm_2_21_0;
  reg act_regs_data_1_12_sva_dfm_2_31;
  reg [4:0] act_regs_data_1_12_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_1_12_sva_dfm_2_21_0;
  reg act_regs_data_1_13_sva_dfm_2_31;
  reg [4:0] act_regs_data_1_13_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_1_13_sva_dfm_2_21_0;
  reg act_regs_data_1_14_sva_dfm_2_31;
  reg [4:0] act_regs_data_1_14_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_1_14_sva_dfm_2_21_0;
  reg act_regs_data_1_15_sva_dfm_2_31;
  reg [4:0] act_regs_data_1_15_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_1_15_sva_dfm_2_21_0;
  reg act_regs_data_2_0_sva_dfm_2_31;
  reg [4:0] act_regs_data_2_0_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_2_0_sva_dfm_2_21_0;
  reg act_regs_data_2_1_sva_dfm_2_31;
  reg [4:0] act_regs_data_2_1_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_2_1_sva_dfm_2_21_0;
  reg act_regs_data_2_2_sva_dfm_2_31;
  reg [4:0] act_regs_data_2_2_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_2_2_sva_dfm_2_21_0;
  reg act_regs_data_2_3_sva_dfm_2_31;
  reg [4:0] act_regs_data_2_3_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_2_3_sva_dfm_2_21_0;
  reg act_regs_data_2_4_sva_dfm_2_31;
  reg [4:0] act_regs_data_2_4_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_2_4_sva_dfm_2_21_0;
  reg act_regs_data_2_5_sva_dfm_2_31;
  reg [4:0] act_regs_data_2_5_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_2_5_sva_dfm_2_21_0;
  reg act_regs_data_2_6_sva_dfm_2_31;
  reg [4:0] act_regs_data_2_6_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_2_6_sva_dfm_2_21_0;
  reg act_regs_data_2_7_sva_dfm_2_31;
  reg [4:0] act_regs_data_2_7_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_2_7_sva_dfm_2_21_0;
  reg act_regs_data_2_8_sva_dfm_2_31;
  reg [4:0] act_regs_data_2_8_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_2_8_sva_dfm_2_21_0;
  reg act_regs_data_2_9_sva_dfm_2_31;
  reg [4:0] act_regs_data_2_9_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_2_9_sva_dfm_2_21_0;
  reg act_regs_data_2_10_sva_dfm_2_31;
  reg [4:0] act_regs_data_2_10_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_2_10_sva_dfm_2_21_0;
  reg act_regs_data_2_11_sva_dfm_2_31;
  reg [4:0] act_regs_data_2_11_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_2_11_sva_dfm_2_21_0;
  reg act_regs_data_2_12_sva_dfm_2_31;
  reg [4:0] act_regs_data_2_12_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_2_12_sva_dfm_2_21_0;
  reg act_regs_data_2_13_sva_dfm_2_31;
  reg [4:0] act_regs_data_2_13_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_2_13_sva_dfm_2_21_0;
  reg act_regs_data_2_14_sva_dfm_2_31;
  reg [4:0] act_regs_data_2_14_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_2_14_sva_dfm_2_21_0;
  reg act_regs_data_2_15_sva_dfm_2_31;
  reg [4:0] act_regs_data_2_15_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_2_15_sva_dfm_2_21_0;
  reg act_regs_data_3_0_sva_dfm_2_31;
  reg [4:0] act_regs_data_3_0_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_3_0_sva_dfm_2_21_0;
  reg act_regs_data_3_1_sva_dfm_2_31;
  reg [4:0] act_regs_data_3_1_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_3_1_sva_dfm_2_21_0;
  reg act_regs_data_3_2_sva_dfm_2_31;
  reg [4:0] act_regs_data_3_2_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_3_2_sva_dfm_2_21_0;
  reg act_regs_data_3_3_sva_dfm_2_31;
  reg [4:0] act_regs_data_3_3_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_3_3_sva_dfm_2_21_0;
  reg act_regs_data_3_4_sva_dfm_2_31;
  reg [4:0] act_regs_data_3_4_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_3_4_sva_dfm_2_21_0;
  reg act_regs_data_3_5_sva_dfm_2_31;
  reg [4:0] act_regs_data_3_5_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_3_5_sva_dfm_2_21_0;
  reg act_regs_data_3_6_sva_dfm_2_31;
  reg [4:0] act_regs_data_3_6_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_3_6_sva_dfm_2_21_0;
  reg act_regs_data_3_7_sva_dfm_2_31;
  reg [4:0] act_regs_data_3_7_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_3_7_sva_dfm_2_21_0;
  reg act_regs_data_3_8_sva_dfm_2_31;
  reg [4:0] act_regs_data_3_8_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_3_8_sva_dfm_2_21_0;
  reg act_regs_data_3_9_sva_dfm_2_31;
  reg [4:0] act_regs_data_3_9_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_3_9_sva_dfm_2_21_0;
  reg act_regs_data_3_10_sva_dfm_2_31;
  reg [4:0] act_regs_data_3_10_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_3_10_sva_dfm_2_21_0;
  reg act_regs_data_3_11_sva_dfm_2_31;
  reg [4:0] act_regs_data_3_11_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_3_11_sva_dfm_2_21_0;
  reg act_regs_data_3_12_sva_dfm_2_31;
  reg [4:0] act_regs_data_3_12_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_3_12_sva_dfm_2_21_0;
  reg act_regs_data_3_13_sva_dfm_2_31;
  reg [4:0] act_regs_data_3_13_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_3_13_sva_dfm_2_21_0;
  reg act_regs_data_3_14_sva_dfm_2_31;
  reg [4:0] act_regs_data_3_14_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_3_14_sva_dfm_2_21_0;
  reg act_regs_data_3_15_sva_dfm_2_31;
  reg [4:0] act_regs_data_3_15_sva_dfm_2_30_26;
  reg [21:0] act_regs_data_3_15_sva_dfm_2_21_0;
  reg [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_511_480;
  reg [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_479_448;
  reg [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_447_416;
  reg [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_415_384;
  reg [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_383_352;
  reg [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_351_320;
  reg [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_319_288;
  reg [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_287_256;
  reg [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_255_224;
  reg [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_223_192;
  reg [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_191_160;
  reg [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_159_128;
  reg [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_127_96;
  reg [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_95_64;
  reg [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_63_32;
  reg [31:0] act_mem_banks_read_read_data_lpi_1_dfm_1_31_0;
  reg act_regs_data_1_15_sva_8_31;
  reg [4:0] act_regs_data_1_15_sva_8_30_26;
  reg [21:0] act_regs_data_1_15_sva_8_21_0;
  reg act_regs_data_2_0_sva_8_31;
  reg [4:0] act_regs_data_2_0_sva_8_30_26;
  reg [21:0] act_regs_data_2_0_sva_8_21_0;
  reg act_regs_data_1_14_sva_8_31;
  reg [4:0] act_regs_data_1_14_sva_8_30_26;
  reg [21:0] act_regs_data_1_14_sva_8_21_0;
  reg act_regs_data_2_1_sva_8_31;
  reg [4:0] act_regs_data_2_1_sva_8_30_26;
  reg [21:0] act_regs_data_2_1_sva_8_21_0;
  reg act_regs_data_1_13_sva_8_31;
  reg [4:0] act_regs_data_1_13_sva_8_30_26;
  reg [21:0] act_regs_data_1_13_sva_8_21_0;
  reg act_regs_data_2_2_sva_8_31;
  reg [4:0] act_regs_data_2_2_sva_8_30_26;
  reg [21:0] act_regs_data_2_2_sva_8_21_0;
  reg act_regs_data_1_12_sva_8_31;
  reg [4:0] act_regs_data_1_12_sva_8_30_26;
  reg [21:0] act_regs_data_1_12_sva_8_21_0;
  reg act_regs_data_2_3_sva_8_31;
  reg [4:0] act_regs_data_2_3_sva_8_30_26;
  reg [21:0] act_regs_data_2_3_sva_8_21_0;
  reg act_regs_data_1_11_sva_8_31;
  reg [4:0] act_regs_data_1_11_sva_8_30_26;
  reg [21:0] act_regs_data_1_11_sva_8_21_0;
  reg act_regs_data_2_4_sva_8_31;
  reg [4:0] act_regs_data_2_4_sva_8_30_26;
  reg [21:0] act_regs_data_2_4_sva_8_21_0;
  reg act_regs_data_1_10_sva_8_31;
  reg [4:0] act_regs_data_1_10_sva_8_30_26;
  reg [21:0] act_regs_data_1_10_sva_8_21_0;
  reg act_regs_data_2_5_sva_8_31;
  reg [4:0] act_regs_data_2_5_sva_8_30_26;
  reg [21:0] act_regs_data_2_5_sva_8_21_0;
  reg act_regs_data_1_9_sva_8_31;
  reg [4:0] act_regs_data_1_9_sva_8_30_26;
  reg [21:0] act_regs_data_1_9_sva_8_21_0;
  reg act_regs_data_2_6_sva_8_31;
  reg [4:0] act_regs_data_2_6_sva_8_30_26;
  reg [21:0] act_regs_data_2_6_sva_8_21_0;
  reg act_regs_data_1_8_sva_8_31;
  reg [4:0] act_regs_data_1_8_sva_8_30_26;
  reg [21:0] act_regs_data_1_8_sva_8_21_0;
  reg act_regs_data_2_7_sva_8_31;
  reg [4:0] act_regs_data_2_7_sva_8_30_26;
  reg [21:0] act_regs_data_2_7_sva_8_21_0;
  reg act_regs_data_1_7_sva_8_31;
  reg [4:0] act_regs_data_1_7_sva_8_30_26;
  reg [21:0] act_regs_data_1_7_sva_8_21_0;
  reg act_regs_data_2_8_sva_8_31;
  reg [4:0] act_regs_data_2_8_sva_8_30_26;
  reg [21:0] act_regs_data_2_8_sva_8_21_0;
  reg act_regs_data_1_6_sva_8_31;
  reg [4:0] act_regs_data_1_6_sva_8_30_26;
  reg [21:0] act_regs_data_1_6_sva_8_21_0;
  reg act_regs_data_2_9_sva_8_31;
  reg [4:0] act_regs_data_2_9_sva_8_30_26;
  reg [21:0] act_regs_data_2_9_sva_8_21_0;
  reg act_regs_data_1_5_sva_8_31;
  reg [4:0] act_regs_data_1_5_sva_8_30_26;
  reg [21:0] act_regs_data_1_5_sva_8_21_0;
  reg act_regs_data_2_10_sva_8_31;
  reg [4:0] act_regs_data_2_10_sva_8_30_26;
  reg [21:0] act_regs_data_2_10_sva_8_21_0;
  reg act_regs_data_1_4_sva_8_31;
  reg [4:0] act_regs_data_1_4_sva_8_30_26;
  reg [21:0] act_regs_data_1_4_sva_8_21_0;
  reg act_regs_data_2_11_sva_8_31;
  reg [4:0] act_regs_data_2_11_sva_8_30_26;
  reg [21:0] act_regs_data_2_11_sva_8_21_0;
  reg act_regs_data_1_3_sva_8_31;
  reg [4:0] act_regs_data_1_3_sva_8_30_26;
  reg [21:0] act_regs_data_1_3_sva_8_21_0;
  reg act_regs_data_2_12_sva_8_31;
  reg [4:0] act_regs_data_2_12_sva_8_30_26;
  reg [21:0] act_regs_data_2_12_sva_8_21_0;
  reg act_regs_data_1_2_sva_8_31;
  reg [4:0] act_regs_data_1_2_sva_8_30_26;
  reg [21:0] act_regs_data_1_2_sva_8_21_0;
  reg act_regs_data_2_13_sva_8_31;
  reg [4:0] act_regs_data_2_13_sva_8_30_26;
  reg [21:0] act_regs_data_2_13_sva_8_21_0;
  reg act_regs_data_1_1_sva_8_31;
  reg [4:0] act_regs_data_1_1_sva_8_30_26;
  reg [21:0] act_regs_data_1_1_sva_8_21_0;
  reg act_regs_data_2_14_sva_8_31;
  reg [4:0] act_regs_data_2_14_sva_8_30_26;
  reg [21:0] act_regs_data_2_14_sva_8_21_0;
  reg act_regs_data_1_0_sva_8_31;
  reg [4:0] act_regs_data_1_0_sva_8_30_26;
  reg [21:0] act_regs_data_1_0_sva_8_21_0;
  reg act_regs_data_2_15_sva_8_31;
  reg [4:0] act_regs_data_2_15_sva_8_30_26;
  reg [21:0] act_regs_data_2_15_sva_8_21_0;
  reg act_regs_data_0_15_sva_8_31;
  reg [4:0] act_regs_data_0_15_sva_8_30_26;
  reg [21:0] act_regs_data_0_15_sva_8_21_0;
  reg act_regs_data_3_0_sva_8_31;
  reg [4:0] act_regs_data_3_0_sva_8_30_26;
  reg [21:0] act_regs_data_3_0_sva_8_21_0;
  reg act_regs_data_0_14_sva_8_31;
  reg [4:0] act_regs_data_0_14_sva_8_30_26;
  reg [21:0] act_regs_data_0_14_sva_8_21_0;
  reg act_regs_data_3_1_sva_8_31;
  reg [4:0] act_regs_data_3_1_sva_8_30_26;
  reg [21:0] act_regs_data_3_1_sva_8_21_0;
  reg act_regs_data_0_13_sva_8_31;
  reg [4:0] act_regs_data_0_13_sva_8_30_26;
  reg [21:0] act_regs_data_0_13_sva_8_21_0;
  reg act_regs_data_3_2_sva_8_31;
  reg [4:0] act_regs_data_3_2_sva_8_30_26;
  reg [21:0] act_regs_data_3_2_sva_8_21_0;
  reg act_regs_data_0_12_sva_8_31;
  reg [4:0] act_regs_data_0_12_sva_8_30_26;
  reg [21:0] act_regs_data_0_12_sva_8_21_0;
  reg act_regs_data_3_3_sva_8_31;
  reg [4:0] act_regs_data_3_3_sva_8_30_26;
  reg [21:0] act_regs_data_3_3_sva_8_21_0;
  reg act_regs_data_0_11_sva_8_31;
  reg [4:0] act_regs_data_0_11_sva_8_30_26;
  reg [21:0] act_regs_data_0_11_sva_8_21_0;
  reg act_regs_data_3_4_sva_8_31;
  reg [4:0] act_regs_data_3_4_sva_8_30_26;
  reg [21:0] act_regs_data_3_4_sva_8_21_0;
  reg act_regs_data_0_10_sva_8_31;
  reg [4:0] act_regs_data_0_10_sva_8_30_26;
  reg [21:0] act_regs_data_0_10_sva_8_21_0;
  reg act_regs_data_3_5_sva_8_31;
  reg [4:0] act_regs_data_3_5_sva_8_30_26;
  reg [21:0] act_regs_data_3_5_sva_8_21_0;
  reg act_regs_data_0_9_sva_8_31;
  reg [4:0] act_regs_data_0_9_sva_8_30_26;
  reg [21:0] act_regs_data_0_9_sva_8_21_0;
  reg act_regs_data_3_6_sva_8_31;
  reg [4:0] act_regs_data_3_6_sva_8_30_26;
  reg [21:0] act_regs_data_3_6_sva_8_21_0;
  reg act_regs_data_0_8_sva_8_31;
  reg [4:0] act_regs_data_0_8_sva_8_30_26;
  reg [21:0] act_regs_data_0_8_sva_8_21_0;
  reg act_regs_data_3_7_sva_8_31;
  reg [4:0] act_regs_data_3_7_sva_8_30_26;
  reg [21:0] act_regs_data_3_7_sva_8_21_0;
  reg act_regs_data_0_7_sva_8_31;
  reg [4:0] act_regs_data_0_7_sva_8_30_26;
  reg [21:0] act_regs_data_0_7_sva_8_21_0;
  reg act_regs_data_3_8_sva_8_31;
  reg [4:0] act_regs_data_3_8_sva_8_30_26;
  reg [21:0] act_regs_data_3_8_sva_8_21_0;
  reg act_regs_data_0_6_sva_8_31;
  reg [4:0] act_regs_data_0_6_sva_8_30_26;
  reg [21:0] act_regs_data_0_6_sva_8_21_0;
  reg act_regs_data_3_9_sva_8_31;
  reg [4:0] act_regs_data_3_9_sva_8_30_26;
  reg [21:0] act_regs_data_3_9_sva_8_21_0;
  reg act_regs_data_0_5_sva_8_31;
  reg [4:0] act_regs_data_0_5_sva_8_30_26;
  reg [21:0] act_regs_data_0_5_sva_8_21_0;
  reg act_regs_data_3_10_sva_8_31;
  reg [4:0] act_regs_data_3_10_sva_8_30_26;
  reg [21:0] act_regs_data_3_10_sva_8_21_0;
  reg act_regs_data_0_4_sva_8_31;
  reg [4:0] act_regs_data_0_4_sva_8_30_26;
  reg [21:0] act_regs_data_0_4_sva_8_21_0;
  reg act_regs_data_3_11_sva_8_31;
  reg [4:0] act_regs_data_3_11_sva_8_30_26;
  reg [21:0] act_regs_data_3_11_sva_8_21_0;
  reg act_regs_data_0_3_sva_8_31;
  reg [4:0] act_regs_data_0_3_sva_8_30_26;
  reg [21:0] act_regs_data_0_3_sva_8_21_0;
  reg act_regs_data_3_12_sva_8_31;
  reg [4:0] act_regs_data_3_12_sva_8_30_26;
  reg [21:0] act_regs_data_3_12_sva_8_21_0;
  reg act_regs_data_0_2_sva_8_31;
  reg [4:0] act_regs_data_0_2_sva_8_30_26;
  reg [21:0] act_regs_data_0_2_sva_8_21_0;
  reg act_regs_data_3_13_sva_8_31;
  reg [4:0] act_regs_data_3_13_sva_8_30_26;
  reg [21:0] act_regs_data_3_13_sva_8_21_0;
  reg act_regs_data_0_1_sva_8_31;
  reg [4:0] act_regs_data_0_1_sva_8_30_26;
  reg [21:0] act_regs_data_0_1_sva_8_21_0;
  reg act_regs_data_3_14_sva_8_31;
  reg [4:0] act_regs_data_3_14_sva_8_30_26;
  reg [21:0] act_regs_data_3_14_sva_8_21_0;
  reg act_regs_data_0_0_sva_8_31;
  reg [4:0] act_regs_data_0_0_sva_8_30_26;
  reg [21:0] act_regs_data_0_0_sva_8_21_0;
  reg act_regs_data_3_15_sva_8_31;
  reg [4:0] act_regs_data_3_15_sva_8_30_26;
  reg [21:0] act_regs_data_3_15_sva_8_21_0;
  reg act_config_inst_regs_16_sva_0;
  reg act_config_inst_regs_17_sva_0;
  reg act_config_inst_regs_1_sva_0;
  reg act_config_inst_regs_0_sva_0;
  wire ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0;
  wire rva_out_reg_data_39_32_sva_dfm_6_mx0c0;
  wire act_config_output_counter_sva_mx0c0;
  wire act_config_output_counter_sva_mx0c1;
  wire act_config_output_counter_sva_mx0c2;
  wire act_config_inst_counter_sva_mx0c1;
  wire [3:0] Gelu_for_1_else_if_acc_itm_mx1w0;
  wire [4:0] nl_Gelu_for_1_else_if_acc_itm_mx1w0;
  wire [3:0] Gelu_for_2_else_if_acc_itm_mx1w0;
  wire [4:0] nl_Gelu_for_2_else_if_acc_itm_mx1w0;
  wire [3:0] Gelu_for_3_else_if_acc_itm_mx1w0;
  wire [4:0] nl_Gelu_for_3_else_if_acc_itm_mx1w0;
  wire [3:0] Gelu_for_4_else_if_acc_itm_mx1w0;
  wire [4:0] nl_Gelu_for_4_else_if_acc_itm_mx1w0;
  wire [3:0] Gelu_for_5_else_if_acc_itm_mx1w0;
  wire [4:0] nl_Gelu_for_5_else_if_acc_itm_mx1w0;
  wire [3:0] Gelu_for_6_else_if_acc_itm_mx1w0;
  wire [4:0] nl_Gelu_for_6_else_if_acc_itm_mx1w0;
  wire [3:0] Gelu_for_7_else_if_acc_itm_mx1w0;
  wire [4:0] nl_Gelu_for_7_else_if_acc_itm_mx1w0;
  wire [3:0] Gelu_for_8_else_if_acc_itm_mx1w0;
  wire [4:0] nl_Gelu_for_8_else_if_acc_itm_mx1w0;
  wire Silu_for_else_and_17_m1c_mx0w1;
  wire Silu_for_else_and_21_m1c_mx0w1;
  wire Silu_for_else_and_23_m1c_mx0w1;
  wire Silu_for_else_and_25_m1c_mx0w1;
  wire Silu_for_else_and_27_m1c_mx0w1;
  wire Silu_for_else_and_29_m1c_mx0w1;
  wire Silu_for_else_and_31_m1c_mx0w1;
  wire [4:0] act_read_addrs_sva_2_mx0w0;
  wire [5:0] nl_act_read_addrs_sva_2_mx0w0;
  wire [4:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_2_mx0w2;
  wire Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs_mx0w0;
  wire Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs_mx0w0;
  wire Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs_mx0w0;
  wire Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs_mx0w0;
  wire Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs_mx0w0;
  wire Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs_mx0w0;
  wire Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs_mx0w0;
  wire Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs_mx0w0;
  wire ActUnit_RunInst_switch_lp_equal_tmp_9;
  wire ActUnit_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva_mx0c4;
  wire ActUnit_PushOutput_if_for_i_4_0_sva_3_0_mx0c0;
  wire [4:0] while_mux_53_ssc_mx0;
  wire [4:0] act_read_addrs_lpi_1_dfm_7;
  wire [31:0] act_write_data_data_0_0_lpi_1_dfm_7;
  wire [31:0] act_write_data_data_0_1_lpi_1_dfm_7;
  wire [31:0] act_write_data_data_0_2_lpi_1_dfm_7;
  wire [31:0] act_write_data_data_0_3_lpi_1_dfm_7;
  wire [31:0] act_write_data_data_0_4_lpi_1_dfm_7;
  wire [31:0] act_write_data_data_0_5_lpi_1_dfm_7;
  wire [31:0] act_write_data_data_0_6_lpi_1_dfm_7;
  wire [31:0] act_write_data_data_0_7_lpi_1_dfm_7;
  wire [31:0] act_write_data_data_0_8_lpi_1_dfm_7;
  wire [31:0] act_write_data_data_0_9_lpi_1_dfm_7;
  wire [31:0] act_write_data_data_0_10_lpi_1_dfm_7;
  wire [31:0] act_write_data_data_0_11_lpi_1_dfm_7;
  wire [31:0] act_write_data_data_0_12_lpi_1_dfm_7;
  wire [31:0] act_write_data_data_0_13_lpi_1_dfm_7;
  wire [31:0] act_write_data_data_0_14_lpi_1_dfm_7;
  wire [31:0] act_write_data_data_0_15_lpi_1_dfm_7;
  wire while_asn_2035;
  wire while_asn_2037;
  wire while_asn_2039;
  wire Silu_for_else_and_ssc_1;
  wire Silu_for_else_else_else_and_1_ssc_1;
  wire Silu_for_else_and_2_ssc_1;
  wire Silu_for_else_else_else_and_3_ssc_1;
  wire Silu_for_else_and_6_ssc_1;
  wire Silu_for_else_else_else_and_7_ssc_1;
  wire Silu_for_else_and_8_ssc_1;
  wire Silu_for_else_else_else_and_9_ssc_1;
  wire Silu_for_else_and_10_ssc_1;
  wire Silu_for_else_else_else_and_11_ssc_1;
  wire Silu_for_else_and_12_ssc_1;
  wire Silu_for_else_else_else_and_13_ssc_1;
  wire Silu_for_else_and_14_ssc_1;
  wire Silu_for_else_else_else_and_15_ssc_1;
  wire Silu_for_else_and_39_ssc_1;
  wire Silu_for_else_else_else_and_14_ssc_1;
  wire Silu_for_else_and_38_ssc_1;
  wire Silu_for_else_else_else_and_12_ssc_1;
  wire Silu_for_else_and_37_ssc_1;
  wire Silu_for_else_else_else_and_10_ssc_1;
  wire Silu_for_else_and_36_ssc_1;
  wire Silu_for_else_else_else_and_8_ssc_1;
  wire Silu_for_else_and_35_ssc_1;
  wire Silu_for_else_else_else_and_6_ssc_1;
  wire Silu_for_else_and_33_ssc_1;
  wire Silu_for_else_else_else_and_2_ssc_1;
  wire Silu_for_else_and_32_ssc_1;
  wire Silu_for_else_else_else_and_ssc_1;
  wire Silu_for_y_lpi_1_dfm_4_31_1;
  wire [21:0] Silu_for_y_lpi_1_dfm_4_21_0_1;
  wire [4:0] Silu_for_y_lpi_1_dfm_4_30_26_1;
  wire Silu_for_y_15_lpi_1_dfm_4_31_1;
  wire [21:0] Silu_for_y_15_lpi_1_dfm_4_21_0_1;
  wire [4:0] Silu_for_y_15_lpi_1_dfm_4_30_26_1;
  wire Silu_for_y_14_lpi_1_dfm_4_31_1;
  wire [21:0] Silu_for_y_14_lpi_1_dfm_4_21_0_1;
  wire [4:0] Silu_for_y_14_lpi_1_dfm_4_30_26_1;
  wire Silu_for_y_13_lpi_1_dfm_4_31_1;
  wire [21:0] Silu_for_y_13_lpi_1_dfm_4_21_0_1;
  wire [4:0] Silu_for_y_13_lpi_1_dfm_4_30_26_1;
  wire Silu_for_y_12_lpi_1_dfm_4_31_1;
  wire [21:0] Silu_for_y_12_lpi_1_dfm_4_21_0_1;
  wire [4:0] Silu_for_y_12_lpi_1_dfm_4_30_26_1;
  wire Silu_for_y_11_lpi_1_dfm_4_31_1;
  wire [21:0] Silu_for_y_11_lpi_1_dfm_4_21_0_1;
  wire [4:0] Silu_for_y_11_lpi_1_dfm_4_30_26_1;
  wire Silu_for_y_10_lpi_1_dfm_4_31_1;
  wire [21:0] Silu_for_y_10_lpi_1_dfm_4_21_0_1;
  wire [4:0] Silu_for_y_10_lpi_1_dfm_4_30_26_1;
  wire Silu_for_y_9_lpi_1_dfm_4_31_1;
  wire [21:0] Silu_for_y_9_lpi_1_dfm_4_21_0_1;
  wire [4:0] Silu_for_y_9_lpi_1_dfm_4_30_26_1;
  wire Gelu_for_y_lpi_1_dfm_4_31_1;
  wire [21:0] Gelu_for_y_lpi_1_dfm_4_21_0_1;
  wire Gelu_for_y_15_lpi_1_dfm_4_31_1;
  wire [21:0] Gelu_for_y_15_lpi_1_dfm_4_21_0_1;
  wire Gelu_for_y_14_lpi_1_dfm_4_31_1;
  wire [21:0] Gelu_for_y_14_lpi_1_dfm_4_21_0_1;
  wire Gelu_for_y_13_lpi_1_dfm_4_31_1;
  wire [21:0] Gelu_for_y_13_lpi_1_dfm_4_21_0_1;
  wire Gelu_for_y_12_lpi_1_dfm_4_31_1;
  wire [21:0] Gelu_for_y_12_lpi_1_dfm_4_21_0_1;
  wire Gelu_for_y_11_lpi_1_dfm_4_31_1;
  wire [21:0] Gelu_for_y_11_lpi_1_dfm_4_21_0_1;
  wire Gelu_for_y_10_lpi_1_dfm_4_31_1;
  wire [21:0] Gelu_for_y_10_lpi_1_dfm_4_21_0_1;
  wire Gelu_for_y_9_lpi_1_dfm_4_31_1;
  wire [21:0] Gelu_for_y_9_lpi_1_dfm_4_21_0_1;
  wire Gelu_for_y_8_lpi_1_dfm_4_31_1;
  wire [21:0] Gelu_for_y_8_lpi_1_dfm_4_21_0_1;
  wire Gelu_for_y_7_lpi_1_dfm_4_31_1;
  wire [21:0] Gelu_for_y_7_lpi_1_dfm_4_21_0_1;
  wire Gelu_for_y_6_lpi_1_dfm_4_31_1;
  wire [21:0] Gelu_for_y_6_lpi_1_dfm_4_21_0_1;
  wire Gelu_for_y_5_lpi_1_dfm_4_31_1;
  wire [21:0] Gelu_for_y_5_lpi_1_dfm_4_21_0_1;
  wire Gelu_for_y_4_lpi_1_dfm_4_31_1;
  wire [21:0] Gelu_for_y_4_lpi_1_dfm_4_21_0_1;
  wire Gelu_for_y_3_lpi_1_dfm_4_31_1;
  wire [21:0] Gelu_for_y_3_lpi_1_dfm_4_21_0_1;
  wire Gelu_for_y_2_lpi_1_dfm_4_31_1;
  wire [21:0] Gelu_for_y_2_lpi_1_dfm_4_21_0_1;
  wire Gelu_for_y_1_lpi_1_dfm_4_31_1;
  wire [21:0] Gelu_for_y_1_lpi_1_dfm_4_21_0_1;
  wire Silu_for_else_and_16_ssc_1;
  wire Silu_for_else_else_else_and_17_ssc_1;
  wire Silu_for_else_and_18_ssc_1;
  wire Silu_for_else_else_else_and_19_ssc_1;
  wire Silu_for_else_and_20_ssc_1;
  wire Silu_for_else_else_else_and_21_ssc_1;
  wire Silu_for_else_and_22_ssc_1;
  wire Silu_for_else_else_else_and_23_ssc_1;
  wire Silu_for_else_and_24_ssc_1;
  wire Silu_for_else_else_else_and_25_ssc_1;
  wire Silu_for_else_and_26_ssc_1;
  wire Silu_for_else_else_else_and_27_ssc_1;
  wire Silu_for_else_and_28_ssc_1;
  wire Silu_for_else_else_else_and_29_ssc_1;
  wire Silu_for_else_and_30_ssc_1;
  wire Silu_for_else_else_else_and_31_ssc_1;
  wire Silu_for_else_and_47_ssc_1;
  wire Silu_for_else_else_else_and_30_ssc_1;
  wire Silu_for_else_and_46_ssc_1;
  wire Silu_for_else_else_else_and_28_ssc_1;
  wire Silu_for_else_and_45_ssc_1;
  wire Silu_for_else_else_else_and_26_ssc_1;
  wire Silu_for_else_and_44_ssc_1;
  wire Silu_for_else_else_else_and_24_ssc_1;
  wire Silu_for_else_and_43_ssc_1;
  wire Silu_for_else_else_else_and_22_ssc_1;
  wire Silu_for_else_and_42_ssc_1;
  wire Silu_for_else_else_else_and_20_ssc_1;
  wire Silu_for_else_and_41_ssc_1;
  wire Silu_for_else_else_else_and_18_ssc_1;
  wire Silu_for_else_and_40_ssc_1;
  wire Silu_for_else_else_else_and_16_ssc_1;
  wire [5:0] Gelu_for_y_1_sva_4_27_22_1;
  wire [6:0] nl_Gelu_for_y_1_sva_4_27_22_1;
  wire [5:0] Gelu_for_y_2_sva_4_27_22_1;
  wire [6:0] nl_Gelu_for_y_2_sva_4_27_22_1;
  wire [5:0] Gelu_for_y_3_sva_4_27_22_1;
  wire [6:0] nl_Gelu_for_y_3_sva_4_27_22_1;
  wire [5:0] Gelu_for_y_4_sva_4_27_22_1;
  wire [6:0] nl_Gelu_for_y_4_sva_4_27_22_1;
  wire [5:0] Gelu_for_y_5_sva_4_27_22_1;
  wire [6:0] nl_Gelu_for_y_5_sva_4_27_22_1;
  wire [5:0] Gelu_for_y_6_sva_4_27_22_1;
  wire [6:0] nl_Gelu_for_y_6_sva_4_27_22_1;
  wire [5:0] Gelu_for_y_7_sva_4_27_22_1;
  wire [6:0] nl_Gelu_for_y_7_sva_4_27_22_1;
  wire [5:0] Gelu_for_y_8_sva_4_27_22_1;
  wire [6:0] nl_Gelu_for_y_8_sva_4_27_22_1;
  wire [5:0] Gelu_for_y_9_sva_4_27_22_1;
  wire [6:0] nl_Gelu_for_y_9_sva_4_27_22_1;
  wire [5:0] Gelu_for_y_10_sva_4_27_22_1;
  wire [6:0] nl_Gelu_for_y_10_sva_4_27_22_1;
  wire [5:0] Gelu_for_y_11_sva_4_27_22_1;
  wire [6:0] nl_Gelu_for_y_11_sva_4_27_22_1;
  wire [5:0] Gelu_for_y_12_sva_4_27_22_1;
  wire [6:0] nl_Gelu_for_y_12_sva_4_27_22_1;
  wire [5:0] Gelu_for_y_13_sva_4_27_22_1;
  wire [6:0] nl_Gelu_for_y_13_sva_4_27_22_1;
  wire [5:0] Gelu_for_y_14_sva_4_27_22_1;
  wire [6:0] nl_Gelu_for_y_14_sva_4_27_22_1;
  wire [5:0] Gelu_for_y_15_sva_4_27_22_1;
  wire [6:0] nl_Gelu_for_y_15_sva_4_27_22_1;
  wire [5:0] Gelu_for_y_sva_4_27_22_1;
  wire [6:0] nl_Gelu_for_y_sva_4_27_22_1;
  wire Gelu_for_else_and_30_ssc_1;
  wire Gelu_for_else_else_else_and_30_ssc_1;
  wire Gelu_for_else_and_47_ssc_1;
  wire Gelu_for_else_else_else_and_31_ssc_1;
  wire Gelu_for_else_and_28_ssc_1;
  wire Gelu_for_else_else_else_and_28_ssc_1;
  wire Gelu_for_else_and_46_ssc_1;
  wire Gelu_for_else_else_else_and_29_ssc_1;
  wire Gelu_for_else_and_26_ssc_1;
  wire Gelu_for_else_else_else_and_26_ssc_1;
  wire Gelu_for_else_and_45_ssc_1;
  wire Gelu_for_else_else_else_and_27_ssc_1;
  wire Gelu_for_else_and_24_ssc_1;
  wire Gelu_for_else_else_else_and_24_ssc_1;
  wire Gelu_for_else_and_44_ssc_1;
  wire Gelu_for_else_else_else_and_25_ssc_1;
  wire Gelu_for_else_and_22_ssc_1;
  wire Gelu_for_else_else_else_and_22_ssc_1;
  wire Gelu_for_else_and_43_ssc_1;
  wire Gelu_for_else_else_else_and_23_ssc_1;
  wire Gelu_for_else_and_20_ssc_1;
  wire Gelu_for_else_else_else_and_20_ssc_1;
  wire Gelu_for_else_and_42_ssc_1;
  wire Gelu_for_else_else_else_and_21_ssc_1;
  wire Gelu_for_else_and_18_ssc_1;
  wire Gelu_for_else_else_else_and_18_ssc_1;
  wire Gelu_for_else_and_41_ssc_1;
  wire Gelu_for_else_else_else_and_19_ssc_1;
  wire Gelu_for_else_and_16_ssc_1;
  wire Gelu_for_else_else_else_and_16_ssc_1;
  wire Gelu_for_else_and_40_ssc_1;
  wire Gelu_for_else_else_else_and_17_ssc_1;
  wire Gelu_for_else_and_14_ssc_1;
  wire Gelu_for_else_else_else_and_14_ssc_1;
  wire Gelu_for_else_and_39_ssc_1;
  wire Gelu_for_else_else_else_and_15_ssc_1;
  wire Gelu_for_else_and_12_ssc_1;
  wire Gelu_for_else_else_else_and_12_ssc_1;
  wire Gelu_for_else_and_38_ssc_1;
  wire Gelu_for_else_else_else_and_13_ssc_1;
  wire Gelu_for_else_and_10_ssc_1;
  wire Gelu_for_else_else_else_and_10_ssc_1;
  wire Gelu_for_else_and_37_ssc_1;
  wire Gelu_for_else_else_else_and_11_ssc_1;
  wire Gelu_for_else_and_8_ssc_1;
  wire Gelu_for_else_else_else_and_8_ssc_1;
  wire Gelu_for_else_and_36_ssc_1;
  wire Gelu_for_else_else_else_and_9_ssc_1;
  wire Gelu_for_else_and_6_ssc_1;
  wire Gelu_for_else_else_else_and_6_ssc_1;
  wire Gelu_for_else_and_35_ssc_1;
  wire Gelu_for_else_else_else_and_7_ssc_1;
  wire Gelu_for_else_and_4_ssc_1;
  wire Gelu_for_else_else_else_and_4_ssc_1;
  wire Gelu_for_else_and_34_ssc_1;
  wire Gelu_for_else_else_else_and_5_ssc_1;
  wire Gelu_for_else_and_2_ssc_1;
  wire Gelu_for_else_else_else_and_2_ssc_1;
  wire Gelu_for_else_and_33_ssc_1;
  wire Gelu_for_else_else_else_and_3_ssc_1;
  wire Gelu_for_else_and_ssc_1;
  wire Gelu_for_else_else_else_and_ssc_1;
  wire Gelu_for_else_and_32_ssc_1;
  wire Gelu_for_else_else_else_and_1_ssc_1;
  wire while_nand_112_ssc_1;
  wire ActUnit_RunInst_switch_lp_and_801_ssc_1;
  wire ActUnit_RunInst_switch_lp_and_545_ssc_1;
  wire ActUnit_RunInst_switch_lp_and_547_ssc_1;
  wire ActUnit_RunInst_switch_lp_and_551_ssc_1;
  wire ActUnit_RunInst_switch_lp_and_553_ssc_1;
  wire ActUnit_RunInst_switch_lp_and_549_ssc_1;
  wire while_nand_96_ssc_1;
  wire ActUnit_RunInst_switch_lp_and_769_ssc_1;
  wire ActUnit_RunInst_switch_lp_and_385_ssc_1;
  wire ActUnit_RunInst_switch_lp_and_387_ssc_1;
  wire ActUnit_RunInst_switch_lp_and_391_ssc_1;
  wire ActUnit_RunInst_switch_lp_and_393_ssc_1;
  wire ActUnit_RunInst_switch_lp_and_389_ssc_1;
  wire while_nand_80_ssc_1;
  wire ActUnit_RunInst_switch_lp_and_737_ssc_1;
  wire ActUnit_RunInst_switch_lp_and_225_ssc_1;
  wire ActUnit_RunInst_switch_lp_and_227_ssc_1;
  wire ActUnit_RunInst_switch_lp_and_231_ssc_1;
  wire ActUnit_RunInst_switch_lp_and_233_ssc_1;
  wire ActUnit_RunInst_switch_lp_and_229_ssc_1;
  wire while_nand_64_ssc_1;
  wire ActUnit_RunInst_switch_lp_and_704_ssc_1;
  wire ActUnit_RunInst_switch_lp_and_65_ssc_1;
  wire ActUnit_RunInst_switch_lp_and_67_ssc_1;
  wire ActUnit_RunInst_switch_lp_and_71_ssc_1;
  wire ActUnit_RunInst_switch_lp_and_73_ssc_1;
  wire ActUnit_RunInst_switch_lp_and_69_ssc_1;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295;
  wire while_nand_ssc_1;
  wire ActUnit_RunLoad_and_ssc_1;
  wire ActUnit_RunLoad_and_1_ssc_1;
  reg act_regs_data_1_15_sva_31;
  reg [4:0] act_regs_data_1_15_sva_30_26;
  reg [21:0] act_regs_data_1_15_sva_21_0;
  reg act_regs_data_2_0_sva_31;
  reg [4:0] act_regs_data_2_0_sva_30_26;
  reg [21:0] act_regs_data_2_0_sva_21_0;
  reg act_regs_data_1_14_sva_31;
  reg [4:0] act_regs_data_1_14_sva_30_26;
  reg [21:0] act_regs_data_1_14_sva_21_0;
  reg act_regs_data_2_1_sva_31;
  reg [4:0] act_regs_data_2_1_sva_30_26;
  reg [21:0] act_regs_data_2_1_sva_21_0;
  reg act_regs_data_1_13_sva_31;
  reg [4:0] act_regs_data_1_13_sva_30_26;
  reg [21:0] act_regs_data_1_13_sva_21_0;
  reg act_regs_data_2_2_sva_31;
  reg [4:0] act_regs_data_2_2_sva_30_26;
  reg [21:0] act_regs_data_2_2_sva_21_0;
  reg act_regs_data_1_12_sva_31;
  reg [4:0] act_regs_data_1_12_sva_30_26;
  reg [21:0] act_regs_data_1_12_sva_21_0;
  reg act_regs_data_2_3_sva_31;
  reg [4:0] act_regs_data_2_3_sva_30_26;
  reg [21:0] act_regs_data_2_3_sva_21_0;
  reg act_regs_data_1_11_sva_31;
  reg [4:0] act_regs_data_1_11_sva_30_26;
  reg [21:0] act_regs_data_1_11_sva_21_0;
  reg act_regs_data_2_4_sva_31;
  reg [4:0] act_regs_data_2_4_sva_30_26;
  reg [21:0] act_regs_data_2_4_sva_21_0;
  reg act_regs_data_1_10_sva_31;
  reg [4:0] act_regs_data_1_10_sva_30_26;
  reg [21:0] act_regs_data_1_10_sva_21_0;
  reg act_regs_data_2_5_sva_31;
  reg [4:0] act_regs_data_2_5_sva_30_26;
  reg [21:0] act_regs_data_2_5_sva_21_0;
  reg act_regs_data_1_9_sva_31;
  reg [4:0] act_regs_data_1_9_sva_30_26;
  reg [21:0] act_regs_data_1_9_sva_21_0;
  reg act_regs_data_2_6_sva_31;
  reg [4:0] act_regs_data_2_6_sva_30_26;
  reg [21:0] act_regs_data_2_6_sva_21_0;
  reg act_regs_data_1_8_sva_31;
  reg [4:0] act_regs_data_1_8_sva_30_26;
  reg [21:0] act_regs_data_1_8_sva_21_0;
  reg act_regs_data_2_7_sva_31;
  reg [4:0] act_regs_data_2_7_sva_30_26;
  reg [21:0] act_regs_data_2_7_sva_21_0;
  reg act_regs_data_1_7_sva_31;
  reg [4:0] act_regs_data_1_7_sva_30_26;
  reg [21:0] act_regs_data_1_7_sva_21_0;
  reg act_regs_data_2_8_sva_31;
  reg [4:0] act_regs_data_2_8_sva_30_26;
  reg [21:0] act_regs_data_2_8_sva_21_0;
  reg act_regs_data_1_6_sva_31;
  reg [4:0] act_regs_data_1_6_sva_30_26;
  reg [21:0] act_regs_data_1_6_sva_21_0;
  reg act_regs_data_2_9_sva_31;
  reg [4:0] act_regs_data_2_9_sva_30_26;
  reg [21:0] act_regs_data_2_9_sva_21_0;
  reg act_regs_data_1_5_sva_31;
  reg [4:0] act_regs_data_1_5_sva_30_26;
  reg [21:0] act_regs_data_1_5_sva_21_0;
  reg act_regs_data_2_10_sva_31;
  reg [4:0] act_regs_data_2_10_sva_30_26;
  reg [21:0] act_regs_data_2_10_sva_21_0;
  reg act_regs_data_1_4_sva_31;
  reg [4:0] act_regs_data_1_4_sva_30_26;
  reg [21:0] act_regs_data_1_4_sva_21_0;
  reg act_regs_data_2_11_sva_31;
  reg [4:0] act_regs_data_2_11_sva_30_26;
  reg [21:0] act_regs_data_2_11_sva_21_0;
  reg act_regs_data_1_3_sva_31;
  reg [4:0] act_regs_data_1_3_sva_30_26;
  reg [21:0] act_regs_data_1_3_sva_21_0;
  reg act_regs_data_2_12_sva_31;
  reg [4:0] act_regs_data_2_12_sva_30_26;
  reg [21:0] act_regs_data_2_12_sva_21_0;
  reg act_regs_data_1_2_sva_31;
  reg [4:0] act_regs_data_1_2_sva_30_26;
  reg [21:0] act_regs_data_1_2_sva_21_0;
  reg act_regs_data_2_13_sva_31;
  reg [4:0] act_regs_data_2_13_sva_30_26;
  reg [21:0] act_regs_data_2_13_sva_21_0;
  reg act_regs_data_1_1_sva_31;
  reg [4:0] act_regs_data_1_1_sva_30_26;
  reg [21:0] act_regs_data_1_1_sva_21_0;
  reg act_regs_data_2_14_sva_31;
  reg [4:0] act_regs_data_2_14_sva_30_26;
  reg [21:0] act_regs_data_2_14_sva_21_0;
  reg act_regs_data_1_0_sva_31;
  reg [4:0] act_regs_data_1_0_sva_30_26;
  reg [21:0] act_regs_data_1_0_sva_21_0;
  reg act_regs_data_2_15_sva_31;
  reg [4:0] act_regs_data_2_15_sva_30_26;
  reg [21:0] act_regs_data_2_15_sva_21_0;
  reg act_regs_data_0_15_sva_31;
  reg [4:0] act_regs_data_0_15_sva_30_26;
  reg [21:0] act_regs_data_0_15_sva_21_0;
  reg act_regs_data_3_0_sva_31;
  reg [4:0] act_regs_data_3_0_sva_30_26;
  reg [21:0] act_regs_data_3_0_sva_21_0;
  reg act_regs_data_0_14_sva_31;
  reg [4:0] act_regs_data_0_14_sva_30_26;
  reg [21:0] act_regs_data_0_14_sva_21_0;
  reg act_regs_data_3_1_sva_31;
  reg [4:0] act_regs_data_3_1_sva_30_26;
  reg [21:0] act_regs_data_3_1_sva_21_0;
  reg act_regs_data_3_2_sva_31;
  reg [4:0] act_regs_data_3_2_sva_30_26;
  reg [21:0] act_regs_data_3_2_sva_21_0;
  reg act_regs_data_3_3_sva_31;
  reg [4:0] act_regs_data_3_3_sva_30_26;
  reg [21:0] act_regs_data_3_3_sva_21_0;
  reg act_regs_data_3_4_sva_31;
  reg [4:0] act_regs_data_3_4_sva_30_26;
  reg [21:0] act_regs_data_3_4_sva_21_0;
  reg act_regs_data_3_5_sva_31;
  reg [4:0] act_regs_data_3_5_sva_30_26;
  reg [21:0] act_regs_data_3_5_sva_21_0;
  reg act_regs_data_0_9_sva_31;
  reg [4:0] act_regs_data_0_9_sva_30_26;
  reg [21:0] act_regs_data_0_9_sva_21_0;
  reg act_regs_data_3_6_sva_31;
  reg [4:0] act_regs_data_3_6_sva_30_26;
  reg [21:0] act_regs_data_3_6_sva_21_0;
  reg act_regs_data_0_8_sva_31;
  reg [4:0] act_regs_data_0_8_sva_30_26;
  reg [21:0] act_regs_data_0_8_sva_21_0;
  reg act_regs_data_3_7_sva_31;
  reg [4:0] act_regs_data_3_7_sva_30_26;
  reg [21:0] act_regs_data_3_7_sva_21_0;
  reg act_regs_data_0_7_sva_31;
  reg [4:0] act_regs_data_0_7_sva_30_26;
  reg [21:0] act_regs_data_0_7_sva_21_0;
  reg act_regs_data_3_8_sva_31;
  reg [4:0] act_regs_data_3_8_sva_30_26;
  reg [21:0] act_regs_data_3_8_sva_21_0;
  reg act_regs_data_0_6_sva_31;
  reg [4:0] act_regs_data_0_6_sva_30_26;
  reg [21:0] act_regs_data_0_6_sva_21_0;
  reg act_regs_data_3_9_sva_31;
  reg [4:0] act_regs_data_3_9_sva_30_26;
  reg [21:0] act_regs_data_3_9_sva_21_0;
  reg act_regs_data_0_5_sva_31;
  reg [4:0] act_regs_data_0_5_sva_30_26;
  reg [21:0] act_regs_data_0_5_sva_21_0;
  reg act_regs_data_3_10_sva_31;
  reg [4:0] act_regs_data_3_10_sva_30_26;
  reg [21:0] act_regs_data_3_10_sva_21_0;
  reg act_regs_data_0_4_sva_31;
  reg [4:0] act_regs_data_0_4_sva_30_26;
  reg [21:0] act_regs_data_0_4_sva_21_0;
  reg act_regs_data_3_11_sva_31;
  reg [4:0] act_regs_data_3_11_sva_30_26;
  reg [21:0] act_regs_data_3_11_sva_21_0;
  reg act_regs_data_0_3_sva_31;
  reg [4:0] act_regs_data_0_3_sva_30_26;
  reg [21:0] act_regs_data_0_3_sva_21_0;
  reg act_regs_data_3_12_sva_31;
  reg [4:0] act_regs_data_3_12_sva_30_26;
  reg [21:0] act_regs_data_3_12_sva_21_0;
  reg act_regs_data_0_2_sva_31;
  reg [4:0] act_regs_data_0_2_sva_30_26;
  reg [21:0] act_regs_data_0_2_sva_21_0;
  reg act_regs_data_3_13_sva_31;
  reg [4:0] act_regs_data_3_13_sva_30_26;
  reg [21:0] act_regs_data_3_13_sva_21_0;
  reg act_regs_data_3_14_sva_31;
  reg [4:0] act_regs_data_3_14_sva_30_26;
  reg [21:0] act_regs_data_3_14_sva_21_0;
  reg act_regs_data_3_15_sva_31;
  reg [4:0] act_regs_data_3_15_sva_30_26;
  reg [21:0] act_regs_data_3_15_sva_21_0;
  reg [2:0] rva_out_reg_data_71_64_sva_dfm_6_7_5;
  reg [3:0] rva_out_reg_data_39_32_sva_dfm_6_7_4;
  reg [1:0] rva_out_reg_data_29_24_sva_dfm_6_5_4;
  reg [2:0] Silu_for_2_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_24_22;
  reg [2:0] Silu_for_3_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_24_22;
  reg [2:0] Silu_for_4_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_24_22;
  reg [2:0] Silu_for_5_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_24_22;
  reg [2:0] Silu_for_6_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_24_22;
  reg [2:0] Silu_for_7_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_24_22;
  reg [2:0] Silu_for_9_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_24_22;
  reg [2:0] Silu_for_y_1_sva_3_24_22;
  reg [2:0] Silu_for_y_8_sva_3_24_22;
  wire ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_31;
  wire [4:0] ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_30_26;
  wire [21:0] ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_21_0;
  reg act_write_data_data_0_7_sva_31;
  reg act_write_data_data_0_8_sva_31;
  reg act_write_data_data_0_6_sva_31;
  reg act_write_data_data_0_9_sva_31;
  reg act_write_data_data_0_5_sva_31;
  reg act_write_data_data_0_10_sva_31;
  reg act_write_data_data_0_4_sva_31;
  reg act_write_data_data_0_11_sva_31;
  reg act_write_data_data_0_3_sva_31;
  reg act_write_data_data_0_12_sva_31;
  reg act_write_data_data_0_2_sva_31;
  reg act_write_data_data_0_13_sva_31;
  reg act_write_data_data_0_1_sva_31;
  reg act_write_data_data_0_14_sva_31;
  reg act_write_data_data_0_0_sva_31;
  reg act_write_data_data_0_15_sva_2_31;
  wire Tanh_for_and_79_ssc;
  wire Tanh_for_and_77_ssc;
  wire Tanh_for_and_75_ssc;
  wire Tanh_for_and_73_ssc;
  wire Tanh_for_and_71_ssc;
  wire Tanh_for_and_69_ssc;
  wire Tanh_for_and_67_ssc;
  wire Tanh_for_and_65_ssc;
  wire Tanh_for_and_63_ssc;
  wire Tanh_for_and_61_ssc;
  wire Tanh_for_and_59_ssc;
  wire Tanh_for_and_57_ssc;
  wire Tanh_for_and_55_ssc;
  wire Tanh_for_and_53_ssc;
  wire Tanh_for_and_51_ssc;
  wire Tanh_for_and_49_ssc;
  wire ActUnit_PushOutput_if_for_and_28_cse;
  wire act_write_data_data_and_15_cse;
  wire ActUnit_RunInst_switch_lp_and_811_cse;
  wire ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_31_3;
  wire act_write_data_data_act_write_data_data_and_26_cse;
  wire Silu_for_else_else_else_if_or_14_cse;
  wire Silu_for_else_else_else_if_or_13_rgt;
  reg [2:0] rva_out_reg_data_71_64_sva_dfm_3_7_5;
  reg [4:0] rva_out_reg_data_71_64_sva_dfm_3_4_0;
  reg [3:0] rva_out_reg_data_39_32_sva_dfm_3_7_4;
  reg [1:0] rva_out_reg_data_29_24_sva_dfm_3_5_4;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31;
  reg [4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26;
  reg [21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0;
  reg [21:0] Tanh_for_y_25_0_1_lpi_1_dfm_1_21_0;
  reg [4:0] Relu_for_y_qr_30_0_1_lpi_1_dfm_30_26;
  reg [21:0] Relu_for_y_qr_30_0_1_lpi_1_dfm_21_0;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31;
  reg [4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26;
  reg [21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0;
  reg [21:0] Tanh_for_y_25_0_2_lpi_1_dfm_1_21_0;
  reg [4:0] Relu_for_y_qr_30_0_2_lpi_1_dfm_30_26;
  reg [21:0] Relu_for_y_qr_30_0_2_lpi_1_dfm_21_0;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31;
  reg [4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26;
  reg [21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0;
  reg [21:0] Tanh_for_y_25_0_3_lpi_1_dfm_1_21_0;
  reg [4:0] Relu_for_y_qr_30_0_3_lpi_1_dfm_30_26;
  reg [21:0] Relu_for_y_qr_30_0_3_lpi_1_dfm_21_0;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31;
  reg [4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26;
  reg [21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0;
  reg [21:0] Tanh_for_y_25_0_4_lpi_1_dfm_1_21_0;
  reg [4:0] Relu_for_y_qr_30_0_4_lpi_1_dfm_30_26;
  reg [21:0] Relu_for_y_qr_30_0_4_lpi_1_dfm_21_0;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31;
  reg [4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26;
  reg [21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0;
  reg [21:0] Tanh_for_y_25_0_5_lpi_1_dfm_1_21_0;
  reg [4:0] Relu_for_y_qr_30_0_5_lpi_1_dfm_30_26;
  reg [21:0] Relu_for_y_qr_30_0_5_lpi_1_dfm_21_0;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31;
  reg [4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26;
  reg [21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0;
  reg [21:0] Tanh_for_y_25_0_6_lpi_1_dfm_1_21_0;
  reg [4:0] Relu_for_y_qr_30_0_6_lpi_1_dfm_30_26;
  reg [21:0] Relu_for_y_qr_30_0_6_lpi_1_dfm_21_0;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31;
  reg [4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26;
  reg [21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0;
  reg [21:0] Tanh_for_y_25_0_7_lpi_1_dfm_1_21_0;
  reg [4:0] Relu_for_y_qr_30_0_7_lpi_1_dfm_30_26;
  reg [21:0] Relu_for_y_qr_30_0_7_lpi_1_dfm_21_0;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31;
  reg [4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26;
  reg [21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0;
  reg [21:0] Tanh_for_y_25_0_8_lpi_1_dfm_1_21_0;
  reg [4:0] Relu_for_y_qr_30_0_8_lpi_1_dfm_30_26;
  reg [21:0] Relu_for_y_qr_30_0_8_lpi_1_dfm_21_0;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31;
  reg [4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26;
  reg [21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0;
  reg [21:0] Tanh_for_y_25_0_9_lpi_1_dfm_1_21_0;
  reg [4:0] Relu_for_y_qr_30_0_9_lpi_1_dfm_30_26;
  reg [21:0] Relu_for_y_qr_30_0_9_lpi_1_dfm_21_0;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31;
  reg [4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26;
  reg [21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0;
  reg [21:0] Tanh_for_y_25_0_10_lpi_1_dfm_1_21_0;
  reg [4:0] Relu_for_y_qr_30_0_10_lpi_1_dfm_30_26;
  reg [21:0] Relu_for_y_qr_30_0_10_lpi_1_dfm_21_0;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31;
  reg [4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26;
  reg [21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0;
  reg [21:0] Tanh_for_y_25_0_11_lpi_1_dfm_1_21_0;
  reg [4:0] Relu_for_y_qr_30_0_11_lpi_1_dfm_30_26;
  reg [21:0] Relu_for_y_qr_30_0_11_lpi_1_dfm_21_0;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31;
  reg [4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26;
  reg [21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0;
  reg [21:0] Tanh_for_y_25_0_12_lpi_1_dfm_1_21_0;
  reg [4:0] Relu_for_y_qr_30_0_12_lpi_1_dfm_30_26;
  reg [21:0] Relu_for_y_qr_30_0_12_lpi_1_dfm_21_0;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31;
  reg [4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26;
  reg [21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0;
  reg [21:0] Tanh_for_y_25_0_13_lpi_1_dfm_1_21_0;
  reg [4:0] Relu_for_y_qr_30_0_13_lpi_1_dfm_30_26;
  reg [21:0] Relu_for_y_qr_30_0_13_lpi_1_dfm_21_0;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31;
  reg [4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26;
  reg [21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0;
  reg [21:0] Tanh_for_y_25_0_14_lpi_1_dfm_1_21_0;
  reg [4:0] Relu_for_y_qr_30_0_14_lpi_1_dfm_30_26;
  reg [21:0] Relu_for_y_qr_30_0_14_lpi_1_dfm_21_0;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31;
  reg [4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26;
  reg [21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0;
  reg [21:0] Tanh_for_y_25_0_15_lpi_1_dfm_1_21_0;
  reg [4:0] Relu_for_y_qr_30_0_15_lpi_1_dfm_30_26;
  reg [21:0] Relu_for_y_qr_30_0_15_lpi_1_dfm_21_0;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31;
  reg [4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26;
  reg [21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0;
  wire Tanh_for_y_and_ssc;
  reg [21:0] Tanh_for_y_25_0_lpi_1_dfm_1_21_0;
  wire Relu_for_y_qelse_and_ssc;
  reg [4:0] Relu_for_y_qr_30_0_lpi_1_dfm_30_26;
  reg [21:0] Relu_for_y_qr_30_0_lpi_1_dfm_21_0;
  reg [4:0] act_write_data_data_0_7_sva_30_26;
  reg [21:0] act_write_data_data_0_7_sva_21_0;
  reg [4:0] act_write_data_data_0_8_sva_30_26;
  reg [21:0] act_write_data_data_0_8_sva_21_0;
  reg [4:0] act_write_data_data_0_6_sva_30_26;
  reg [21:0] act_write_data_data_0_6_sva_21_0;
  reg [4:0] act_write_data_data_0_9_sva_30_26;
  reg [21:0] act_write_data_data_0_9_sva_21_0;
  reg [4:0] act_write_data_data_0_5_sva_30_26;
  reg [21:0] act_write_data_data_0_5_sva_21_0;
  reg [4:0] act_write_data_data_0_10_sva_30_26;
  reg [21:0] act_write_data_data_0_10_sva_21_0;
  reg [4:0] act_write_data_data_0_4_sva_30_26;
  reg [21:0] act_write_data_data_0_4_sva_21_0;
  reg [4:0] act_write_data_data_0_11_sva_30_26;
  reg [21:0] act_write_data_data_0_11_sva_21_0;
  reg [4:0] act_write_data_data_0_3_sva_30_26;
  reg [21:0] act_write_data_data_0_3_sva_21_0;
  reg [4:0] act_write_data_data_0_12_sva_30_26;
  reg [21:0] act_write_data_data_0_12_sva_21_0;
  reg [4:0] act_write_data_data_0_2_sva_30_26;
  reg [21:0] act_write_data_data_0_2_sva_21_0;
  reg [4:0] act_write_data_data_0_13_sva_30_26;
  reg [21:0] act_write_data_data_0_13_sva_21_0;
  reg [4:0] act_write_data_data_0_1_sva_30_26;
  reg [21:0] act_write_data_data_0_1_sva_21_0;
  reg [4:0] act_write_data_data_0_14_sva_30_26;
  reg [21:0] act_write_data_data_0_14_sva_21_0;
  wire act_write_data_data_and_16_ssc;
  reg [4:0] act_write_data_data_0_0_sva_30_26;
  reg [21:0] act_write_data_data_0_0_sva_21_0;
  reg [4:0] act_write_data_data_0_15_sva_2_30_26;
  reg [21:0] act_write_data_data_0_15_sva_2_21_0;
  reg [21:0] reg_nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1;
  reg [4:0] reg_nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26;
  reg [21:0] reg_nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1;
  reg [4:0] reg_nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26;
  reg [21:0] reg_nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1;
  reg [4:0] reg_nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26;
  reg [21:0] reg_nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1;
  reg [4:0] reg_nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26;
  reg [21:0] reg_nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1;
  reg [4:0] reg_nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26;
  reg [21:0] reg_nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1;
  reg [4:0] reg_nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26;
  reg [21:0] reg_nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1;
  reg [4:0] reg_nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26;
  reg [21:0] reg_nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1;
  reg [4:0] reg_nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26;
  reg [21:0] reg_nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1;
  reg [4:0] reg_nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26;
  reg [21:0] reg_nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1;
  reg [4:0] reg_nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26;
  reg [21:0] reg_nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1;
  reg [4:0] reg_nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26;
  reg [21:0] reg_nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1;
  reg [4:0] reg_nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26;
  reg [21:0] reg_nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1;
  reg [4:0] reg_nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26;
  reg [21:0] reg_nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1;
  reg [4:0] reg_nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26;
  reg [21:0] reg_nv_scvector_cctor_nv_scvector_5_for_2_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1;
  reg [4:0] reg_nv_scvector_cctor_nv_scvector_5_for_2_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26;
  reg [21:0] reg_ActUnit_RunInst_case_14_nv_scvector_cctor_data_0_1_ftd_1;
  reg [4:0] reg_ActUnit_RunInst_case_14_nv_scvector_cctor_data_0_ftd_1_30_26;
  reg [21:0] reg_ActUnit_RunInst_case_15_nv_scvector_cctor_data_0_ftd_1;
  reg [4:0] ActUnit_RunInst_case_15_nv_scvector_cctor_data_0_sva_30_26;
  reg [21:0] reg_nv_scvector_cctor_nv_scvector_6_for_16_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1;
  reg [4:0] nv_scvector_cctor_nv_scvector_6_for_16_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26;
  reg [21:0] reg_nv_scvector_cctor_nv_scvector_6_for_15_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1;
  reg [4:0] nv_scvector_cctor_nv_scvector_6_for_15_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26;
  reg [21:0] reg_nv_scvector_cctor_nv_scvector_6_for_14_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1;
  reg [4:0] nv_scvector_cctor_nv_scvector_6_for_14_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26;
  reg [21:0] reg_nv_scvector_cctor_nv_scvector_6_for_13_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1;
  reg [4:0] nv_scvector_cctor_nv_scvector_6_for_13_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26;
  reg [21:0] reg_nv_scvector_cctor_nv_scvector_6_for_12_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1;
  reg [4:0] nv_scvector_cctor_nv_scvector_6_for_12_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26;
  reg [21:0] reg_nv_scvector_cctor_nv_scvector_6_for_11_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1;
  reg [4:0] nv_scvector_cctor_nv_scvector_6_for_11_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26;
  reg [21:0] reg_nv_scvector_cctor_nv_scvector_6_for_10_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1;
  reg [4:0] nv_scvector_cctor_nv_scvector_6_for_10_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26;
  reg [21:0] reg_nv_scvector_cctor_nv_scvector_6_for_9_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1;
  reg [4:0] nv_scvector_cctor_nv_scvector_6_for_9_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26;
  reg [21:0] reg_nv_scvector_cctor_nv_scvector_6_for_8_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1;
  reg [4:0] nv_scvector_cctor_nv_scvector_6_for_8_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26;
  reg [21:0] reg_nv_scvector_cctor_nv_scvector_6_for_7_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1;
  reg [4:0] nv_scvector_cctor_nv_scvector_6_for_7_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26;
  reg [21:0] reg_nv_scvector_cctor_nv_scvector_6_for_6_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1;
  reg [4:0] nv_scvector_cctor_nv_scvector_6_for_6_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26;
  reg [21:0] reg_nv_scvector_cctor_nv_scvector_6_for_5_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1;
  reg [4:0] nv_scvector_cctor_nv_scvector_6_for_5_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26;
  reg [21:0] reg_nv_scvector_cctor_nv_scvector_6_for_4_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1;
  reg [4:0] nv_scvector_cctor_nv_scvector_6_for_4_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26;
  reg [21:0] reg_nv_scvector_cctor_nv_scvector_6_for_3_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1;
  reg [4:0] nv_scvector_cctor_nv_scvector_6_for_3_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26;
  reg [21:0] reg_nv_scvector_cctor_nv_scvector_6_for_2_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1;
  reg [4:0] nv_scvector_cctor_nv_scvector_6_for_2_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26;
  wire [4:0] Gelu_for_y_1_lpi_1_dfm_4_30_26;
  wire [4:0] Gelu_for_y_2_lpi_1_dfm_4_30_26;
  wire [4:0] Gelu_for_y_3_lpi_1_dfm_4_30_26;
  wire [4:0] Gelu_for_y_4_lpi_1_dfm_4_30_26;
  wire [4:0] Gelu_for_y_5_lpi_1_dfm_4_30_26;
  wire [4:0] Gelu_for_y_6_lpi_1_dfm_4_30_26;
  wire [4:0] Gelu_for_y_7_lpi_1_dfm_4_30_26;
  wire [4:0] Gelu_for_y_8_lpi_1_dfm_4_30_26;
  wire [4:0] Gelu_for_y_9_lpi_1_dfm_4_30_26;
  wire [4:0] Gelu_for_y_10_lpi_1_dfm_4_30_26;
  wire [4:0] Gelu_for_y_11_lpi_1_dfm_4_30_26;
  wire [4:0] Gelu_for_y_12_lpi_1_dfm_4_30_26;
  wire [4:0] Gelu_for_y_13_lpi_1_dfm_4_30_26;
  wire [4:0] Gelu_for_y_14_lpi_1_dfm_4_30_26;
  wire [4:0] Gelu_for_y_15_lpi_1_dfm_4_30_26;
  wire [4:0] Gelu_for_y_lpi_1_dfm_4_30_26;
  wire act_write_data_data_and_96_cse;
  wire Gelu_for_y_1_lpi_1_dfm_4_25;
  wire [2:0] Gelu_for_y_1_lpi_1_dfm_4_24_22;
  wire Gelu_for_y_2_lpi_1_dfm_4_25;
  wire [2:0] Gelu_for_y_2_lpi_1_dfm_4_24_22;
  wire Gelu_for_y_3_lpi_1_dfm_4_25;
  wire [2:0] Gelu_for_y_3_lpi_1_dfm_4_24_22;
  wire Gelu_for_y_4_lpi_1_dfm_4_25;
  wire [2:0] Gelu_for_y_4_lpi_1_dfm_4_24_22;
  wire Gelu_for_y_5_lpi_1_dfm_4_25;
  wire [2:0] Gelu_for_y_5_lpi_1_dfm_4_24_22;
  wire Gelu_for_y_6_lpi_1_dfm_4_25;
  wire [2:0] Gelu_for_y_6_lpi_1_dfm_4_24_22;
  wire Gelu_for_y_7_lpi_1_dfm_4_25;
  wire [2:0] Gelu_for_y_7_lpi_1_dfm_4_24_22;
  wire Gelu_for_y_8_lpi_1_dfm_4_25;
  wire [2:0] Gelu_for_y_8_lpi_1_dfm_4_24_22;
  wire Gelu_for_y_9_lpi_1_dfm_4_25;
  wire [2:0] Gelu_for_y_9_lpi_1_dfm_4_24_22;
  wire Gelu_for_y_10_lpi_1_dfm_4_25;
  wire [2:0] Gelu_for_y_10_lpi_1_dfm_4_24_22;
  wire Gelu_for_y_11_lpi_1_dfm_4_25;
  wire [2:0] Gelu_for_y_11_lpi_1_dfm_4_24_22;
  wire Gelu_for_y_12_lpi_1_dfm_4_25;
  wire [2:0] Gelu_for_y_12_lpi_1_dfm_4_24_22;
  wire Gelu_for_y_13_lpi_1_dfm_4_25;
  wire [2:0] Gelu_for_y_13_lpi_1_dfm_4_24_22;
  wire Gelu_for_y_14_lpi_1_dfm_4_25;
  wire [2:0] Gelu_for_y_14_lpi_1_dfm_4_24_22;
  wire Gelu_for_y_15_lpi_1_dfm_4_25;
  wire [2:0] Gelu_for_y_15_lpi_1_dfm_4_24_22;
  wire Gelu_for_y_lpi_1_dfm_4_25;
  wire [2:0] Gelu_for_y_lpi_1_dfm_4_24_22;
  wire ActUnit_DecodeAxi_if_and_37_cse;
  wire act_config_inst_regs_and_36_cse;
  wire operator_32_8_true_AC_TRN_AC_WRAP_2_and_16_cse;
  wire operator_32_8_true_AC_TRN_AC_WRAP_and_cse;
  wire operator_32_8_true_AC_TRN_AC_WRAP_and_23_cse;
  wire Gelu_for_if_and_cse;
  wire act_mem_banks_read_for_and_cse;
  wire rva_out_reg_data_and_62_cse;
  wire act_regs_data_and_832_cse;
  wire act_regs_data_and_892_cse;
  wire act_regs_data_and_893_cse;
  wire act_regs_data_and_898_cse;
  wire act_regs_data_and_899_cse;
  wire act_regs_data_and_904_cse;
  wire act_regs_data_and_905_cse;
  wire act_regs_data_and_910_cse;
  wire act_regs_data_and_911_cse;
  wire act_regs_data_and_916_cse;
  wire act_regs_data_and_917_cse;
  wire act_regs_data_and_922_cse;
  wire act_regs_data_and_923_cse;
  wire act_regs_data_and_928_cse;
  wire act_regs_data_and_929_cse;
  wire act_regs_data_and_934_cse;
  wire act_regs_data_and_935_cse;
  wire act_regs_data_and_940_cse;
  wire act_regs_data_and_941_cse;
  wire act_regs_data_and_946_cse;
  wire act_regs_data_and_947_cse;
  wire act_regs_data_and_952_cse;
  wire act_regs_data_and_953_cse;
  wire act_regs_data_and_958_cse;
  wire act_regs_data_and_959_cse;
  wire act_regs_data_and_964_cse;
  wire act_regs_data_and_965_cse;
  wire act_regs_data_and_970_cse;
  wire act_regs_data_and_971_cse;
  wire act_regs_data_and_976_cse;
  wire act_regs_data_and_977_cse;
  wire act_regs_data_and_982_cse;
  wire act_regs_data_and_983_cse;
  wire act_regs_data_and_988_cse;
  wire act_regs_data_and_989_cse;
  wire act_regs_data_and_994_cse;
  wire act_regs_data_and_995_cse;
  wire act_regs_data_and_1000_cse;
  wire act_regs_data_and_1001_cse;
  wire act_regs_data_and_1006_cse;
  wire act_regs_data_and_1007_cse;
  wire act_regs_data_and_1012_cse;
  wire act_regs_data_and_1013_cse;
  wire act_regs_data_and_1018_cse;
  wire act_regs_data_and_1019_cse;
  wire act_regs_data_and_1024_cse;
  wire act_regs_data_and_1025_cse;
  wire act_regs_data_and_1030_cse;
  wire act_regs_data_and_1031_cse;
  wire act_regs_data_and_1036_cse;
  wire act_regs_data_and_1037_cse;
  wire act_regs_data_and_1042_cse;
  wire act_regs_data_and_1043_cse;
  wire act_regs_data_and_1048_cse;
  wire act_regs_data_and_1049_cse;
  wire act_regs_data_and_1054_cse;
  wire act_regs_data_and_1055_cse;
  wire act_regs_data_and_1060_cse;
  wire act_regs_data_and_1061_cse;
  wire act_regs_data_and_1066_cse;
  wire act_regs_data_and_1067_cse;
  wire act_regs_data_and_1072_cse;
  wire act_regs_data_and_1073_cse;
  wire act_regs_data_and_1078_cse;
  wire act_regs_data_and_1079_cse;
  wire act_regs_data_and_1084_cse;
  wire act_regs_data_and_1085_cse;
  wire act_regs_data_and_1090_cse;
  wire act_regs_data_and_1091_cse;
  wire act_regs_data_and_1096_cse;
  wire act_regs_data_and_1097_cse;
  wire act_regs_data_and_1102_cse;
  wire act_regs_data_and_1103_cse;
  wire act_regs_data_and_1108_cse;
  wire act_regs_data_and_1109_cse;
  wire act_regs_data_and_1114_cse;
  wire act_regs_data_and_1115_cse;
  wire act_regs_data_and_1120_cse;
  wire act_regs_data_and_1121_cse;
  wire act_regs_data_and_1126_cse;
  wire act_regs_data_and_1127_cse;
  wire act_regs_data_and_1132_cse;
  wire act_regs_data_and_1133_cse;
  wire act_regs_data_and_1138_cse;
  wire act_regs_data_and_1139_cse;
  wire act_regs_data_and_1144_cse;
  wire act_regs_data_and_1145_cse;
  wire act_regs_data_and_1150_cse;
  wire act_regs_data_and_1151_cse;
  wire act_regs_data_and_1156_cse;
  wire act_regs_data_and_1157_cse;
  wire act_regs_data_and_1162_cse;
  wire act_regs_data_and_1163_cse;
  wire act_regs_data_and_1168_cse;
  wire act_regs_data_and_1169_cse;
  wire act_regs_data_and_1174_cse;
  wire act_regs_data_and_1175_cse;
  wire act_regs_data_and_1180_cse;
  wire act_regs_data_and_1181_cse;
  wire Silu_for_y_and_2_cse;
  wire act_regs_data_and_1186_cse;
  wire act_regs_data_and_1187_cse;
  wire act_regs_data_and_1188_cse;
  wire act_regs_data_and_1189_cse;
  wire act_regs_data_and_1190_cse;
  wire act_regs_data_and_1191_cse;
  wire act_regs_data_and_1192_cse;
  wire act_regs_data_and_1298_cse;
  wire act_regs_data_and_1299_cse;
  wire act_regs_data_and_1300_cse;
  wire act_regs_data_and_1301_cse;
  wire act_regs_data_and_1302_cse;
  wire act_regs_data_and_1303_cse;
  wire act_regs_data_and_1304_cse;
  wire act_regs_data_and_1410_cse;
  wire act_regs_data_and_1411_cse;
  wire act_regs_data_and_1412_cse;
  wire act_regs_data_and_1413_cse;
  wire act_regs_data_and_1414_cse;
  wire act_regs_data_and_1415_cse;
  wire act_regs_data_and_1416_cse;
  wire act_regs_data_and_1522_cse;
  wire act_regs_data_and_1523_cse;
  wire act_regs_data_and_1524_cse;
  wire act_regs_data_and_1525_cse;
  wire act_regs_data_and_1526_cse;
  wire act_regs_data_and_1527_cse;
  wire act_regs_data_and_1528_cse;
  wire Silu_for_else_if_and_1_cse;
  wire Silu_for_else_if_and_2_cse;
  wire or_tmp_552;
  wire or_tmp_555;
  wire or_tmp_653;
  wire or_tmp_871;
  wire or_tmp_873;
  wire or_tmp_938;
  wire or_tmp_999;
  wire nand_tmp_41;
  wire or_tmp_1057;
  wire or_tmp_1113;
  wire or_tmp_1178;
  wire nand_tmp_73;
  wire or_tmp_1297;
  wire nand_tmp_104;
  wire or_tmp_1408;
  wire nor_tmp_635;
  wire nand_tmp_120;
  wire or_tmp_1529;
  wire nand_tmp_136;
  wire or_tmp_1648;
  wire nor_tmp_771;
  wire nand_tmp_152;
  wire or_tmp_1769;
  wire not_tmp_2198;
  wire nor_1405_cse;
  wire and_1809_cse;
  wire and_1821_cse;
  wire nor_1484_cse;
  wire or_3396_cse;
  wire nor_1479_cse;
  wire or_1702_cse;
  wire or_1714_cse;
  wire and_2344_cse;
  wire or_1726_cse;
  wire or_1738_cse;
  wire or_1750_cse;
  wire or_1762_cse;
  wire or_1798_cse;
  wire or_1810_cse;
  wire and_2350_cse;
  wire or_3395_cse;
  wire or_1831_cse;
  wire nand_533_cse;
  wire mux_746_cse;
  wire nand_cse;
  wire and_2367_cse;
  wire and_2372_cse;
  wire and_2354_cse;
  wire nand_542_cse;
  wire and_2412_cse;
  wire and_2484_cse;
  wire and_2494_cse;
  wire or_1905_cse;
  wire or_1913_cse;
  wire or_1921_cse;
  wire or_1929_cse;
  wire or_1937_cse;
  wire or_1945_cse;
  wire or_1953_cse;
  wire or_1961_cse;
  wire or_1969_cse;
  wire or_1977_cse;
  wire or_1985_cse;
  wire or_1993_cse;
  wire or_2001_cse;
  wire or_2009_cse;
  wire or_2017_cse;
  wire or_2025_cse;
  wire or_2033_cse;
  wire or_2040_cse;
  wire or_2047_cse;
  wire or_2054_cse;
  wire or_2061_cse;
  wire or_2068_cse;
  wire or_2075_cse;
  wire or_2082_cse;
  wire or_2089_cse;
  wire or_2096_cse;
  wire or_2103_cse;
  wire or_2110_cse;
  wire or_2117_cse;
  wire or_2124_cse;
  wire or_2131_cse;
  wire or_2138_cse;
  wire or_2145_cse;
  wire or_2153_cse;
  wire or_2161_cse;
  wire or_2169_cse;
  wire or_2177_cse;
  wire or_2185_cse;
  wire or_2193_cse;
  wire or_2201_cse;
  wire or_2209_cse;
  wire or_2217_cse;
  wire or_2225_cse;
  wire or_2233_cse;
  wire or_2241_cse;
  wire or_2249_cse;
  wire or_2257_cse;
  wire and_2497_cse;
  wire or_2265_cse;
  wire or_2273_cse;
  wire or_2280_cse;
  wire or_2287_cse;
  wire or_2294_cse;
  wire or_2301_cse;
  wire or_2308_cse;
  wire or_2315_cse;
  wire nand_685_cse;
  wire or_2329_cse;
  wire or_2336_cse;
  wire or_2343_cse;
  wire or_2350_cse;
  wire or_2357_cse;
  wire or_2364_cse;
  wire or_2371_cse;
  wire and_2533_cse;
  wire nor_1441_cse;
  wire or_1872_cse;
  wire and_2371_cse;
  wire nor_1553_cse;
  wire nor_320_cse;
  wire or_1579_cse;
  wire nor_1406_cse;
  wire and_2824_cse;
  wire and_2825_cse;
  wire and_2936_cse;
  wire and_2937_cse;
  wire and_2872_cse;
  wire and_2984_cse;
  wire and_1824_cse;
  wire and_1827_cse;
  wire and_1830_cse;
  wire and_1833_cse;
  wire and_1836_cse;
  wire and_1839_cse;
  wire and_1842_cse;
  wire and_1845_cse;
  wire and_1848_cse;
  wire and_1851_cse;
  wire and_1854_cse;
  wire and_1857_cse;
  wire and_1860_cse;
  wire and_2364_cse;
  wire mux_438_cse;
  wire mux_827_cse;
  wire nor_1562_cse;
  wire mux_939_cse;
  wire nor_1578_cse;
  wire nor_1654_cse;
  wire nand_583_cse;
  wire nand_663_cse;
  wire mux_771_cse;
  wire nor_1554_cse;
  wire mux_883_cse;
  wire nor_1570_cse;
  wire mux_995_cse;
  wire nor_1586_cse;
  wire mux_1052_cse;
  wire nor_1594_cse;
  wire mux_1123_cse;
  wire nor_1602_cse;
  wire mux_1180_cse;
  wire nor_1610_cse;
  wire nand_543_cse;
  wire nand_623_cse;
  wire nand_704_cse;
  wire nand_744_cse;
  wire nand_784_cse;
  wire nand_824_cse;
  wire and_1935_cse;
  wire and_1937_cse;
  wire and_1939_cse;
  wire and_1941_cse;
  wire and_1943_cse;
  wire and_1945_cse;
  wire and_1947_cse;
  wire and_1949_cse;
  wire and_1999_cse;
  wire and_2001_cse;
  wire and_2003_cse;
  wire and_2005_cse;
  wire and_2007_cse;
  wire and_2009_cse;
  wire and_2011_cse;
  wire and_2013_cse;
  wire and_1951_cse;
  wire and_1953_cse;
  wire and_1955_cse;
  wire and_1957_cse;
  wire and_1959_cse;
  wire and_1961_cse;
  wire and_1963_cse;
  wire and_1965_cse;
  wire and_1967_cse;
  wire and_1969_cse;
  wire and_1971_cse;
  wire and_1973_cse;
  wire and_1975_cse;
  wire and_1977_cse;
  wire and_1979_cse;
  wire and_1981_cse;
  wire and_1983_cse;
  wire and_1985_cse;
  wire and_1987_cse;
  wire and_1989_cse;
  wire and_1991_cse;
  wire and_1993_cse;
  wire and_1995_cse;
  wire and_1997_cse;
  wire and_2015_cse;
  wire and_2017_cse;
  wire and_2019_cse;
  wire and_2021_cse;
  wire and_2023_cse;
  wire and_2025_cse;
  wire and_2027_cse;
  wire and_2029_cse;
  wire and_2031_cse;
  wire and_2033_cse;
  wire and_2035_cse;
  wire and_2037_cse;
  wire and_2039_cse;
  wire and_2041_cse;
  wire and_2043_cse;
  wire and_2045_cse;
  wire and_2047_cse;
  wire and_2049_cse;
  wire and_2051_cse;
  wire and_2053_cse;
  wire and_2055_cse;
  wire and_2057_cse;
  wire and_2059_cse;
  wire and_2061_cse;
  wire or_dcpl;
  reg reg_is_start_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo;
  reg reg_act_regs_data_3_15_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo;
  reg reg_act_regs_data_3_15_sva_8_30_26_enexo;
  reg reg_act_regs_data_2_2_sva_8_30_26_enexo;
  reg reg_is_start_enexo_1;
  reg reg_act_regs_data_3_15_sva_dfm_2_25_22_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_1;
  reg reg_w_load_lpi_1_dfm_1_enexo_1;
  reg reg_act_regs_data_3_15_sva_8_25_22_enexo;
  reg reg_act_regs_data_2_2_sva_8_25_22_enexo;
  reg reg_is_start_enexo_2;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_2;
  reg reg_act_regs_data_3_15_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_2;
  reg reg_act_regs_data_3_15_sva_8_21_0_enexo;
  reg reg_act_regs_data_2_2_sva_8_21_0_enexo;
  reg reg_is_start_enexo_3;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_3;
  reg reg_act_regs_data_2_15_sva_8_30_26_enexo;
  reg reg_act_regs_data_3_14_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_3;
  reg reg_act_regs_data_3_14_sva_8_30_26_enexo;
  reg reg_is_start_enexo_4;
  reg reg_act_regs_data_3_14_sva_dfm_2_25_22_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_4;
  reg reg_act_regs_data_2_15_sva_8_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_4;
  reg reg_act_regs_data_3_14_sva_8_25_22_enexo;
  reg reg_is_start_enexo_5;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_5;
  reg reg_act_regs_data_2_15_sva_8_21_0_enexo;
  reg reg_act_regs_data_3_14_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_5;
  reg reg_act_regs_data_3_14_sva_8_21_0_enexo;
  reg reg_is_start_enexo_6;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_6;
  reg reg_act_regs_data_2_14_sva_8_30_26_enexo;
  reg reg_act_regs_data_3_13_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_6;
  reg reg_act_regs_data_3_13_sva_8_30_26_enexo;
  reg reg_is_start_enexo_7;
  reg reg_act_regs_data_3_13_sva_dfm_2_25_22_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_7;
  reg reg_act_regs_data_2_14_sva_8_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_7;
  reg reg_act_regs_data_3_13_sva_8_25_22_enexo;
  reg reg_is_start_enexo_8;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_8;
  reg reg_act_regs_data_2_14_sva_8_21_0_enexo;
  reg reg_act_regs_data_3_13_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_8;
  reg reg_act_regs_data_3_13_sva_8_21_0_enexo;
  reg reg_is_start_enexo_9;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_9;
  reg reg_act_regs_data_2_13_sva_8_30_26_enexo;
  reg reg_act_regs_data_3_12_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_9;
  reg reg_act_regs_data_3_12_sva_8_30_26_enexo;
  reg reg_is_start_enexo_10;
  reg reg_act_regs_data_3_12_sva_dfm_2_25_22_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_10;
  reg reg_act_regs_data_2_13_sva_8_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_10;
  reg reg_act_regs_data_3_12_sva_8_25_22_enexo;
  reg reg_is_start_enexo_11;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_11;
  reg reg_act_regs_data_2_13_sva_8_21_0_enexo;
  reg reg_act_regs_data_3_12_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_11;
  reg reg_act_regs_data_3_12_sva_8_21_0_enexo;
  reg reg_is_start_enexo_12;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_12;
  reg reg_act_regs_data_2_12_sva_8_30_26_enexo;
  reg reg_act_regs_data_3_11_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_12;
  reg reg_act_regs_data_3_11_sva_8_30_26_enexo;
  reg reg_is_start_enexo_13;
  reg reg_act_regs_data_3_11_sva_dfm_2_25_22_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_13;
  reg reg_act_regs_data_2_12_sva_8_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_13;
  reg reg_act_regs_data_3_11_sva_8_25_22_enexo;
  reg reg_is_start_enexo_14;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_14;
  reg reg_act_regs_data_2_12_sva_8_21_0_enexo;
  reg reg_act_regs_data_3_11_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_14;
  reg reg_act_regs_data_3_11_sva_8_21_0_enexo;
  reg reg_is_start_enexo_15;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_15;
  reg reg_act_regs_data_2_11_sva_8_30_26_enexo;
  reg reg_act_regs_data_3_10_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_15;
  reg reg_act_regs_data_3_10_sva_8_30_26_enexo;
  reg reg_is_start_enexo_16;
  reg reg_act_regs_data_3_10_sva_dfm_2_25_22_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_16;
  reg reg_act_regs_data_2_11_sva_8_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_16;
  reg reg_act_regs_data_3_10_sva_8_25_22_enexo;
  reg reg_is_start_enexo_17;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_17;
  reg reg_act_regs_data_2_11_sva_8_21_0_enexo;
  reg reg_act_regs_data_3_10_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_17;
  reg reg_act_regs_data_3_10_sva_8_21_0_enexo;
  reg reg_is_start_enexo_18;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_18;
  reg reg_act_regs_data_3_0_sva_8_30_26_enexo;
  reg reg_act_regs_data_3_9_sva_dfm_2_30_26_enexo;
  reg reg_act_regs_data_3_9_sva_8_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_18;
  reg reg_is_start_enexo_19;
  reg reg_act_regs_data_3_9_sva_dfm_2_25_22_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_19;
  reg reg_act_regs_data_3_0_sva_8_25_22_enexo;
  reg reg_act_regs_data_3_9_sva_8_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_19;
  reg reg_is_start_enexo_20;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_20;
  reg reg_act_regs_data_3_0_sva_8_21_0_enexo;
  reg reg_act_regs_data_3_9_sva_dfm_2_21_0_enexo;
  reg reg_act_regs_data_3_9_sva_8_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_20;
  reg reg_is_start_enexo_21;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_21;
  reg reg_act_regs_data_2_9_sva_8_30_26_enexo;
  reg reg_act_regs_data_3_8_sva_dfm_2_30_26_enexo;
  reg reg_act_regs_data_3_8_sva_8_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_21;
  reg reg_is_start_enexo_22;
  reg reg_act_regs_data_3_8_sva_dfm_2_25_22_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_22;
  reg reg_act_regs_data_2_9_sva_8_25_22_enexo;
  reg reg_act_regs_data_3_8_sva_8_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_22;
  reg reg_is_start_enexo_23;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_23;
  reg reg_act_regs_data_2_9_sva_8_21_0_enexo;
  reg reg_act_regs_data_3_8_sva_dfm_2_21_0_enexo;
  reg reg_act_regs_data_3_8_sva_8_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_23;
  reg reg_is_start_enexo_24;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_24;
  reg reg_act_regs_data_2_8_sva_8_30_26_enexo;
  reg reg_act_regs_data_3_7_sva_dfm_2_30_26_enexo;
  reg reg_act_regs_data_3_7_sva_8_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_24;
  reg reg_is_start_enexo_25;
  reg reg_act_regs_data_3_7_sva_dfm_2_25_22_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_25;
  reg reg_act_regs_data_2_8_sva_8_25_22_enexo;
  reg reg_act_regs_data_3_7_sva_8_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_25;
  reg reg_is_start_enexo_26;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_26;
  reg reg_act_regs_data_2_8_sva_8_21_0_enexo;
  reg reg_act_regs_data_3_7_sva_dfm_2_21_0_enexo;
  reg reg_act_regs_data_3_7_sva_8_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_26;
  reg reg_is_start_enexo_27;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_27;
  reg reg_act_regs_data_2_7_sva_8_30_26_enexo;
  reg reg_act_regs_data_3_6_sva_dfm_2_30_26_enexo;
  reg reg_act_regs_data_3_6_sva_8_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_27;
  reg reg_is_start_enexo_28;
  reg reg_act_regs_data_3_6_sva_dfm_2_25_22_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_28;
  reg reg_act_regs_data_2_7_sva_8_25_22_enexo;
  reg reg_act_regs_data_3_6_sva_8_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_28;
  reg reg_is_start_enexo_29;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_29;
  reg reg_act_regs_data_2_7_sva_8_21_0_enexo;
  reg reg_act_regs_data_3_6_sva_dfm_2_21_0_enexo;
  reg reg_act_regs_data_3_6_sva_8_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_29;
  reg reg_is_start_enexo_30;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_30;
  reg reg_act_regs_data_2_6_sva_8_30_26_enexo;
  reg reg_act_regs_data_3_5_sva_dfm_2_30_26_enexo;
  reg reg_act_regs_data_3_5_sva_8_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_30;
  reg reg_is_start_enexo_31;
  reg reg_act_regs_data_3_5_sva_dfm_2_25_22_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_31;
  reg reg_act_regs_data_2_6_sva_8_25_22_enexo;
  reg reg_act_regs_data_3_5_sva_8_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_31;
  reg reg_is_start_enexo_32;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_32;
  reg reg_act_regs_data_2_6_sva_8_21_0_enexo;
  reg reg_act_regs_data_3_5_sva_dfm_2_21_0_enexo;
  reg reg_act_regs_data_3_5_sva_8_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_32;
  reg reg_is_start_enexo_33;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_33;
  reg reg_act_regs_data_2_5_sva_8_30_26_enexo;
  reg reg_act_regs_data_3_4_sva_dfm_2_30_26_enexo;
  reg reg_act_regs_data_3_4_sva_8_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_33;
  reg reg_is_start_enexo_34;
  reg reg_act_regs_data_3_4_sva_dfm_2_25_22_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_34;
  reg reg_act_regs_data_2_5_sva_8_25_22_enexo;
  reg reg_act_regs_data_3_4_sva_8_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_34;
  reg reg_is_start_enexo_35;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_35;
  reg reg_act_regs_data_3_4_sva_dfm_2_21_0_enexo;
  reg reg_act_regs_data_3_4_sva_8_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_35;
  reg reg_act_regs_data_2_5_sva_8_21_0_enexo;
  reg reg_is_start_enexo_36;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_36;
  reg reg_act_regs_data_3_3_sva_dfm_2_30_26_enexo;
  reg reg_act_regs_data_3_3_sva_8_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_36;
  reg reg_act_regs_data_2_4_sva_8_30_26_enexo;
  reg reg_is_start_enexo_37;
  reg reg_act_regs_data_3_3_sva_dfm_2_25_22_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_37;
  reg reg_act_regs_data_3_3_sva_8_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_37;
  reg reg_act_regs_data_2_4_sva_8_25_22_enexo;
  reg reg_is_start_enexo_38;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_38;
  reg reg_act_regs_data_3_3_sva_dfm_2_21_0_enexo;
  reg reg_act_regs_data_3_3_sva_8_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_38;
  reg reg_act_regs_data_2_4_sva_8_21_0_enexo;
  reg reg_is_start_enexo_39;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_39;
  reg reg_act_regs_data_3_2_sva_dfm_2_30_26_enexo;
  reg reg_act_regs_data_3_2_sva_8_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_39;
  reg reg_act_regs_data_2_3_sva_8_30_26_enexo;
  reg reg_is_start_enexo_40;
  reg reg_act_regs_data_3_2_sva_dfm_2_25_22_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_40;
  reg reg_act_regs_data_3_2_sva_8_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_40;
  reg reg_act_regs_data_2_3_sva_8_25_22_enexo;
  reg reg_is_start_enexo_41;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_41;
  reg reg_act_regs_data_3_2_sva_dfm_2_21_0_enexo;
  reg reg_act_regs_data_3_2_sva_8_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_41;
  reg reg_act_regs_data_2_3_sva_8_21_0_enexo;
  reg reg_is_start_enexo_42;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_42;
  reg reg_act_regs_data_2_10_sva_8_30_26_enexo;
  reg reg_act_regs_data_3_1_sva_dfm_2_30_26_enexo;
  reg reg_act_regs_data_3_1_sva_8_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_42;
  reg reg_is_start_enexo_43;
  reg reg_act_regs_data_3_1_sva_dfm_2_25_22_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_43;
  reg reg_act_regs_data_2_10_sva_8_25_22_enexo;
  reg reg_act_regs_data_3_1_sva_8_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_43;
  reg reg_is_start_enexo_44;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_44;
  reg reg_act_regs_data_2_10_sva_8_21_0_enexo;
  reg reg_act_regs_data_3_1_sva_dfm_2_21_0_enexo;
  reg reg_act_regs_data_3_1_sva_8_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_44;
  reg reg_is_start_enexo_45;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_45;
  reg reg_act_regs_data_3_0_sva_8_30_26_enexo_1;
  reg reg_act_regs_data_3_0_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_45;
  reg reg_act_regs_data_2_1_sva_8_30_26_enexo;
  reg reg_is_start_enexo_46;
  reg reg_act_regs_data_3_0_sva_dfm_2_25_22_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_46;
  reg reg_act_regs_data_3_0_sva_8_25_22_enexo_1;
  reg reg_w_load_lpi_1_dfm_1_enexo_46;
  reg reg_act_regs_data_2_1_sva_8_25_22_enexo;
  reg reg_is_start_enexo_47;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_47;
  reg reg_act_regs_data_3_0_sva_8_21_0_enexo_1;
  reg reg_act_regs_data_3_0_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_47;
  reg reg_act_regs_data_2_1_sva_8_21_0_enexo;
  reg reg_is_start_enexo_48;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_48;
  reg reg_act_regs_data_1_2_sva_8_30_26_enexo;
  reg reg_act_regs_data_2_15_sva_8_30_26_enexo_1;
  reg reg_act_regs_data_2_15_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_48;
  reg reg_is_start_enexo_49;
  reg reg_act_regs_data_2_15_sva_dfm_2_25_22_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_49;
  reg reg_act_regs_data_1_2_sva_8_25_22_enexo;
  reg reg_act_regs_data_2_15_sva_8_25_22_enexo_1;
  reg reg_w_load_lpi_1_dfm_1_enexo_49;
  reg reg_is_start_enexo_50;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_50;
  reg reg_act_regs_data_1_2_sva_8_21_0_enexo;
  reg reg_act_regs_data_2_15_sva_8_21_0_enexo_1;
  reg reg_act_regs_data_2_15_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_50;
  reg reg_is_start_enexo_51;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_51;
  reg reg_act_regs_data_2_14_sva_8_30_26_enexo_1;
  reg reg_act_regs_data_2_14_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_51;
  reg reg_act_regs_data_1_15_sva_8_30_26_enexo;
  reg reg_is_start_enexo_52;
  reg reg_act_regs_data_2_14_sva_dfm_2_25_22_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_52;
  reg reg_act_regs_data_2_14_sva_8_25_22_enexo_1;
  reg reg_w_load_lpi_1_dfm_1_enexo_52;
  reg reg_act_regs_data_1_15_sva_8_25_22_enexo;
  reg reg_is_start_enexo_53;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_53;
  reg reg_act_regs_data_2_14_sva_8_21_0_enexo_1;
  reg reg_act_regs_data_2_14_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_53;
  reg reg_act_regs_data_1_15_sva_8_21_0_enexo;
  reg reg_is_start_enexo_54;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_54;
  reg reg_act_regs_data_2_13_sva_8_30_26_enexo_1;
  reg reg_act_regs_data_2_13_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_54;
  reg reg_act_regs_data_1_14_sva_8_30_26_enexo;
  reg reg_is_start_enexo_55;
  reg reg_act_regs_data_2_13_sva_dfm_2_25_22_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_55;
  reg reg_act_regs_data_2_13_sva_8_25_22_enexo_1;
  reg reg_w_load_lpi_1_dfm_1_enexo_55;
  reg reg_act_regs_data_1_14_sva_8_25_22_enexo;
  reg reg_is_start_enexo_56;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_56;
  reg reg_act_regs_data_2_13_sva_8_21_0_enexo_1;
  reg reg_act_regs_data_2_13_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_56;
  reg reg_act_regs_data_1_14_sva_8_21_0_enexo;
  reg reg_is_start_enexo_57;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_57;
  reg reg_act_regs_data_2_12_sva_8_30_26_enexo_1;
  reg reg_act_regs_data_2_12_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_57;
  reg reg_act_regs_data_1_13_sva_8_30_26_enexo;
  reg reg_is_start_enexo_58;
  reg reg_act_regs_data_2_12_sva_dfm_2_25_22_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_58;
  reg reg_act_regs_data_2_12_sva_8_25_22_enexo_1;
  reg reg_w_load_lpi_1_dfm_1_enexo_58;
  reg reg_act_regs_data_1_13_sva_8_25_22_enexo;
  reg reg_is_start_enexo_59;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_59;
  reg reg_act_regs_data_2_12_sva_8_21_0_enexo_1;
  reg reg_act_regs_data_2_12_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_59;
  reg reg_act_regs_data_1_13_sva_8_21_0_enexo;
  reg reg_is_start_enexo_60;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_60;
  reg reg_act_regs_data_2_11_sva_8_30_26_enexo_1;
  reg reg_act_regs_data_2_11_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_60;
  reg reg_act_regs_data_1_12_sva_8_30_26_enexo;
  reg reg_is_start_enexo_61;
  reg reg_act_regs_data_2_11_sva_dfm_2_25_22_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_61;
  reg reg_act_regs_data_2_11_sva_8_25_22_enexo_1;
  reg reg_w_load_lpi_1_dfm_1_enexo_61;
  reg reg_act_regs_data_1_12_sva_8_25_22_enexo;
  reg reg_is_start_enexo_62;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_62;
  reg reg_act_regs_data_2_11_sva_8_21_0_enexo_1;
  reg reg_act_regs_data_2_11_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_62;
  reg reg_act_regs_data_1_12_sva_8_21_0_enexo;
  reg reg_is_start_enexo_63;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_63;
  reg reg_act_regs_data_2_10_sva_8_30_26_enexo_1;
  reg reg_act_regs_data_2_10_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_63;
  reg reg_act_regs_data_1_11_sva_8_30_26_enexo;
  reg reg_is_start_enexo_64;
  reg reg_act_regs_data_2_10_sva_dfm_2_25_22_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_64;
  reg reg_act_regs_data_2_10_sva_8_25_22_enexo_1;
  reg reg_w_load_lpi_1_dfm_1_enexo_64;
  reg reg_act_regs_data_1_11_sva_8_25_22_enexo;
  reg reg_is_start_enexo_65;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_65;
  reg reg_act_regs_data_2_10_sva_8_21_0_enexo_1;
  reg reg_act_regs_data_2_10_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_65;
  reg reg_act_regs_data_1_11_sva_8_21_0_enexo;
  reg reg_is_start_enexo_66;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_66;
  reg reg_act_regs_data_2_9_sva_8_30_26_enexo_1;
  reg reg_act_regs_data_2_9_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_66;
  reg reg_act_regs_data_2_0_sva_8_30_26_enexo;
  reg reg_is_start_enexo_67;
  reg reg_act_regs_data_2_9_sva_dfm_2_25_22_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_67;
  reg reg_act_regs_data_2_9_sva_8_25_22_enexo_1;
  reg reg_w_load_lpi_1_dfm_1_enexo_67;
  reg reg_act_regs_data_2_0_sva_8_25_22_enexo;
  reg reg_is_start_enexo_68;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_68;
  reg reg_act_regs_data_2_9_sva_8_21_0_enexo_1;
  reg reg_act_regs_data_2_9_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_68;
  reg reg_act_regs_data_2_0_sva_8_21_0_enexo;
  reg reg_is_start_enexo_69;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_69;
  reg reg_act_regs_data_2_8_sva_8_30_26_enexo_1;
  reg reg_act_regs_data_2_8_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_69;
  reg reg_act_regs_data_1_9_sva_8_30_26_enexo;
  reg reg_is_start_enexo_70;
  reg reg_act_regs_data_2_8_sva_dfm_2_25_22_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_70;
  reg reg_act_regs_data_1_9_sva_8_25_22_enexo;
  reg reg_act_regs_data_2_8_sva_8_25_22_enexo_1;
  reg reg_w_load_lpi_1_dfm_1_enexo_70;
  reg reg_is_start_enexo_71;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_71;
  reg reg_act_regs_data_1_9_sva_8_21_0_enexo;
  reg reg_act_regs_data_2_8_sva_8_21_0_enexo_1;
  reg reg_act_regs_data_2_8_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_71;
  reg reg_is_start_enexo_72;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_72;
  reg reg_act_regs_data_1_8_sva_8_30_26_enexo;
  reg reg_act_regs_data_2_7_sva_8_30_26_enexo_1;
  reg reg_act_regs_data_2_7_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_72;
  reg reg_is_start_enexo_73;
  reg reg_act_regs_data_2_7_sva_dfm_2_25_22_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_73;
  reg reg_act_regs_data_1_8_sva_8_25_22_enexo;
  reg reg_act_regs_data_2_7_sva_8_25_22_enexo_1;
  reg reg_w_load_lpi_1_dfm_1_enexo_73;
  reg reg_is_start_enexo_74;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_74;
  reg reg_act_regs_data_1_8_sva_8_21_0_enexo;
  reg reg_act_regs_data_2_7_sva_8_21_0_enexo_1;
  reg reg_act_regs_data_2_7_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_74;
  reg reg_is_start_enexo_75;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_75;
  reg reg_act_regs_data_1_7_sva_8_30_26_enexo;
  reg reg_act_regs_data_2_6_sva_8_30_26_enexo_1;
  reg reg_act_regs_data_2_6_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_75;
  reg reg_is_start_enexo_76;
  reg reg_act_regs_data_2_6_sva_dfm_2_25_22_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_76;
  reg reg_act_regs_data_1_7_sva_8_25_22_enexo;
  reg reg_act_regs_data_2_6_sva_8_25_22_enexo_1;
  reg reg_w_load_lpi_1_dfm_1_enexo_76;
  reg reg_is_start_enexo_77;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_77;
  reg reg_act_regs_data_1_7_sva_8_21_0_enexo;
  reg reg_act_regs_data_2_6_sva_8_21_0_enexo_1;
  reg reg_act_regs_data_2_6_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_77;
  reg reg_is_start_enexo_78;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_78;
  reg reg_act_regs_data_1_6_sva_8_30_26_enexo;
  reg reg_act_regs_data_2_5_sva_8_30_26_enexo_1;
  reg reg_act_regs_data_2_5_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_78;
  reg reg_is_start_enexo_79;
  reg reg_act_regs_data_2_5_sva_dfm_2_25_22_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_79;
  reg reg_act_regs_data_1_6_sva_8_25_22_enexo;
  reg reg_act_regs_data_2_5_sva_8_25_22_enexo_1;
  reg reg_w_load_lpi_1_dfm_1_enexo_79;
  reg reg_is_start_enexo_80;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_80;
  reg reg_act_regs_data_1_6_sva_8_21_0_enexo;
  reg reg_act_regs_data_2_5_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_80;
  reg reg_act_regs_data_2_5_sva_8_21_0_enexo_1;
  reg reg_is_start_enexo_81;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_81;
  reg reg_act_regs_data_1_5_sva_8_30_26_enexo;
  reg reg_act_regs_data_2_4_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_81;
  reg reg_act_regs_data_2_4_sva_8_30_26_enexo_1;
  reg reg_is_start_enexo_82;
  reg reg_act_regs_data_2_4_sva_dfm_2_25_22_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_82;
  reg reg_act_regs_data_1_5_sva_8_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_82;
  reg reg_act_regs_data_2_4_sva_8_25_22_enexo_1;
  reg reg_is_start_enexo_83;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_83;
  reg reg_act_regs_data_1_5_sva_8_21_0_enexo;
  reg reg_act_regs_data_2_4_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_83;
  reg reg_act_regs_data_2_4_sva_8_21_0_enexo_1;
  reg reg_is_start_enexo_84;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_84;
  reg reg_act_regs_data_1_4_sva_8_30_26_enexo;
  reg reg_act_regs_data_2_3_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_84;
  reg reg_act_regs_data_2_3_sva_8_30_26_enexo_1;
  reg reg_is_start_enexo_85;
  reg reg_act_regs_data_2_3_sva_dfm_2_25_22_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_85;
  reg reg_act_regs_data_1_4_sva_8_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_85;
  reg reg_act_regs_data_2_3_sva_8_25_22_enexo_1;
  reg reg_is_start_enexo_86;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_86;
  reg reg_act_regs_data_1_4_sva_8_21_0_enexo;
  reg reg_act_regs_data_2_3_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_86;
  reg reg_act_regs_data_2_3_sva_8_21_0_enexo_1;
  reg reg_is_start_enexo_87;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_87;
  reg reg_act_regs_data_1_3_sva_8_30_26_enexo;
  reg reg_act_regs_data_2_2_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_87;
  reg reg_act_regs_data_2_2_sva_8_30_26_enexo_1;
  reg reg_is_start_enexo_88;
  reg reg_act_regs_data_2_2_sva_dfm_2_25_22_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_88;
  reg reg_act_regs_data_1_3_sva_8_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_88;
  reg reg_act_regs_data_2_2_sva_8_25_22_enexo_1;
  reg reg_is_start_enexo_89;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_89;
  reg reg_act_regs_data_1_3_sva_8_21_0_enexo;
  reg reg_act_regs_data_2_2_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_89;
  reg reg_act_regs_data_2_2_sva_8_21_0_enexo_1;
  reg reg_is_start_enexo_90;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_90;
  reg reg_act_regs_data_2_1_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_90;
  reg reg_act_regs_data_2_1_sva_8_30_26_enexo_1;
  reg reg_act_regs_data_1_10_sva_8_30_26_enexo;
  reg reg_is_start_enexo_91;
  reg reg_act_regs_data_2_1_sva_dfm_2_25_22_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_91;
  reg reg_w_load_lpi_1_dfm_1_enexo_91;
  reg reg_act_regs_data_2_1_sva_8_25_22_enexo_1;
  reg reg_act_regs_data_1_10_sva_8_25_22_enexo;
  reg reg_is_start_enexo_92;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_92;
  reg reg_act_regs_data_2_1_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_92;
  reg reg_act_regs_data_2_1_sva_8_21_0_enexo_1;
  reg reg_act_regs_data_1_10_sva_8_21_0_enexo;
  reg reg_is_start_enexo_93;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_93;
  reg reg_act_regs_data_1_1_sva_8_30_26_enexo;
  reg reg_act_regs_data_2_0_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_93;
  reg reg_act_regs_data_2_0_sva_8_30_26_enexo_1;
  reg reg_is_start_enexo_94;
  reg reg_act_regs_data_2_0_sva_dfm_2_25_22_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_94;
  reg reg_act_regs_data_1_1_sva_8_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_94;
  reg reg_act_regs_data_2_0_sva_8_25_22_enexo_1;
  reg reg_is_start_enexo_95;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_95;
  reg reg_act_regs_data_1_1_sva_8_21_0_enexo;
  reg reg_act_regs_data_2_0_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_95;
  reg reg_act_regs_data_2_0_sva_8_21_0_enexo_1;
  reg reg_is_start_enexo_96;
  reg reg_act_regs_data_0_2_sva_8_30_26_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_96;
  reg reg_act_regs_data_1_15_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_96;
  reg reg_act_regs_data_1_15_sva_8_30_26_enexo_1;
  reg reg_is_start_enexo_97;
  reg reg_act_regs_data_1_15_sva_dfm_2_25_22_enexo;
  reg reg_act_regs_data_0_2_sva_8_25_22_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_97;
  reg reg_w_load_lpi_1_dfm_1_enexo_97;
  reg reg_act_regs_data_1_15_sva_8_25_22_enexo_1;
  reg reg_is_start_enexo_98;
  reg reg_act_regs_data_0_2_sva_8_21_0_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_98;
  reg reg_act_regs_data_1_15_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_98;
  reg reg_act_regs_data_1_15_sva_8_21_0_enexo_1;
  reg reg_is_start_enexo_99;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_99;
  reg reg_act_regs_data_0_15_sva_8_30_26_enexo;
  reg reg_act_regs_data_1_14_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_99;
  reg reg_act_regs_data_1_14_sva_8_30_26_enexo_1;
  reg reg_is_start_enexo_100;
  reg reg_act_regs_data_1_14_sva_dfm_2_25_22_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_100;
  reg reg_act_regs_data_0_15_sva_8_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_100;
  reg reg_act_regs_data_1_14_sva_8_25_22_enexo_1;
  reg reg_is_start_enexo_101;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_101;
  reg reg_act_regs_data_0_15_sva_8_21_0_enexo;
  reg reg_act_regs_data_1_14_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_101;
  reg reg_act_regs_data_1_14_sva_8_21_0_enexo_1;
  reg reg_is_start_enexo_102;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_102;
  reg reg_act_regs_data_0_14_sva_8_30_26_enexo;
  reg reg_act_regs_data_1_13_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_102;
  reg reg_act_regs_data_1_13_sva_8_30_26_enexo_1;
  reg reg_is_start_enexo_103;
  reg reg_act_regs_data_1_13_sva_dfm_2_25_22_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_103;
  reg reg_act_regs_data_0_14_sva_8_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_103;
  reg reg_act_regs_data_1_13_sva_8_25_22_enexo_1;
  reg reg_is_start_enexo_104;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_104;
  reg reg_act_regs_data_0_14_sva_8_21_0_enexo;
  reg reg_act_regs_data_1_13_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_104;
  reg reg_act_regs_data_1_13_sva_8_21_0_enexo_1;
  reg reg_is_start_enexo_105;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_105;
  reg reg_act_regs_data_0_13_sva_8_30_26_enexo;
  reg reg_act_regs_data_1_12_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_105;
  reg reg_act_regs_data_1_12_sva_8_30_26_enexo_1;
  reg reg_is_start_enexo_106;
  reg reg_act_regs_data_1_12_sva_dfm_2_25_22_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_106;
  reg reg_act_regs_data_0_13_sva_8_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_106;
  reg reg_act_regs_data_1_12_sva_8_25_22_enexo_1;
  reg reg_is_start_enexo_107;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_107;
  reg reg_act_regs_data_0_13_sva_8_21_0_enexo;
  reg reg_act_regs_data_1_12_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_107;
  reg reg_act_regs_data_1_12_sva_8_21_0_enexo_1;
  reg reg_is_start_enexo_108;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_108;
  reg reg_act_regs_data_0_12_sva_8_30_26_enexo;
  reg reg_act_regs_data_1_11_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_108;
  reg reg_act_regs_data_1_11_sva_8_30_26_enexo_1;
  reg reg_is_start_enexo_109;
  reg reg_act_regs_data_1_11_sva_dfm_2_25_22_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_109;
  reg reg_act_regs_data_0_12_sva_8_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_109;
  reg reg_act_regs_data_1_11_sva_8_25_22_enexo_1;
  reg reg_is_start_enexo_110;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_110;
  reg reg_act_regs_data_0_12_sva_8_21_0_enexo;
  reg reg_act_regs_data_1_11_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_110;
  reg reg_act_regs_data_1_11_sva_8_21_0_enexo_1;
  reg reg_is_start_enexo_111;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_111;
  reg reg_act_regs_data_0_11_sva_8_30_26_enexo;
  reg reg_act_regs_data_1_10_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_111;
  reg reg_act_regs_data_1_10_sva_8_30_26_enexo_1;
  reg reg_is_start_enexo_112;
  reg reg_act_regs_data_1_10_sva_dfm_2_25_22_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_112;
  reg reg_act_regs_data_0_11_sva_8_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_112;
  reg reg_act_regs_data_1_10_sva_8_25_22_enexo_1;
  reg reg_is_start_enexo_113;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_113;
  reg reg_act_regs_data_0_11_sva_8_21_0_enexo;
  reg reg_act_regs_data_1_10_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_113;
  reg reg_act_regs_data_1_10_sva_8_21_0_enexo_1;
  reg reg_is_start_enexo_114;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_114;
  reg reg_act_regs_data_1_0_sva_8_30_26_enexo;
  reg reg_act_regs_data_1_9_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_114;
  reg reg_act_regs_data_1_9_sva_8_30_26_enexo_1;
  reg reg_is_start_enexo_115;
  reg reg_act_regs_data_1_9_sva_dfm_2_25_22_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_115;
  reg reg_act_regs_data_1_9_sva_8_25_22_enexo_1;
  reg reg_act_regs_data_1_0_sva_8_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_115;
  reg reg_is_start_enexo_116;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_116;
  reg reg_act_regs_data_1_9_sva_8_21_0_enexo_1;
  reg reg_act_regs_data_1_0_sva_8_21_0_enexo;
  reg reg_act_regs_data_1_9_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_116;
  reg reg_is_start_enexo_117;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_117;
  reg reg_act_regs_data_1_8_sva_8_30_26_enexo_1;
  reg reg_act_regs_data_0_9_sva_8_30_26_enexo;
  reg reg_act_regs_data_1_8_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_117;
  reg reg_is_start_enexo_118;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_118;
  reg reg_act_regs_data_1_8_sva_8_25_22_enexo_1;
  reg reg_act_regs_data_0_9_sva_8_25_22_enexo;
  reg reg_act_regs_data_1_8_sva_dfm_2_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_118;
  reg reg_is_start_enexo_119;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_119;
  reg reg_act_regs_data_1_8_sva_8_21_0_enexo_1;
  reg reg_act_regs_data_0_9_sva_8_21_0_enexo;
  reg reg_act_regs_data_1_8_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_119;
  reg reg_is_start_enexo_120;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_120;
  reg reg_act_regs_data_1_7_sva_8_30_26_enexo_1;
  reg reg_act_regs_data_0_8_sva_8_30_26_enexo;
  reg reg_act_regs_data_1_7_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_120;
  reg reg_is_start_enexo_121;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_121;
  reg reg_act_regs_data_1_7_sva_8_25_22_enexo_1;
  reg reg_act_regs_data_0_8_sva_8_25_22_enexo;
  reg reg_act_regs_data_1_7_sva_dfm_2_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_121;
  reg reg_is_start_enexo_122;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_122;
  reg reg_act_regs_data_1_7_sva_8_21_0_enexo_1;
  reg reg_act_regs_data_0_8_sva_8_21_0_enexo;
  reg reg_act_regs_data_1_7_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_122;
  reg reg_is_start_enexo_123;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_123;
  reg reg_act_regs_data_1_6_sva_8_30_26_enexo_1;
  reg reg_act_regs_data_0_7_sva_8_30_26_enexo;
  reg reg_act_regs_data_1_6_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_123;
  reg reg_is_start_enexo_124;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_124;
  reg reg_act_regs_data_1_6_sva_8_25_22_enexo_1;
  reg reg_act_regs_data_0_7_sva_8_25_22_enexo;
  reg reg_act_regs_data_1_6_sva_dfm_2_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_124;
  reg reg_is_start_enexo_125;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_125;
  reg reg_act_regs_data_1_6_sva_8_21_0_enexo_1;
  reg reg_act_regs_data_0_7_sva_8_21_0_enexo;
  reg reg_act_regs_data_1_6_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_125;
  reg reg_is_start_enexo_126;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_126;
  reg reg_act_regs_data_1_5_sva_8_30_26_enexo_1;
  reg reg_act_regs_data_0_6_sva_8_30_26_enexo;
  reg reg_act_regs_data_1_5_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_126;
  reg reg_is_start_enexo_127;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_127;
  reg reg_act_regs_data_1_5_sva_8_25_22_enexo_1;
  reg reg_act_regs_data_0_6_sva_8_25_22_enexo;
  reg reg_act_regs_data_1_5_sva_dfm_2_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_127;
  reg reg_is_start_enexo_128;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_128;
  reg reg_act_regs_data_1_5_sva_8_21_0_enexo_1;
  reg reg_act_regs_data_0_6_sva_8_21_0_enexo;
  reg reg_act_regs_data_1_5_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_128;
  reg reg_is_start_enexo_129;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_129;
  reg reg_act_regs_data_1_4_sva_8_30_26_enexo_1;
  reg reg_act_regs_data_0_5_sva_8_30_26_enexo;
  reg reg_act_regs_data_1_4_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_129;
  reg reg_is_start_enexo_130;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_130;
  reg reg_act_regs_data_1_4_sva_8_25_22_enexo_1;
  reg reg_act_regs_data_0_5_sva_8_25_22_enexo;
  reg reg_act_regs_data_1_4_sva_dfm_2_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_130;
  reg reg_is_start_enexo_131;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_131;
  reg reg_act_regs_data_1_4_sva_8_21_0_enexo_1;
  reg reg_act_regs_data_0_5_sva_8_21_0_enexo;
  reg reg_act_regs_data_1_4_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_131;
  reg reg_is_start_enexo_132;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_132;
  reg reg_act_regs_data_1_3_sva_8_30_26_enexo_1;
  reg reg_act_regs_data_0_4_sva_8_30_26_enexo;
  reg reg_act_regs_data_1_3_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_132;
  reg reg_is_start_enexo_133;
  reg reg_act_regs_data_0_4_sva_8_25_22_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_133;
  reg reg_act_regs_data_1_3_sva_8_25_22_enexo_1;
  reg reg_act_regs_data_1_3_sva_dfm_2_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_133;
  reg reg_is_start_enexo_134;
  reg reg_act_regs_data_0_4_sva_8_21_0_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_134;
  reg reg_act_regs_data_1_3_sva_8_21_0_enexo_1;
  reg reg_act_regs_data_1_3_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_134;
  reg reg_is_start_enexo_135;
  reg reg_act_regs_data_0_3_sva_8_30_26_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_135;
  reg reg_act_regs_data_1_2_sva_8_30_26_enexo_1;
  reg reg_act_regs_data_1_2_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_135;
  reg reg_is_start_enexo_136;
  reg reg_act_regs_data_0_3_sva_8_25_22_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_136;
  reg reg_act_regs_data_1_2_sva_8_25_22_enexo_1;
  reg reg_act_regs_data_1_2_sva_dfm_2_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_136;
  reg reg_is_start_enexo_137;
  reg reg_act_regs_data_0_3_sva_8_21_0_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_137;
  reg reg_act_regs_data_1_2_sva_8_21_0_enexo_1;
  reg reg_act_regs_data_1_2_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_137;
  reg reg_is_start_enexo_138;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_138;
  reg reg_act_regs_data_1_1_sva_8_30_26_enexo_1;
  reg reg_act_regs_data_0_10_sva_8_30_26_enexo;
  reg reg_act_regs_data_1_1_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_138;
  reg reg_is_start_enexo_139;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_139;
  reg reg_act_regs_data_1_1_sva_8_25_22_enexo_1;
  reg reg_act_regs_data_0_10_sva_8_25_22_enexo;
  reg reg_act_regs_data_1_1_sva_dfm_2_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_139;
  reg reg_is_start_enexo_140;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_140;
  reg reg_act_regs_data_1_1_sva_8_21_0_enexo_1;
  reg reg_act_regs_data_0_10_sva_8_21_0_enexo;
  reg reg_act_regs_data_1_1_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_140;
  reg reg_is_start_enexo_141;
  reg reg_act_regs_data_0_1_sva_8_30_26_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_141;
  reg reg_act_regs_data_1_0_sva_8_30_26_enexo_1;
  reg reg_act_regs_data_1_0_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_141;
  reg reg_is_start_enexo_142;
  reg reg_act_regs_data_0_1_sva_8_25_22_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_142;
  reg reg_act_regs_data_1_0_sva_8_25_22_enexo_1;
  reg reg_act_regs_data_1_0_sva_dfm_2_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_142;
  reg reg_is_start_enexo_143;
  reg reg_act_regs_data_0_1_sva_8_21_0_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_143;
  reg reg_act_regs_data_1_0_sva_8_21_0_enexo_1;
  reg reg_act_regs_data_1_0_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_143;
  reg reg_is_start_enexo_144;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_144;
  reg reg_act_regs_data_0_15_sva_8_30_26_enexo_1;
  reg reg_ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_1_30_26_enexo;
  reg reg_act_regs_data_0_15_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_144;
  reg reg_is_start_enexo_145;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_145;
  reg reg_ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_1_25_22_enexo;
  reg reg_act_regs_data_0_15_sva_8_25_22_enexo_1;
  reg reg_act_regs_data_0_15_sva_dfm_2_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_145;
  reg reg_is_start_enexo_146;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_146;
  reg reg_act_regs_data_0_15_sva_8_21_0_enexo_1;
  reg reg_act_regs_data_0_15_sva_dfm_2_21_0_enexo;
  reg reg_Silu_for_3_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_146;
  reg reg_is_start_enexo_147;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_147;
  reg reg_act_regs_data_0_14_sva_8_30_26_enexo_1;
  reg reg_ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_1_30_26_enexo;
  reg reg_act_regs_data_0_14_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_147;
  reg reg_is_start_enexo_148;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_148;
  reg reg_ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_1_25_22_enexo;
  reg reg_act_regs_data_0_14_sva_8_25_22_enexo_1;
  reg reg_act_regs_data_0_14_sva_dfm_2_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_148;
  reg reg_is_start_enexo_149;
  reg reg_Silu_for_2_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_149;
  reg reg_act_regs_data_0_14_sva_8_21_0_enexo_1;
  reg reg_act_regs_data_0_14_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_149;
  reg reg_is_start_enexo_150;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_150;
  reg reg_act_regs_data_0_9_sva_8_30_26_enexo_1;
  reg reg_act_regs_data_0_0_sva_8_30_26_enexo;
  reg reg_act_regs_data_0_9_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_150;
  reg reg_is_start_enexo_151;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_151;
  reg reg_act_regs_data_0_9_sva_8_25_22_enexo_1;
  reg reg_act_regs_data_0_0_sva_8_25_22_enexo;
  reg reg_act_regs_data_0_9_sva_dfm_2_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_151;
  reg reg_is_start_enexo_152;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_152;
  reg reg_act_regs_data_0_9_sva_8_21_0_enexo_1;
  reg reg_act_regs_data_0_0_sva_8_21_0_enexo;
  reg reg_act_regs_data_0_9_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_152;
  reg reg_is_start_enexo_153;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_153;
  reg reg_act_regs_data_0_8_sva_8_30_26_enexo_1;
  reg reg_act_regs_data_0_8_sva_dfm_2_30_26_enexo;
  reg reg_ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_1_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_153;
  reg reg_is_start_enexo_154;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_154;
  reg reg_act_regs_data_0_8_sva_8_25_22_enexo_1;
  reg reg_act_regs_data_0_8_sva_dfm_2_25_22_enexo;
  reg reg_ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_1_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_154;
  reg reg_is_start_enexo_155;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_155;
  reg reg_Silu_for_y_8_sva_3_24_0_1_enexo;
  reg reg_act_regs_data_0_8_sva_8_21_0_enexo_1;
  reg reg_act_regs_data_0_8_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_155;
  reg reg_is_start_enexo_156;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_156;
  reg reg_act_regs_data_0_7_sva_8_30_26_enexo_1;
  reg reg_act_regs_data_0_7_sva_dfm_2_30_26_enexo;
  reg reg_ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_1_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_156;
  reg reg_is_start_enexo_157;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_157;
  reg reg_act_regs_data_0_7_sva_8_25_22_enexo_1;
  reg reg_act_regs_data_0_7_sva_dfm_2_25_22_enexo;
  reg reg_ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_1_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_157;
  reg reg_is_start_enexo_158;
  reg reg_Silu_for_y_1_sva_3_24_0_1_enexo;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_158;
  reg reg_act_regs_data_0_7_sva_8_21_0_enexo_1;
  reg reg_act_regs_data_0_7_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_158;
  reg reg_is_start_enexo_159;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_159;
  reg reg_act_regs_data_0_6_sva_8_30_26_enexo_1;
  reg reg_act_regs_data_0_6_sva_dfm_2_30_26_enexo;
  reg reg_ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_1_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_159;
  reg reg_is_start_enexo_160;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_160;
  reg reg_act_regs_data_0_6_sva_8_25_22_enexo_1;
  reg reg_act_regs_data_0_6_sva_dfm_2_25_22_enexo;
  reg reg_ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_1_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_160;
  reg reg_is_start_enexo_161;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_161;
  reg reg_Silu_for_9_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo;
  reg reg_act_regs_data_0_6_sva_8_21_0_enexo_1;
  reg reg_act_regs_data_0_6_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_161;
  reg reg_is_start_enexo_162;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_162;
  reg reg_act_regs_data_0_5_sva_8_30_26_enexo_1;
  reg reg_act_regs_data_0_5_sva_dfm_2_30_26_enexo;
  reg reg_ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_1_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_162;
  reg reg_is_start_enexo_163;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_163;
  reg reg_act_regs_data_0_5_sva_8_25_22_enexo_1;
  reg reg_act_regs_data_0_5_sva_dfm_2_25_22_enexo;
  reg reg_ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_1_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_163;
  reg reg_is_start_enexo_164;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_164;
  reg reg_Silu_for_7_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo;
  reg reg_act_regs_data_0_5_sva_8_21_0_enexo_1;
  reg reg_act_regs_data_0_5_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_164;
  reg reg_is_start_enexo_165;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_165;
  reg reg_act_regs_data_0_4_sva_8_30_26_enexo_1;
  reg reg_act_regs_data_0_4_sva_dfm_2_30_26_enexo;
  reg reg_ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_1_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_165;
  reg reg_is_start_enexo_166;
  reg reg_act_regs_data_0_4_sva_8_25_22_enexo_1;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_166;
  reg reg_ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_1_25_22_enexo;
  reg reg_act_regs_data_0_4_sva_dfm_2_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_166;
  reg reg_is_start_enexo_167;
  reg reg_act_regs_data_0_4_sva_8_21_0_enexo_1;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_167;
  reg reg_act_regs_data_0_4_sva_dfm_2_21_0_enexo;
  reg reg_Silu_for_6_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_167;
  reg reg_is_start_enexo_168;
  reg reg_act_regs_data_0_3_sva_8_30_26_enexo_1;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_168;
  reg reg_act_regs_data_0_3_sva_dfm_2_30_26_enexo;
  reg reg_ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_1_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_168;
  reg reg_is_start_enexo_169;
  reg reg_act_regs_data_0_3_sva_8_25_22_enexo_1;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_169;
  reg reg_ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_1_25_22_enexo;
  reg reg_act_regs_data_0_3_sva_dfm_2_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_169;
  reg reg_is_start_enexo_170;
  reg reg_act_regs_data_0_3_sva_8_21_0_enexo_1;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_170;
  reg reg_act_regs_data_0_3_sva_dfm_2_21_0_enexo;
  reg reg_Silu_for_5_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_170;
  reg reg_is_start_enexo_171;
  reg reg_act_regs_data_0_2_sva_8_30_26_enexo_1;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_171;
  reg reg_ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_1_30_26_enexo;
  reg reg_act_regs_data_0_2_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_171;
  reg reg_is_start_enexo_172;
  reg reg_act_regs_data_0_2_sva_8_25_22_enexo_1;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_172;
  reg reg_ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_1_25_22_enexo;
  reg reg_act_regs_data_0_2_sva_dfm_2_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_172;
  reg reg_is_start_enexo_173;
  reg reg_act_regs_data_0_2_sva_8_21_0_enexo_1;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_173;
  reg reg_act_regs_data_0_2_sva_dfm_2_21_0_enexo;
  reg reg_Silu_for_4_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_173;
  reg reg_act_mem_banks_read_for_mux_15_enexo;
  reg reg_act_mem_banks_read_for_mux_14_enexo;
  reg reg_act_mem_banks_read_for_mux_13_enexo;
  reg reg_act_mem_banks_read_for_mux_12_enexo;
  reg reg_act_mem_banks_read_for_mux_11_enexo;
  reg reg_act_mem_banks_read_for_mux_10_enexo;
  reg reg_act_mem_banks_read_for_mux_9_enexo;
  reg reg_act_mem_banks_read_for_mux_8_enexo;
  reg reg_act_mem_banks_read_for_mux_7_enexo;
  reg reg_act_mem_banks_read_for_mux_6_enexo;
  reg reg_act_mem_banks_read_for_mux_5_enexo;
  reg reg_act_mem_banks_read_for_mux_4_enexo;
  reg reg_act_mem_banks_read_for_mux_3_enexo;
  reg reg_act_mem_banks_read_for_mux_2_enexo;
  reg reg_act_mem_banks_read_for_mux_1_enexo;
  reg reg_act_mem_banks_read_for_mux_enexo;
  reg reg_act_mem_banks_read_for_mux_15_enexo_1;
  reg reg_act_write_req_valid_lpi_1_dfm_5_enexo;
  reg reg_act_mem_banks_read_read_data_lpi_1_dfm_1_31_0_enexo;
  reg reg_act_mem_banks_read_read_data_lpi_1_dfm_1_63_32_enexo;
  reg reg_act_write_req_valid_lpi_1_dfm_5_enexo_1;
  reg reg_act_mem_banks_read_for_mux_14_enexo_1;
  reg reg_act_write_req_valid_lpi_1_dfm_5_enexo_2;
  reg reg_act_mem_banks_read_for_mux_13_enexo_1;
  reg reg_act_mem_banks_read_read_data_lpi_1_dfm_1_95_64_enexo;
  reg reg_act_write_req_valid_lpi_1_dfm_5_enexo_3;
  reg reg_act_mem_banks_read_for_mux_12_enexo_1;
  reg reg_act_mem_banks_read_read_data_lpi_1_dfm_1_127_96_enexo;
  reg reg_act_mem_banks_read_for_mux_11_enexo_1;
  reg reg_act_write_req_valid_lpi_1_dfm_5_enexo_4;
  reg reg_act_mem_banks_read_read_data_lpi_1_dfm_1_159_128_enexo;
  reg reg_act_mem_banks_read_read_data_lpi_1_dfm_1_191_160_enexo;
  reg reg_act_mem_banks_read_for_mux_10_enexo_1;
  reg reg_act_write_req_valid_lpi_1_dfm_5_enexo_5;
  reg reg_act_mem_banks_read_for_mux_9_enexo_1;
  reg reg_act_write_req_valid_lpi_1_dfm_5_enexo_6;
  reg reg_act_mem_banks_read_read_data_lpi_1_dfm_1_223_192_enexo;
  reg reg_act_mem_banks_read_read_data_lpi_1_dfm_1_255_224_enexo;
  reg reg_act_mem_banks_read_for_mux_8_enexo_1;
  reg reg_act_write_req_valid_lpi_1_dfm_5_enexo_7;
  reg reg_act_mem_banks_read_read_data_lpi_1_dfm_1_287_256_enexo;
  reg reg_act_mem_banks_read_for_mux_7_enexo_1;
  reg reg_act_write_req_valid_lpi_1_dfm_5_enexo_8;
  reg reg_act_mem_banks_read_read_data_lpi_1_dfm_1_319_288_enexo;
  reg reg_act_mem_banks_read_for_mux_6_enexo_1;
  reg reg_act_write_req_valid_lpi_1_dfm_5_enexo_9;
  reg reg_act_mem_banks_read_read_data_lpi_1_dfm_1_351_320_enexo;
  reg reg_act_write_req_valid_lpi_1_dfm_5_enexo_10;
  reg reg_act_mem_banks_read_for_mux_5_enexo_1;
  reg reg_act_mem_banks_read_read_data_lpi_1_dfm_1_383_352_enexo;
  reg reg_act_write_req_valid_lpi_1_dfm_5_enexo_11;
  reg reg_act_mem_banks_read_for_mux_4_enexo_1;
  reg reg_act_mem_banks_read_read_data_lpi_1_dfm_1_415_384_enexo;
  reg reg_act_write_req_valid_lpi_1_dfm_5_enexo_12;
  reg reg_act_mem_banks_read_for_mux_3_enexo_1;
  reg reg_act_mem_banks_read_for_mux_2_enexo_1;
  reg reg_act_write_req_valid_lpi_1_dfm_5_enexo_13;
  reg reg_act_mem_banks_read_read_data_lpi_1_dfm_1_447_416_enexo;
  reg reg_act_mem_banks_read_for_mux_1_enexo_1;
  reg reg_act_mem_banks_read_read_data_lpi_1_dfm_1_479_448_enexo;
  reg reg_act_write_req_valid_lpi_1_dfm_5_enexo_14;
  reg reg_act_mem_banks_read_for_mux_enexo_1;
  reg reg_act_mem_banks_read_read_data_lpi_1_dfm_1_511_480_enexo;
  reg reg_act_write_req_valid_lpi_1_dfm_5_enexo_15;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo;
  reg reg_act_config_inst_counter_enexo;
  reg reg_act_regs_data_0_15_1_enexo;
  reg reg_act_regs_data_1_15_1_enexo;
  reg reg_act_regs_data_2_15_1_enexo;
  reg reg_act_regs_data_3_15_1_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_1;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_1;
  reg reg_act_config_inst_counter_enexo_1;
  reg reg_act_regs_data_3_15_2_enexo;
  reg reg_act_regs_data_2_15_2_enexo;
  reg reg_act_regs_data_0_15_2_enexo;
  reg reg_act_regs_data_1_15_2_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_2;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_2;
  reg reg_act_regs_data_2_15_3_enexo;
  reg reg_act_config_inst_counter_enexo_2;
  reg reg_act_regs_data_0_15_3_enexo;
  reg reg_act_regs_data_1_15_3_enexo;
  reg reg_act_regs_data_3_15_3_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_3;
  reg reg_act_regs_data_1_14_1_enexo;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_3;
  reg reg_act_config_inst_counter_enexo_3;
  reg reg_act_regs_data_2_14_1_enexo;
  reg reg_act_regs_data_3_14_1_enexo;
  reg reg_act_regs_data_0_14_1_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_4;
  reg reg_act_regs_data_0_14_2_enexo;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_4;
  reg reg_act_config_inst_counter_enexo_4;
  reg reg_act_regs_data_2_14_2_enexo;
  reg reg_act_regs_data_3_14_2_enexo;
  reg reg_act_regs_data_1_14_2_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_5;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_5;
  reg reg_act_config_inst_counter_enexo_5;
  reg reg_act_regs_data_0_14_3_enexo;
  reg reg_act_regs_data_2_14_3_enexo;
  reg reg_act_regs_data_3_14_3_enexo;
  reg reg_act_regs_data_1_14_3_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_6;
  reg reg_act_regs_data_1_13_1_enexo;
  reg reg_act_regs_data_2_13_1_enexo;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_6;
  reg reg_act_config_inst_counter_enexo_6;
  reg reg_act_regs_data_0_13_1_enexo;
  reg reg_act_regs_data_3_13_1_enexo;
  reg reg_act_regs_data_3_13_2_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_7;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_7;
  reg reg_act_regs_data_0_13_2_enexo;
  reg reg_act_config_inst_counter_enexo_7;
  reg reg_act_regs_data_1_13_2_enexo;
  reg reg_act_regs_data_2_13_2_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_8;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_8;
  reg reg_act_config_inst_counter_enexo_8;
  reg reg_act_regs_data_2_13_3_enexo;
  reg reg_act_regs_data_3_13_3_enexo;
  reg reg_act_regs_data_1_13_3_enexo;
  reg reg_act_regs_data_0_13_3_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_9;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_9;
  reg reg_act_config_inst_counter_enexo_9;
  reg reg_act_regs_data_2_12_1_enexo;
  reg reg_act_regs_data_0_12_1_enexo;
  reg reg_act_regs_data_1_12_1_enexo;
  reg reg_act_regs_data_3_12_1_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_10;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_10;
  reg reg_act_regs_data_2_12_2_enexo;
  reg reg_act_config_inst_counter_enexo_10;
  reg reg_act_regs_data_0_12_2_enexo;
  reg reg_act_regs_data_3_12_2_enexo;
  reg reg_act_regs_data_1_12_2_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_11;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_11;
  reg reg_act_config_inst_counter_enexo_11;
  reg reg_act_regs_data_0_12_3_enexo;
  reg reg_act_regs_data_2_12_3_enexo;
  reg reg_act_regs_data_3_12_3_enexo;
  reg reg_act_regs_data_1_12_3_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_12;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_12;
  reg reg_act_config_inst_counter_enexo_12;
  reg reg_act_regs_data_2_11_1_enexo;
  reg reg_act_regs_data_3_11_1_enexo;
  reg reg_act_regs_data_0_11_1_enexo;
  reg reg_act_regs_data_1_11_1_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_13;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_13;
  reg reg_act_config_inst_counter_enexo_13;
  reg reg_act_regs_data_2_11_2_enexo;
  reg reg_act_regs_data_0_11_2_enexo;
  reg reg_act_regs_data_3_11_2_enexo;
  reg reg_act_regs_data_1_11_2_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_14;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_14;
  reg reg_act_config_inst_counter_enexo_14;
  reg reg_act_regs_data_0_11_3_enexo;
  reg reg_act_regs_data_1_11_3_enexo;
  reg reg_act_regs_data_2_11_3_enexo;
  reg reg_act_regs_data_3_11_3_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_15;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_15;
  reg reg_act_config_inst_counter_enexo_15;
  reg reg_act_regs_data_1_10_1_enexo;
  reg reg_act_regs_data_2_10_1_enexo;
  reg reg_act_regs_data_3_10_1_enexo;
  reg reg_act_regs_data_0_10_1_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_16;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_16;
  reg reg_act_config_inst_counter_enexo_16;
  reg reg_act_regs_data_1_10_2_enexo;
  reg reg_act_regs_data_0_10_2_enexo;
  reg reg_act_regs_data_3_10_2_enexo;
  reg reg_act_regs_data_2_10_2_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_17;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_17;
  reg reg_act_config_inst_counter_enexo_17;
  reg reg_act_regs_data_3_10_3_enexo;
  reg reg_act_regs_data_0_10_3_enexo;
  reg reg_act_regs_data_2_10_3_enexo;
  reg reg_act_regs_data_1_10_3_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_18;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_18;
  reg reg_act_config_inst_counter_enexo_18;
  reg reg_act_regs_data_1_9_1_enexo;
  reg reg_act_regs_data_3_9_1_enexo;
  reg reg_act_regs_data_0_9_1_enexo;
  reg reg_act_regs_data_2_9_1_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_19;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_19;
  reg reg_act_config_inst_counter_enexo_19;
  reg reg_act_regs_data_0_9_2_enexo;
  reg reg_act_regs_data_2_9_2_enexo;
  reg reg_act_regs_data_1_9_2_enexo;
  reg reg_act_regs_data_3_9_2_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_20;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_20;
  reg reg_act_config_inst_counter_enexo_20;
  reg reg_act_regs_data_1_9_3_enexo;
  reg reg_act_regs_data_0_9_3_enexo;
  reg reg_act_regs_data_2_9_3_enexo;
  reg reg_act_regs_data_3_9_3_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_21;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_21;
  reg reg_act_config_inst_counter_enexo_21;
  reg reg_act_regs_data_2_8_1_enexo;
  reg reg_act_regs_data_0_8_1_enexo;
  reg reg_act_regs_data_3_8_1_enexo;
  reg reg_act_regs_data_1_8_1_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_22;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_22;
  reg reg_act_config_inst_counter_enexo_22;
  reg reg_act_regs_data_0_8_2_enexo;
  reg reg_act_regs_data_1_8_2_enexo;
  reg reg_act_regs_data_2_8_2_enexo;
  reg reg_act_regs_data_3_8_2_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_23;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_23;
  reg reg_act_config_inst_counter_enexo_23;
  reg reg_act_regs_data_0_8_3_enexo;
  reg reg_act_regs_data_2_8_3_enexo;
  reg reg_act_regs_data_1_8_3_enexo;
  reg reg_act_regs_data_3_8_3_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_24;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_24;
  reg reg_act_config_inst_counter_enexo_24;
  reg reg_act_regs_data_3_7_1_enexo;
  reg reg_act_regs_data_1_7_1_enexo;
  reg reg_act_regs_data_0_7_1_enexo;
  reg reg_act_regs_data_2_7_1_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_25;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_25;
  reg reg_act_config_inst_counter_enexo_25;
  reg reg_act_regs_data_0_7_2_enexo;
  reg reg_act_regs_data_2_7_2_enexo;
  reg reg_act_regs_data_3_7_2_enexo;
  reg reg_act_regs_data_1_7_2_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_26;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_26;
  reg reg_act_config_inst_counter_enexo_26;
  reg reg_act_regs_data_0_7_3_enexo;
  reg reg_act_regs_data_1_7_3_enexo;
  reg reg_act_regs_data_3_7_3_enexo;
  reg reg_act_regs_data_2_7_3_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_27;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_27;
  reg reg_act_config_inst_counter_enexo_27;
  reg reg_act_regs_data_3_6_1_enexo;
  reg reg_act_regs_data_1_6_1_enexo;
  reg reg_act_regs_data_2_6_1_enexo;
  reg reg_act_regs_data_0_6_1_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_28;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_28;
  reg reg_act_config_inst_counter_enexo_28;
  reg reg_act_regs_data_2_6_2_enexo;
  reg reg_act_regs_data_1_6_2_enexo;
  reg reg_act_regs_data_3_6_2_enexo;
  reg reg_act_regs_data_0_6_2_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_29;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_29;
  reg reg_act_config_inst_counter_enexo_29;
  reg reg_act_regs_data_2_6_3_enexo;
  reg reg_act_regs_data_3_6_3_enexo;
  reg reg_act_regs_data_0_6_3_enexo;
  reg reg_act_regs_data_1_6_3_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_30;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_30;
  reg reg_act_config_inst_counter_enexo_30;
  reg reg_act_regs_data_3_5_1_enexo;
  reg reg_act_regs_data_0_5_1_enexo;
  reg reg_act_regs_data_1_5_1_enexo;
  reg reg_act_regs_data_2_5_1_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_31;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_31;
  reg reg_act_config_inst_counter_enexo_31;
  reg reg_act_regs_data_2_5_2_enexo;
  reg reg_act_regs_data_1_5_2_enexo;
  reg reg_act_regs_data_3_5_2_enexo;
  reg reg_act_regs_data_0_5_2_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_32;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_32;
  reg reg_act_regs_data_0_5_3_enexo;
  reg reg_act_config_inst_counter_enexo_32;
  reg reg_act_regs_data_1_5_3_enexo;
  reg reg_act_regs_data_3_5_3_enexo;
  reg reg_act_regs_data_2_5_3_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_33;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_33;
  reg reg_act_config_inst_counter_enexo_33;
  reg reg_act_regs_data_3_4_1_enexo;
  reg reg_act_regs_data_0_4_1_enexo;
  reg reg_act_regs_data_2_4_1_enexo;
  reg reg_act_regs_data_1_4_1_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_34;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_34;
  reg reg_act_config_inst_counter_enexo_34;
  reg reg_act_regs_data_3_4_2_enexo;
  reg reg_act_regs_data_1_4_2_enexo;
  reg reg_act_regs_data_0_4_2_enexo;
  reg reg_act_regs_data_2_4_2_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_35;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_35;
  reg reg_act_config_inst_counter_enexo_35;
  reg reg_act_regs_data_0_4_3_enexo;
  reg reg_act_regs_data_1_4_3_enexo;
  reg reg_act_regs_data_3_4_3_enexo;
  reg reg_act_regs_data_2_4_3_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_36;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_36;
  reg reg_act_config_inst_counter_enexo_36;
  reg reg_act_regs_data_0_3_1_enexo;
  reg reg_act_regs_data_3_3_1_enexo;
  reg reg_act_regs_data_1_3_1_enexo;
  reg reg_act_regs_data_2_3_1_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_37;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_37;
  reg reg_act_config_inst_counter_enexo_37;
  reg reg_act_regs_data_0_3_2_enexo;
  reg reg_act_regs_data_1_3_2_enexo;
  reg reg_act_regs_data_3_3_2_enexo;
  reg reg_act_regs_data_2_3_2_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_38;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_38;
  reg reg_act_config_inst_counter_enexo_38;
  reg reg_act_regs_data_0_3_3_enexo;
  reg reg_act_regs_data_3_3_3_enexo;
  reg reg_act_regs_data_1_3_3_enexo;
  reg reg_act_regs_data_2_3_3_enexo;
  reg reg_act_regs_data_2_2_1_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_39;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_39;
  reg reg_act_config_inst_counter_enexo_39;
  reg reg_act_regs_data_3_2_1_enexo;
  reg reg_act_regs_data_1_2_1_enexo;
  reg reg_act_regs_data_0_2_1_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_40;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_40;
  reg reg_act_config_inst_counter_enexo_40;
  reg reg_act_regs_data_0_2_2_enexo;
  reg reg_act_regs_data_1_2_2_enexo;
  reg reg_act_regs_data_3_2_2_enexo;
  reg reg_act_regs_data_2_2_2_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_41;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_41;
  reg reg_act_config_inst_counter_enexo_41;
  reg reg_act_regs_data_3_2_3_enexo;
  reg reg_act_regs_data_2_2_3_enexo;
  reg reg_act_regs_data_0_2_3_enexo;
  reg reg_act_regs_data_1_2_3_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_42;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_42;
  reg reg_act_regs_data_2_1_1_enexo;
  reg reg_act_config_inst_counter_enexo_42;
  reg reg_act_regs_data_3_1_1_enexo;
  reg reg_act_regs_data_0_1_1_enexo;
  reg reg_act_regs_data_1_1_1_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_43;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_43;
  reg reg_act_config_inst_counter_enexo_43;
  reg reg_act_regs_data_1_1_2_enexo;
  reg reg_act_regs_data_3_1_2_enexo;
  reg reg_act_regs_data_0_1_2_enexo;
  reg reg_act_regs_data_2_1_2_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_44;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_44;
  reg reg_act_config_inst_counter_enexo_44;
  reg reg_act_regs_data_0_1_3_enexo;
  reg reg_act_regs_data_3_1_3_enexo;
  reg reg_act_regs_data_1_1_3_enexo;
  reg reg_act_regs_data_2_1_3_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_45;
  reg reg_act_regs_data_3_0_1_enexo;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_45;
  reg reg_act_config_inst_counter_enexo_45;
  reg reg_act_regs_data_0_0_1_enexo;
  reg reg_act_regs_data_2_0_1_enexo;
  reg reg_act_regs_data_1_0_1_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_46;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_46;
  reg reg_act_config_inst_counter_enexo_46;
  reg reg_act_regs_data_3_0_2_enexo;
  reg reg_act_regs_data_0_0_2_enexo;
  reg reg_act_regs_data_1_0_2_enexo;
  reg reg_act_regs_data_2_0_2_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_47;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_47;
  reg reg_act_config_inst_counter_enexo_47;
  reg reg_act_regs_data_3_0_3_enexo;
  reg reg_act_regs_data_0_0_3_enexo;
  reg reg_act_regs_data_2_0_3_enexo;
  reg reg_act_regs_data_1_0_3_enexo;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_48;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_48;
  reg reg_act_regs_data_2_15_3_enexo_1;
  reg reg_act_config_inst_counter_enexo_48;
  reg reg_act_regs_data_1_15_enexo;
  reg reg_act_regs_data_0_15_1_enexo_1;
  reg reg_act_regs_data_1_15_1_enexo_1;
  reg reg_act_regs_data_0_15_3_enexo_1;
  reg reg_act_regs_data_1_15_3_enexo_1;
  reg reg_act_regs_data_3_15_2_enexo_1;
  reg reg_act_regs_data_3_15_3_enexo_1;
  reg reg_act_regs_data_2_15_2_enexo_1;
  reg reg_act_regs_data_0_15_2_enexo_1;
  reg reg_act_regs_data_2_15_1_enexo_1;
  reg reg_act_regs_data_3_15_1_enexo_1;
  reg reg_act_regs_data_1_15_2_enexo_1;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_49;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_49;
  reg reg_act_regs_data_2_15_3_enexo_2;
  reg reg_act_config_inst_counter_enexo_49;
  reg reg_act_regs_data_1_15_enexo_1;
  reg reg_act_regs_data_0_15_1_enexo_2;
  reg reg_act_regs_data_1_15_1_enexo_2;
  reg reg_act_regs_data_0_15_3_enexo_2;
  reg reg_act_regs_data_1_15_3_enexo_2;
  reg reg_act_regs_data_3_15_2_enexo_2;
  reg reg_act_regs_data_3_15_3_enexo_2;
  reg reg_act_regs_data_2_15_2_enexo_2;
  reg reg_act_regs_data_0_15_2_enexo_2;
  reg reg_act_regs_data_2_15_1_enexo_2;
  reg reg_act_regs_data_3_15_1_enexo_2;
  reg reg_act_regs_data_1_15_2_enexo_2;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_50;
  reg reg_act_regs_data_0_14_2_enexo_1;
  reg reg_act_regs_data_1_14_1_enexo_1;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_50;
  reg reg_act_config_inst_counter_enexo_50;
  reg reg_act_regs_data_0_14_enexo;
  reg reg_act_regs_data_2_14_2_enexo_1;
  reg reg_act_regs_data_0_14_3_enexo_1;
  reg reg_act_regs_data_3_14_2_enexo_1;
  reg reg_act_regs_data_2_14_1_enexo_1;
  reg reg_act_regs_data_1_14_2_enexo_1;
  reg reg_act_regs_data_3_14_1_enexo_1;
  reg reg_act_regs_data_2_14_3_enexo_1;
  reg reg_act_regs_data_0_14_1_enexo_1;
  reg reg_act_regs_data_3_14_3_enexo_1;
  reg reg_act_regs_data_1_14_3_enexo_1;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_51;
  reg reg_act_regs_data_0_14_2_enexo_2;
  reg reg_act_regs_data_1_14_1_enexo_2;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_51;
  reg reg_act_config_inst_counter_enexo_51;
  reg reg_act_regs_data_0_14_enexo_1;
  reg reg_act_regs_data_2_14_2_enexo_2;
  reg reg_act_regs_data_0_14_3_enexo_2;
  reg reg_act_regs_data_3_14_2_enexo_2;
  reg reg_act_regs_data_2_14_1_enexo_2;
  reg reg_act_regs_data_1_14_2_enexo_2;
  reg reg_act_regs_data_3_14_1_enexo_2;
  reg reg_act_regs_data_2_14_3_enexo_2;
  reg reg_act_regs_data_0_14_1_enexo_2;
  reg reg_act_regs_data_3_14_3_enexo_2;
  reg reg_act_regs_data_1_14_3_enexo_2;
  reg reg_act_regs_data_3_13_2_enexo_1;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_52;
  reg reg_act_regs_data_1_13_1_enexo_1;
  reg reg_act_regs_data_2_13_1_enexo_1;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_52;
  reg reg_act_regs_data_0_13_2_enexo_1;
  reg reg_act_config_inst_counter_enexo_52;
  reg reg_act_regs_data_0_13_1_enexo_1;
  reg reg_act_regs_data_1_13_2_enexo_1;
  reg reg_act_regs_data_3_13_enexo;
  reg reg_act_regs_data_2_13_3_enexo_1;
  reg reg_act_regs_data_2_13_2_enexo_1;
  reg reg_act_regs_data_3_13_3_enexo_1;
  reg reg_act_regs_data_3_13_1_enexo_1;
  reg reg_act_regs_data_1_13_3_enexo_1;
  reg reg_act_regs_data_0_13_3_enexo_1;
  reg reg_act_regs_data_3_13_2_enexo_2;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_53;
  reg reg_act_regs_data_1_13_1_enexo_2;
  reg reg_act_regs_data_2_13_1_enexo_2;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_53;
  reg reg_act_regs_data_0_13_2_enexo_2;
  reg reg_act_config_inst_counter_enexo_53;
  reg reg_act_regs_data_0_13_1_enexo_2;
  reg reg_act_regs_data_1_13_2_enexo_2;
  reg reg_act_regs_data_3_13_enexo_1;
  reg reg_act_regs_data_2_13_3_enexo_2;
  reg reg_act_regs_data_2_13_2_enexo_2;
  reg reg_act_regs_data_3_13_3_enexo_2;
  reg reg_act_regs_data_3_13_1_enexo_2;
  reg reg_act_regs_data_1_13_3_enexo_2;
  reg reg_act_regs_data_0_13_3_enexo_2;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_54;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_54;
  reg reg_act_regs_data_2_12_2_enexo_1;
  reg reg_act_config_inst_counter_enexo_54;
  reg reg_act_regs_data_2_12_1_enexo_1;
  reg reg_act_regs_data_0_12_enexo;
  reg reg_act_regs_data_0_12_1_enexo_1;
  reg reg_act_regs_data_1_12_1_enexo_1;
  reg reg_act_regs_data_0_12_2_enexo_1;
  reg reg_act_regs_data_0_12_3_enexo_1;
  reg reg_act_regs_data_3_12_2_enexo_1;
  reg reg_act_regs_data_2_12_3_enexo_1;
  reg reg_act_regs_data_3_12_3_enexo_1;
  reg reg_act_regs_data_1_12_2_enexo_1;
  reg reg_act_regs_data_1_12_3_enexo_1;
  reg reg_act_regs_data_3_12_1_enexo_1;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_55;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_55;
  reg reg_act_regs_data_2_12_2_enexo_2;
  reg reg_act_config_inst_counter_enexo_55;
  reg reg_act_regs_data_2_12_1_enexo_2;
  reg reg_act_regs_data_0_12_enexo_1;
  reg reg_act_regs_data_0_12_1_enexo_2;
  reg reg_act_regs_data_1_12_1_enexo_2;
  reg reg_act_regs_data_0_12_2_enexo_2;
  reg reg_act_regs_data_0_12_3_enexo_2;
  reg reg_act_regs_data_3_12_2_enexo_2;
  reg reg_act_regs_data_2_12_3_enexo_2;
  reg reg_act_regs_data_3_12_3_enexo_2;
  reg reg_act_regs_data_1_12_2_enexo_2;
  reg reg_act_regs_data_1_12_3_enexo_2;
  reg reg_act_regs_data_3_12_1_enexo_2;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_56;
  reg reg_act_regs_data_2_11_enexo;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_56;
  reg reg_act_config_inst_counter_enexo_56;
  reg reg_act_regs_data_0_11_3_enexo_1;
  reg reg_act_regs_data_2_11_1_enexo_1;
  reg reg_act_regs_data_1_11_3_enexo_1;
  reg reg_act_regs_data_2_11_2_enexo_1;
  reg reg_act_regs_data_0_11_2_enexo_1;
  reg reg_act_regs_data_2_11_3_enexo_1;
  reg reg_act_regs_data_3_11_1_enexo_1;
  reg reg_act_regs_data_0_11_1_enexo_1;
  reg reg_act_regs_data_3_11_3_enexo_1;
  reg reg_act_regs_data_3_11_2_enexo_1;
  reg reg_act_regs_data_1_11_1_enexo_1;
  reg reg_act_regs_data_1_11_2_enexo_1;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_57;
  reg reg_act_regs_data_2_11_enexo_1;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_57;
  reg reg_act_config_inst_counter_enexo_57;
  reg reg_act_regs_data_0_11_3_enexo_2;
  reg reg_act_regs_data_2_11_1_enexo_2;
  reg reg_act_regs_data_1_11_3_enexo_2;
  reg reg_act_regs_data_2_11_2_enexo_2;
  reg reg_act_regs_data_0_11_2_enexo_2;
  reg reg_act_regs_data_2_11_3_enexo_2;
  reg reg_act_regs_data_3_11_1_enexo_2;
  reg reg_act_regs_data_0_11_1_enexo_2;
  reg reg_act_regs_data_3_11_3_enexo_2;
  reg reg_act_regs_data_3_11_2_enexo_2;
  reg reg_act_regs_data_1_11_1_enexo_2;
  reg reg_act_regs_data_1_11_2_enexo_2;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_58;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_58;
  reg reg_act_config_inst_counter_enexo_58;
  reg reg_act_regs_data_1_10_1_enexo_1;
  reg reg_act_regs_data_1_10_2_enexo_1;
  reg reg_act_regs_data_3_10_3_enexo_1;
  reg reg_act_regs_data_2_10_1_enexo_1;
  reg reg_act_regs_data_0_10_enexo;
  reg reg_act_regs_data_0_10_2_enexo_1;
  reg reg_act_regs_data_0_10_3_enexo_1;
  reg reg_act_regs_data_3_10_1_enexo_1;
  reg reg_act_regs_data_2_10_3_enexo_1;
  reg reg_act_regs_data_1_10_3_enexo_1;
  reg reg_act_regs_data_0_10_1_enexo_1;
  reg reg_act_regs_data_3_10_2_enexo_1;
  reg reg_act_regs_data_2_10_2_enexo_1;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_59;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_59;
  reg reg_act_config_inst_counter_enexo_59;
  reg reg_act_regs_data_1_10_1_enexo_2;
  reg reg_act_regs_data_1_10_2_enexo_2;
  reg reg_act_regs_data_3_10_3_enexo_2;
  reg reg_act_regs_data_2_10_1_enexo_2;
  reg reg_act_regs_data_0_10_enexo_1;
  reg reg_act_regs_data_0_10_2_enexo_2;
  reg reg_act_regs_data_0_10_3_enexo_2;
  reg reg_act_regs_data_3_10_1_enexo_2;
  reg reg_act_regs_data_2_10_3_enexo_2;
  reg reg_act_regs_data_1_10_3_enexo_2;
  reg reg_act_regs_data_0_10_1_enexo_2;
  reg reg_act_regs_data_3_10_2_enexo_2;
  reg reg_act_regs_data_2_10_2_enexo_2;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_60;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_60;
  reg reg_act_config_inst_counter_enexo_60;
  reg reg_act_regs_data_1_9_3_enexo_1;
  reg reg_act_regs_data_0_9_2_enexo_1;
  reg reg_act_regs_data_1_9_1_enexo_1;
  reg reg_act_regs_data_1_9_enexo;
  reg reg_act_regs_data_0_9_3_enexo_1;
  reg reg_act_regs_data_2_9_3_enexo_1;
  reg reg_act_regs_data_2_9_2_enexo_1;
  reg reg_act_regs_data_3_9_1_enexo_1;
  reg reg_act_regs_data_1_9_2_enexo_1;
  reg reg_act_regs_data_3_9_2_enexo_1;
  reg reg_act_regs_data_0_9_1_enexo_1;
  reg reg_act_regs_data_3_9_3_enexo_1;
  reg reg_act_regs_data_2_9_1_enexo_1;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_61;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_61;
  reg reg_act_config_inst_counter_enexo_61;
  reg reg_act_regs_data_1_9_3_enexo_2;
  reg reg_act_regs_data_0_9_2_enexo_2;
  reg reg_act_regs_data_1_9_1_enexo_2;
  reg reg_act_regs_data_1_9_enexo_1;
  reg reg_act_regs_data_0_9_3_enexo_2;
  reg reg_act_regs_data_2_9_3_enexo_2;
  reg reg_act_regs_data_2_9_2_enexo_2;
  reg reg_act_regs_data_3_9_1_enexo_2;
  reg reg_act_regs_data_1_9_2_enexo_2;
  reg reg_act_regs_data_3_9_2_enexo_2;
  reg reg_act_regs_data_0_9_1_enexo_2;
  reg reg_act_regs_data_3_9_3_enexo_2;
  reg reg_act_regs_data_2_9_1_enexo_2;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_62;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_62;
  reg reg_act_config_inst_counter_enexo_62;
  reg reg_act_regs_data_2_8_enexo;
  reg reg_act_regs_data_0_8_2_enexo_1;
  reg reg_act_regs_data_1_8_2_enexo_1;
  reg reg_act_regs_data_2_8_1_enexo_1;
  reg reg_act_regs_data_0_8_1_enexo_1;
  reg reg_act_regs_data_0_8_3_enexo_1;
  reg reg_act_regs_data_2_8_2_enexo_1;
  reg reg_act_regs_data_3_8_1_enexo_1;
  reg reg_act_regs_data_2_8_3_enexo_1;
  reg reg_act_regs_data_3_8_2_enexo_1;
  reg reg_act_regs_data_1_8_1_enexo_1;
  reg reg_act_regs_data_1_8_3_enexo_1;
  reg reg_act_regs_data_3_8_3_enexo_1;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_63;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_63;
  reg reg_act_config_inst_counter_enexo_63;
  reg reg_act_regs_data_2_8_enexo_1;
  reg reg_act_regs_data_0_8_2_enexo_2;
  reg reg_act_regs_data_1_8_2_enexo_2;
  reg reg_act_regs_data_2_8_1_enexo_2;
  reg reg_act_regs_data_0_8_1_enexo_2;
  reg reg_act_regs_data_0_8_3_enexo_2;
  reg reg_act_regs_data_2_8_2_enexo_2;
  reg reg_act_regs_data_3_8_1_enexo_2;
  reg reg_act_regs_data_2_8_3_enexo_2;
  reg reg_act_regs_data_3_8_2_enexo_2;
  reg reg_act_regs_data_1_8_1_enexo_2;
  reg reg_act_regs_data_1_8_3_enexo_2;
  reg reg_act_regs_data_3_8_3_enexo_2;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_64;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_64;
  reg reg_act_config_inst_counter_enexo_64;
  reg reg_act_regs_data_0_7_3_enexo_1;
  reg reg_act_regs_data_1_7_3_enexo_1;
  reg reg_act_regs_data_3_7_3_enexo_1;
  reg reg_act_regs_data_1_7_enexo;
  reg reg_act_regs_data_0_7_2_enexo_1;
  reg reg_act_regs_data_2_7_2_enexo_1;
  reg reg_act_regs_data_2_7_3_enexo_1;
  reg reg_act_regs_data_3_7_2_enexo_1;
  reg reg_act_regs_data_3_7_1_enexo_1;
  reg reg_act_regs_data_1_7_1_enexo_1;
  reg reg_act_regs_data_1_7_2_enexo_1;
  reg reg_act_regs_data_0_7_1_enexo_1;
  reg reg_act_regs_data_2_7_1_enexo_1;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_65;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_65;
  reg reg_act_config_inst_counter_enexo_65;
  reg reg_act_regs_data_0_7_3_enexo_2;
  reg reg_act_regs_data_1_7_3_enexo_2;
  reg reg_act_regs_data_3_7_3_enexo_2;
  reg reg_act_regs_data_1_7_enexo_1;
  reg reg_act_regs_data_0_7_2_enexo_2;
  reg reg_act_regs_data_2_7_2_enexo_2;
  reg reg_act_regs_data_2_7_3_enexo_2;
  reg reg_act_regs_data_3_7_2_enexo_2;
  reg reg_act_regs_data_3_7_1_enexo_2;
  reg reg_act_regs_data_1_7_1_enexo_2;
  reg reg_act_regs_data_1_7_2_enexo_2;
  reg reg_act_regs_data_0_7_1_enexo_2;
  reg reg_act_regs_data_2_7_1_enexo_2;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_66;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_66;
  reg reg_act_config_inst_counter_enexo_66;
  reg reg_act_regs_data_3_6_1_enexo_1;
  reg reg_act_regs_data_1_6_1_enexo_1;
  reg reg_act_regs_data_2_6_3_enexo_1;
  reg reg_act_regs_data_3_6_3_enexo_1;
  reg reg_act_regs_data_3_6_enexo;
  reg reg_act_regs_data_2_6_1_enexo_1;
  reg reg_act_regs_data_2_6_2_enexo_1;
  reg reg_act_regs_data_0_6_3_enexo_1;
  reg reg_act_regs_data_1_6_3_enexo_1;
  reg reg_act_regs_data_1_6_2_enexo_1;
  reg reg_act_regs_data_0_6_1_enexo_1;
  reg reg_act_regs_data_3_6_2_enexo_1;
  reg reg_act_regs_data_0_6_2_enexo_1;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_67;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_67;
  reg reg_act_config_inst_counter_enexo_67;
  reg reg_act_regs_data_3_6_1_enexo_2;
  reg reg_act_regs_data_1_6_1_enexo_2;
  reg reg_act_regs_data_2_6_3_enexo_2;
  reg reg_act_regs_data_3_6_3_enexo_2;
  reg reg_act_regs_data_3_6_enexo_1;
  reg reg_act_regs_data_2_6_1_enexo_2;
  reg reg_act_regs_data_2_6_2_enexo_2;
  reg reg_act_regs_data_0_6_3_enexo_2;
  reg reg_act_regs_data_1_6_3_enexo_2;
  reg reg_act_regs_data_1_6_2_enexo_2;
  reg reg_act_regs_data_0_6_1_enexo_2;
  reg reg_act_regs_data_3_6_2_enexo_2;
  reg reg_act_regs_data_0_6_2_enexo_2;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_68;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_68;
  reg reg_act_regs_data_0_5_3_enexo_1;
  reg reg_act_config_inst_counter_enexo_68;
  reg reg_act_regs_data_2_5_2_enexo_1;
  reg reg_act_regs_data_3_5_1_enexo_1;
  reg reg_act_regs_data_0_5_1_enexo_1;
  reg reg_act_regs_data_1_5_enexo;
  reg reg_act_regs_data_1_5_1_enexo_1;
  reg reg_act_regs_data_1_5_2_enexo_1;
  reg reg_act_regs_data_3_5_2_enexo_1;
  reg reg_act_regs_data_0_5_2_enexo_1;
  reg reg_act_regs_data_1_5_3_enexo_1;
  reg reg_act_regs_data_3_5_3_enexo_1;
  reg reg_act_regs_data_2_5_1_enexo_1;
  reg reg_act_regs_data_2_5_3_enexo_1;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_69;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_69;
  reg reg_act_regs_data_0_5_3_enexo_2;
  reg reg_act_config_inst_counter_enexo_69;
  reg reg_act_regs_data_2_5_2_enexo_2;
  reg reg_act_regs_data_3_5_1_enexo_2;
  reg reg_act_regs_data_0_5_1_enexo_2;
  reg reg_act_regs_data_1_5_enexo_1;
  reg reg_act_regs_data_1_5_1_enexo_2;
  reg reg_act_regs_data_1_5_2_enexo_2;
  reg reg_act_regs_data_3_5_2_enexo_2;
  reg reg_act_regs_data_0_5_2_enexo_2;
  reg reg_act_regs_data_1_5_3_enexo_2;
  reg reg_act_regs_data_3_5_3_enexo_2;
  reg reg_act_regs_data_2_5_1_enexo_2;
  reg reg_act_regs_data_2_5_3_enexo_2;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_70;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_70;
  reg reg_act_config_inst_counter_enexo_70;
  reg reg_act_regs_data_0_4_3_enexo_1;
  reg reg_act_regs_data_3_4_1_enexo_1;
  reg reg_act_regs_data_3_4_2_enexo_1;
  reg reg_act_regs_data_1_4_3_enexo_1;
  reg reg_act_regs_data_0_4_1_enexo_1;
  reg reg_act_regs_data_2_4_1_enexo_1;
  reg reg_act_regs_data_3_4_3_enexo_1;
  reg reg_act_regs_data_1_4_2_enexo_1;
  reg reg_act_regs_data_3_4_enexo;
  reg reg_act_regs_data_2_4_3_enexo_1;
  reg reg_act_regs_data_1_4_1_enexo_1;
  reg reg_act_regs_data_0_4_2_enexo_1;
  reg reg_act_regs_data_2_4_2_enexo_1;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_71;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_71;
  reg reg_act_config_inst_counter_enexo_71;
  reg reg_act_regs_data_0_4_3_enexo_2;
  reg reg_act_regs_data_3_4_1_enexo_2;
  reg reg_act_regs_data_3_4_2_enexo_2;
  reg reg_act_regs_data_1_4_3_enexo_2;
  reg reg_act_regs_data_0_4_1_enexo_2;
  reg reg_act_regs_data_2_4_1_enexo_2;
  reg reg_act_regs_data_3_4_3_enexo_2;
  reg reg_act_regs_data_1_4_2_enexo_2;
  reg reg_act_regs_data_3_4_enexo_1;
  reg reg_act_regs_data_2_4_3_enexo_2;
  reg reg_act_regs_data_1_4_1_enexo_2;
  reg reg_act_regs_data_0_4_2_enexo_2;
  reg reg_act_regs_data_2_4_2_enexo_2;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_72;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_72;
  reg reg_act_config_inst_counter_enexo_72;
  reg reg_act_regs_data_0_3_3_enexo_1;
  reg reg_act_regs_data_3_3_3_enexo_1;
  reg reg_act_regs_data_0_3_1_enexo_1;
  reg reg_act_regs_data_3_3_enexo;
  reg reg_act_regs_data_3_3_1_enexo_1;
  reg reg_act_regs_data_1_3_1_enexo_1;
  reg reg_act_regs_data_0_3_2_enexo_1;
  reg reg_act_regs_data_1_3_3_enexo_1;
  reg reg_act_regs_data_1_3_2_enexo_1;
  reg reg_act_regs_data_3_3_2_enexo_1;
  reg reg_act_regs_data_2_3_1_enexo_1;
  reg reg_act_regs_data_2_3_3_enexo_1;
  reg reg_act_regs_data_2_3_2_enexo_1;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_73;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_73;
  reg reg_act_config_inst_counter_enexo_73;
  reg reg_act_regs_data_0_3_3_enexo_2;
  reg reg_act_regs_data_3_3_3_enexo_2;
  reg reg_act_regs_data_0_3_1_enexo_2;
  reg reg_act_regs_data_3_3_enexo_1;
  reg reg_act_regs_data_3_3_1_enexo_2;
  reg reg_act_regs_data_1_3_1_enexo_2;
  reg reg_act_regs_data_0_3_2_enexo_2;
  reg reg_act_regs_data_1_3_3_enexo_2;
  reg reg_act_regs_data_1_3_2_enexo_2;
  reg reg_act_regs_data_3_3_2_enexo_2;
  reg reg_act_regs_data_2_3_1_enexo_2;
  reg reg_act_regs_data_2_3_3_enexo_2;
  reg reg_act_regs_data_2_3_2_enexo_2;
  reg reg_act_regs_data_2_2_1_enexo_1;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_74;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_74;
  reg reg_act_config_inst_counter_enexo_74;
  reg reg_act_regs_data_3_2_enexo;
  reg reg_act_regs_data_0_2_2_enexo_1;
  reg reg_act_regs_data_3_2_1_enexo_1;
  reg reg_act_regs_data_3_2_3_enexo_1;
  reg reg_act_regs_data_2_2_3_enexo_1;
  reg reg_act_regs_data_1_2_1_enexo_1;
  reg reg_act_regs_data_1_2_2_enexo_1;
  reg reg_act_regs_data_3_2_2_enexo_1;
  reg reg_act_regs_data_2_2_2_enexo_1;
  reg reg_act_regs_data_0_2_3_enexo_1;
  reg reg_act_regs_data_0_2_1_enexo_1;
  reg reg_act_regs_data_1_2_3_enexo_1;
  reg reg_act_regs_data_2_2_1_enexo_2;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_75;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_75;
  reg reg_act_config_inst_counter_enexo_75;
  reg reg_act_regs_data_3_2_enexo_1;
  reg reg_act_regs_data_0_2_2_enexo_2;
  reg reg_act_regs_data_3_2_1_enexo_2;
  reg reg_act_regs_data_3_2_3_enexo_2;
  reg reg_act_regs_data_2_2_3_enexo_2;
  reg reg_act_regs_data_1_2_1_enexo_2;
  reg reg_act_regs_data_1_2_2_enexo_2;
  reg reg_act_regs_data_3_2_2_enexo_2;
  reg reg_act_regs_data_2_2_2_enexo_2;
  reg reg_act_regs_data_0_2_3_enexo_2;
  reg reg_act_regs_data_0_2_1_enexo_2;
  reg reg_act_regs_data_1_2_3_enexo_2;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_76;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_76;
  reg reg_act_regs_data_2_1_1_enexo_1;
  reg reg_act_config_inst_counter_enexo_76;
  reg reg_act_regs_data_1_1_2_enexo_1;
  reg reg_act_regs_data_0_1_3_enexo_1;
  reg reg_act_regs_data_3_1_1_enexo_1;
  reg reg_act_regs_data_2_1_enexo;
  reg reg_act_regs_data_0_1_1_enexo_1;
  reg reg_act_regs_data_3_1_2_enexo_1;
  reg reg_act_regs_data_1_1_1_enexo_1;
  reg reg_act_regs_data_0_1_2_enexo_1;
  reg reg_act_regs_data_2_1_2_enexo_1;
  reg reg_act_regs_data_3_1_3_enexo_1;
  reg reg_act_regs_data_1_1_3_enexo_1;
  reg reg_act_regs_data_2_1_3_enexo_1;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_77;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_77;
  reg reg_act_regs_data_2_1_1_enexo_2;
  reg reg_act_config_inst_counter_enexo_77;
  reg reg_act_regs_data_1_1_2_enexo_2;
  reg reg_act_regs_data_0_1_3_enexo_2;
  reg reg_act_regs_data_3_1_1_enexo_2;
  reg reg_act_regs_data_2_1_enexo_1;
  reg reg_act_regs_data_0_1_1_enexo_2;
  reg reg_act_regs_data_3_1_2_enexo_2;
  reg reg_act_regs_data_1_1_1_enexo_2;
  reg reg_act_regs_data_0_1_2_enexo_2;
  reg reg_act_regs_data_2_1_2_enexo_2;
  reg reg_act_regs_data_3_1_3_enexo_2;
  reg reg_act_regs_data_1_1_3_enexo_2;
  reg reg_act_regs_data_2_1_3_enexo_2;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_78;
  reg reg_act_regs_data_3_0_1_enexo_1;
  reg reg_act_regs_data_3_0_enexo;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_78;
  reg reg_act_config_inst_counter_enexo_78;
  reg reg_act_regs_data_3_0_3_enexo_1;
  reg reg_act_regs_data_0_0_3_enexo_1;
  reg reg_act_regs_data_0_0_1_enexo_1;
  reg reg_act_regs_data_3_0_2_enexo_1;
  reg reg_act_regs_data_2_0_1_enexo_1;
  reg reg_act_regs_data_0_0_2_enexo_1;
  reg reg_act_regs_data_1_0_2_enexo_1;
  reg reg_act_regs_data_2_0_3_enexo_1;
  reg reg_act_regs_data_1_0_1_enexo_1;
  reg reg_act_regs_data_2_0_2_enexo_1;
  reg reg_act_regs_data_1_0_3_enexo_1;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_79;
  reg reg_act_regs_data_3_0_1_enexo_2;
  reg reg_act_regs_data_3_0_enexo_1;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_79;
  reg reg_act_config_inst_counter_enexo_79;
  reg reg_act_regs_data_3_0_3_enexo_2;
  reg reg_act_regs_data_0_0_3_enexo_2;
  reg reg_act_regs_data_0_0_1_enexo_2;
  reg reg_act_regs_data_3_0_2_enexo_2;
  reg reg_act_regs_data_2_0_1_enexo_2;
  reg reg_act_regs_data_0_0_2_enexo_2;
  reg reg_act_regs_data_1_0_2_enexo_2;
  reg reg_act_regs_data_2_0_3_enexo_2;
  reg reg_act_regs_data_1_0_1_enexo_2;
  reg reg_act_regs_data_2_0_2_enexo_2;
  reg reg_act_regs_data_1_0_3_enexo_2;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_80;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_80;
  reg reg_act_config_inst_counter_enexo_80;
  reg reg_act_regs_data_1_15_enexo_2;
  reg reg_act_regs_data_0_15_1_enexo_3;
  reg reg_act_regs_data_1_15_1_enexo_3;
  reg reg_act_regs_data_2_15_1_enexo_3;
  reg reg_act_regs_data_3_15_1_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_81;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_81;
  reg reg_act_config_inst_counter_enexo_81;
  reg reg_act_regs_data_1_15_enexo_3;
  reg reg_act_regs_data_3_15_2_enexo_3;
  reg reg_act_regs_data_2_15_2_enexo_3;
  reg reg_act_regs_data_0_15_2_enexo_3;
  reg reg_act_regs_data_1_15_2_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_82;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_82;
  reg reg_act_regs_data_2_15_3_enexo_3;
  reg reg_act_config_inst_counter_enexo_82;
  reg reg_act_regs_data_1_15_enexo_4;
  reg reg_act_regs_data_0_15_3_enexo_3;
  reg reg_act_regs_data_1_15_3_enexo_3;
  reg reg_act_regs_data_3_15_3_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_83;
  reg reg_act_regs_data_1_14_1_enexo_3;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_83;
  reg reg_act_config_inst_counter_enexo_83;
  reg reg_act_regs_data_0_14_enexo_2;
  reg reg_act_regs_data_2_14_1_enexo_3;
  reg reg_act_regs_data_3_14_1_enexo_3;
  reg reg_act_regs_data_0_14_1_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_84;
  reg reg_act_regs_data_0_14_2_enexo_3;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_84;
  reg reg_act_config_inst_counter_enexo_84;
  reg reg_act_regs_data_0_14_enexo_3;
  reg reg_act_regs_data_2_14_2_enexo_3;
  reg reg_act_regs_data_3_14_2_enexo_3;
  reg reg_act_regs_data_1_14_2_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_85;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_85;
  reg reg_act_config_inst_counter_enexo_85;
  reg reg_act_regs_data_0_14_enexo_4;
  reg reg_act_regs_data_0_14_3_enexo_3;
  reg reg_act_regs_data_2_14_3_enexo_3;
  reg reg_act_regs_data_3_14_3_enexo_3;
  reg reg_act_regs_data_1_14_3_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_86;
  reg reg_act_regs_data_1_13_1_enexo_3;
  reg reg_act_regs_data_2_13_1_enexo_3;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_86;
  reg reg_act_config_inst_counter_enexo_86;
  reg reg_act_regs_data_0_13_1_enexo_3;
  reg reg_act_regs_data_3_13_enexo_2;
  reg reg_act_regs_data_3_13_1_enexo_3;
  reg reg_act_regs_data_3_13_2_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_87;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_87;
  reg reg_act_regs_data_0_13_2_enexo_3;
  reg reg_act_config_inst_counter_enexo_87;
  reg reg_act_regs_data_1_13_2_enexo_3;
  reg reg_act_regs_data_3_13_enexo_3;
  reg reg_act_regs_data_2_13_2_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_88;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_88;
  reg reg_act_config_inst_counter_enexo_88;
  reg reg_act_regs_data_3_13_enexo_4;
  reg reg_act_regs_data_2_13_3_enexo_3;
  reg reg_act_regs_data_3_13_3_enexo_3;
  reg reg_act_regs_data_1_13_3_enexo_3;
  reg reg_act_regs_data_0_13_3_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_89;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_89;
  reg reg_act_config_inst_counter_enexo_89;
  reg reg_act_regs_data_2_12_1_enexo_3;
  reg reg_act_regs_data_0_12_enexo_2;
  reg reg_act_regs_data_0_12_1_enexo_3;
  reg reg_act_regs_data_1_12_1_enexo_3;
  reg reg_act_regs_data_3_12_1_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_90;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_90;
  reg reg_act_regs_data_2_12_2_enexo_3;
  reg reg_act_config_inst_counter_enexo_90;
  reg reg_act_regs_data_0_12_enexo_3;
  reg reg_act_regs_data_0_12_2_enexo_3;
  reg reg_act_regs_data_3_12_2_enexo_3;
  reg reg_act_regs_data_1_12_2_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_91;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_91;
  reg reg_act_config_inst_counter_enexo_91;
  reg reg_act_regs_data_0_12_enexo_4;
  reg reg_act_regs_data_0_12_3_enexo_3;
  reg reg_act_regs_data_2_12_3_enexo_3;
  reg reg_act_regs_data_3_12_3_enexo_3;
  reg reg_act_regs_data_1_12_3_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_92;
  reg reg_act_regs_data_2_11_enexo_2;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_92;
  reg reg_act_config_inst_counter_enexo_92;
  reg reg_act_regs_data_2_11_1_enexo_3;
  reg reg_act_regs_data_3_11_1_enexo_3;
  reg reg_act_regs_data_0_11_1_enexo_3;
  reg reg_act_regs_data_1_11_1_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_93;
  reg reg_act_regs_data_2_11_enexo_3;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_93;
  reg reg_act_config_inst_counter_enexo_93;
  reg reg_act_regs_data_2_11_2_enexo_3;
  reg reg_act_regs_data_0_11_2_enexo_3;
  reg reg_act_regs_data_3_11_2_enexo_3;
  reg reg_act_regs_data_1_11_2_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_94;
  reg reg_act_regs_data_2_11_enexo_4;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_94;
  reg reg_act_config_inst_counter_enexo_94;
  reg reg_act_regs_data_0_11_3_enexo_3;
  reg reg_act_regs_data_1_11_3_enexo_3;
  reg reg_act_regs_data_2_11_3_enexo_3;
  reg reg_act_regs_data_3_11_3_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_95;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_95;
  reg reg_act_config_inst_counter_enexo_95;
  reg reg_act_regs_data_1_10_1_enexo_3;
  reg reg_act_regs_data_2_10_1_enexo_3;
  reg reg_act_regs_data_0_10_enexo_2;
  reg reg_act_regs_data_3_10_1_enexo_3;
  reg reg_act_regs_data_0_10_1_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_96;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_96;
  reg reg_act_config_inst_counter_enexo_96;
  reg reg_act_regs_data_1_10_2_enexo_3;
  reg reg_act_regs_data_0_10_enexo_3;
  reg reg_act_regs_data_0_10_2_enexo_3;
  reg reg_act_regs_data_3_10_2_enexo_3;
  reg reg_act_regs_data_2_10_2_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_97;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_97;
  reg reg_act_config_inst_counter_enexo_97;
  reg reg_act_regs_data_3_10_3_enexo_3;
  reg reg_act_regs_data_0_10_enexo_4;
  reg reg_act_regs_data_0_10_3_enexo_3;
  reg reg_act_regs_data_2_10_3_enexo_3;
  reg reg_act_regs_data_1_10_3_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_98;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_98;
  reg reg_act_config_inst_counter_enexo_98;
  reg reg_act_regs_data_1_9_1_enexo_3;
  reg reg_act_regs_data_1_9_enexo_2;
  reg reg_act_regs_data_3_9_1_enexo_3;
  reg reg_act_regs_data_0_9_1_enexo_3;
  reg reg_act_regs_data_2_9_1_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_99;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_99;
  reg reg_act_config_inst_counter_enexo_99;
  reg reg_act_regs_data_0_9_2_enexo_3;
  reg reg_act_regs_data_1_9_enexo_3;
  reg reg_act_regs_data_2_9_2_enexo_3;
  reg reg_act_regs_data_1_9_2_enexo_3;
  reg reg_act_regs_data_3_9_2_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_100;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_100;
  reg reg_act_config_inst_counter_enexo_100;
  reg reg_act_regs_data_1_9_3_enexo_3;
  reg reg_act_regs_data_1_9_enexo_4;
  reg reg_act_regs_data_0_9_3_enexo_3;
  reg reg_act_regs_data_2_9_3_enexo_3;
  reg reg_act_regs_data_3_9_3_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_101;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_101;
  reg reg_act_config_inst_counter_enexo_101;
  reg reg_act_regs_data_2_8_enexo_2;
  reg reg_act_regs_data_2_8_1_enexo_3;
  reg reg_act_regs_data_0_8_1_enexo_3;
  reg reg_act_regs_data_3_8_1_enexo_3;
  reg reg_act_regs_data_1_8_1_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_102;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_102;
  reg reg_act_config_inst_counter_enexo_102;
  reg reg_act_regs_data_2_8_enexo_3;
  reg reg_act_regs_data_0_8_2_enexo_3;
  reg reg_act_regs_data_1_8_2_enexo_3;
  reg reg_act_regs_data_2_8_2_enexo_3;
  reg reg_act_regs_data_3_8_2_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_103;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_103;
  reg reg_act_config_inst_counter_enexo_103;
  reg reg_act_regs_data_2_8_enexo_4;
  reg reg_act_regs_data_0_8_3_enexo_3;
  reg reg_act_regs_data_2_8_3_enexo_3;
  reg reg_act_regs_data_1_8_3_enexo_3;
  reg reg_act_regs_data_3_8_3_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_104;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_104;
  reg reg_act_config_inst_counter_enexo_104;
  reg reg_act_regs_data_1_7_enexo_2;
  reg reg_act_regs_data_3_7_1_enexo_3;
  reg reg_act_regs_data_1_7_1_enexo_3;
  reg reg_act_regs_data_0_7_1_enexo_3;
  reg reg_act_regs_data_2_7_1_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_105;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_105;
  reg reg_act_config_inst_counter_enexo_105;
  reg reg_act_regs_data_1_7_enexo_3;
  reg reg_act_regs_data_0_7_2_enexo_3;
  reg reg_act_regs_data_2_7_2_enexo_3;
  reg reg_act_regs_data_3_7_2_enexo_3;
  reg reg_act_regs_data_1_7_2_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_106;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_106;
  reg reg_act_config_inst_counter_enexo_106;
  reg reg_act_regs_data_0_7_3_enexo_3;
  reg reg_act_regs_data_1_7_3_enexo_3;
  reg reg_act_regs_data_3_7_3_enexo_3;
  reg reg_act_regs_data_1_7_enexo_4;
  reg reg_act_regs_data_2_7_3_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_107;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_107;
  reg reg_act_config_inst_counter_enexo_107;
  reg reg_act_regs_data_3_6_1_enexo_3;
  reg reg_act_regs_data_1_6_1_enexo_3;
  reg reg_act_regs_data_3_6_enexo_2;
  reg reg_act_regs_data_2_6_1_enexo_3;
  reg reg_act_regs_data_0_6_1_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_108;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_108;
  reg reg_act_config_inst_counter_enexo_108;
  reg reg_act_regs_data_3_6_enexo_3;
  reg reg_act_regs_data_2_6_2_enexo_3;
  reg reg_act_regs_data_1_6_2_enexo_3;
  reg reg_act_regs_data_3_6_2_enexo_3;
  reg reg_act_regs_data_0_6_2_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_109;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_109;
  reg reg_act_config_inst_counter_enexo_109;
  reg reg_act_regs_data_2_6_3_enexo_3;
  reg reg_act_regs_data_3_6_3_enexo_3;
  reg reg_act_regs_data_3_6_enexo_4;
  reg reg_act_regs_data_0_6_3_enexo_3;
  reg reg_act_regs_data_1_6_3_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_110;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_110;
  reg reg_act_config_inst_counter_enexo_110;
  reg reg_act_regs_data_3_5_1_enexo_3;
  reg reg_act_regs_data_0_5_1_enexo_3;
  reg reg_act_regs_data_1_5_enexo_2;
  reg reg_act_regs_data_1_5_1_enexo_3;
  reg reg_act_regs_data_2_5_1_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_111;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_111;
  reg reg_act_config_inst_counter_enexo_111;
  reg reg_act_regs_data_2_5_2_enexo_3;
  reg reg_act_regs_data_1_5_enexo_3;
  reg reg_act_regs_data_1_5_2_enexo_3;
  reg reg_act_regs_data_3_5_2_enexo_3;
  reg reg_act_regs_data_0_5_2_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_112;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_112;
  reg reg_act_regs_data_0_5_3_enexo_3;
  reg reg_act_config_inst_counter_enexo_112;
  reg reg_act_regs_data_1_5_enexo_4;
  reg reg_act_regs_data_1_5_3_enexo_3;
  reg reg_act_regs_data_3_5_3_enexo_3;
  reg reg_act_regs_data_2_5_3_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_113;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_113;
  reg reg_act_config_inst_counter_enexo_113;
  reg reg_act_regs_data_3_4_1_enexo_3;
  reg reg_act_regs_data_0_4_1_enexo_3;
  reg reg_act_regs_data_2_4_1_enexo_3;
  reg reg_act_regs_data_3_4_enexo_2;
  reg reg_act_regs_data_1_4_1_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_114;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_114;
  reg reg_act_config_inst_counter_enexo_114;
  reg reg_act_regs_data_3_4_2_enexo_3;
  reg reg_act_regs_data_1_4_2_enexo_3;
  reg reg_act_regs_data_3_4_enexo_3;
  reg reg_act_regs_data_0_4_2_enexo_3;
  reg reg_act_regs_data_2_4_2_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_115;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_115;
  reg reg_act_config_inst_counter_enexo_115;
  reg reg_act_regs_data_0_4_3_enexo_3;
  reg reg_act_regs_data_1_4_3_enexo_3;
  reg reg_act_regs_data_3_4_3_enexo_3;
  reg reg_act_regs_data_3_4_enexo_4;
  reg reg_act_regs_data_2_4_3_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_116;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_116;
  reg reg_act_config_inst_counter_enexo_116;
  reg reg_act_regs_data_0_3_1_enexo_3;
  reg reg_act_regs_data_3_3_enexo_2;
  reg reg_act_regs_data_3_3_1_enexo_3;
  reg reg_act_regs_data_1_3_1_enexo_3;
  reg reg_act_regs_data_2_3_1_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_117;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_117;
  reg reg_act_config_inst_counter_enexo_117;
  reg reg_act_regs_data_3_3_enexo_3;
  reg reg_act_regs_data_0_3_2_enexo_3;
  reg reg_act_regs_data_1_3_2_enexo_3;
  reg reg_act_regs_data_3_3_2_enexo_3;
  reg reg_act_regs_data_2_3_2_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_118;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_118;
  reg reg_act_config_inst_counter_enexo_118;
  reg reg_act_regs_data_0_3_3_enexo_3;
  reg reg_act_regs_data_3_3_3_enexo_3;
  reg reg_act_regs_data_3_3_enexo_4;
  reg reg_act_regs_data_1_3_3_enexo_3;
  reg reg_act_regs_data_2_3_3_enexo_3;
  reg reg_act_regs_data_2_2_1_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_119;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_119;
  reg reg_act_config_inst_counter_enexo_119;
  reg reg_act_regs_data_3_2_enexo_2;
  reg reg_act_regs_data_3_2_1_enexo_3;
  reg reg_act_regs_data_1_2_1_enexo_3;
  reg reg_act_regs_data_0_2_1_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_120;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_120;
  reg reg_act_config_inst_counter_enexo_120;
  reg reg_act_regs_data_3_2_enexo_3;
  reg reg_act_regs_data_0_2_2_enexo_3;
  reg reg_act_regs_data_1_2_2_enexo_3;
  reg reg_act_regs_data_3_2_2_enexo_3;
  reg reg_act_regs_data_2_2_2_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_121;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_121;
  reg reg_act_config_inst_counter_enexo_121;
  reg reg_act_regs_data_3_2_enexo_4;
  reg reg_act_regs_data_3_2_3_enexo_3;
  reg reg_act_regs_data_2_2_3_enexo_3;
  reg reg_act_regs_data_0_2_3_enexo_3;
  reg reg_act_regs_data_1_2_3_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_122;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_122;
  reg reg_act_regs_data_2_1_1_enexo_3;
  reg reg_act_config_inst_counter_enexo_122;
  reg reg_act_regs_data_3_1_1_enexo_3;
  reg reg_act_regs_data_2_1_enexo_2;
  reg reg_act_regs_data_0_1_1_enexo_3;
  reg reg_act_regs_data_1_1_1_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_123;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_123;
  reg reg_act_config_inst_counter_enexo_123;
  reg reg_act_regs_data_1_1_2_enexo_3;
  reg reg_act_regs_data_2_1_enexo_3;
  reg reg_act_regs_data_3_1_2_enexo_3;
  reg reg_act_regs_data_0_1_2_enexo_3;
  reg reg_act_regs_data_2_1_2_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_124;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_124;
  reg reg_act_config_inst_counter_enexo_124;
  reg reg_act_regs_data_0_1_3_enexo_3;
  reg reg_act_regs_data_2_1_enexo_4;
  reg reg_act_regs_data_3_1_3_enexo_3;
  reg reg_act_regs_data_1_1_3_enexo_3;
  reg reg_act_regs_data_2_1_3_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_125;
  reg reg_act_regs_data_3_0_1_enexo_3;
  reg reg_act_regs_data_3_0_enexo_2;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_125;
  reg reg_act_config_inst_counter_enexo_125;
  reg reg_act_regs_data_0_0_1_enexo_3;
  reg reg_act_regs_data_2_0_1_enexo_3;
  reg reg_act_regs_data_1_0_1_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_126;
  reg reg_act_regs_data_3_0_enexo_3;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_126;
  reg reg_act_config_inst_counter_enexo_126;
  reg reg_act_regs_data_3_0_2_enexo_3;
  reg reg_act_regs_data_0_0_2_enexo_3;
  reg reg_act_regs_data_1_0_2_enexo_3;
  reg reg_act_regs_data_2_0_2_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_127;
  reg reg_act_regs_data_3_0_enexo_4;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_127;
  reg reg_act_config_inst_counter_enexo_127;
  reg reg_act_regs_data_3_0_3_enexo_3;
  reg reg_act_regs_data_0_0_3_enexo_3;
  reg reg_act_regs_data_2_0_3_enexo_3;
  reg reg_act_regs_data_1_0_3_enexo_3;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_128;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_128;
  reg reg_act_config_inst_counter_enexo_128;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_129;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_129;
  reg reg_act_config_inst_counter_enexo_129;
  reg reg_act_regs_data_3_0_2_enexo_4;
  reg reg_act_regs_data_0_0_2_enexo_4;
  reg reg_act_regs_data_1_0_2_enexo_4;
  reg reg_act_regs_data_2_0_2_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_130;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_130;
  reg reg_act_config_inst_counter_enexo_130;
  reg reg_act_regs_data_3_0_3_enexo_4;
  reg reg_act_regs_data_0_0_3_enexo_4;
  reg reg_act_regs_data_2_0_3_enexo_4;
  reg reg_act_regs_data_1_0_3_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_131;
  reg reg_act_regs_data_3_0_1_enexo_4;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_131;
  reg reg_act_config_inst_counter_enexo_131;
  reg reg_act_regs_data_0_0_1_enexo_4;
  reg reg_act_regs_data_2_0_1_enexo_4;
  reg reg_act_regs_data_1_0_1_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_132;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_132;
  reg reg_act_config_inst_counter_enexo_132;
  reg reg_act_regs_data_1_1_2_enexo_4;
  reg reg_act_regs_data_3_1_2_enexo_4;
  reg reg_act_regs_data_0_1_2_enexo_4;
  reg reg_act_regs_data_2_1_2_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_133;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_133;
  reg reg_act_config_inst_counter_enexo_133;
  reg reg_act_regs_data_0_1_3_enexo_4;
  reg reg_act_regs_data_3_1_3_enexo_4;
  reg reg_act_regs_data_1_1_3_enexo_4;
  reg reg_act_regs_data_2_1_3_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_134;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_134;
  reg reg_act_regs_data_2_1_1_enexo_4;
  reg reg_act_config_inst_counter_enexo_134;
  reg reg_act_regs_data_3_1_1_enexo_4;
  reg reg_act_regs_data_0_1_1_enexo_4;
  reg reg_act_regs_data_1_1_1_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_135;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_135;
  reg reg_act_config_inst_counter_enexo_135;
  reg reg_act_regs_data_0_2_2_enexo_4;
  reg reg_act_regs_data_1_2_2_enexo_4;
  reg reg_act_regs_data_3_2_2_enexo_4;
  reg reg_act_regs_data_2_2_2_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_136;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_136;
  reg reg_act_config_inst_counter_enexo_136;
  reg reg_act_regs_data_3_2_3_enexo_4;
  reg reg_act_regs_data_2_2_3_enexo_4;
  reg reg_act_regs_data_0_2_3_enexo_4;
  reg reg_act_regs_data_1_2_3_enexo_4;
  reg reg_act_regs_data_2_2_1_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_137;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_137;
  reg reg_act_config_inst_counter_enexo_137;
  reg reg_act_regs_data_3_2_1_enexo_4;
  reg reg_act_regs_data_1_2_1_enexo_4;
  reg reg_act_regs_data_0_2_1_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_138;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_138;
  reg reg_act_config_inst_counter_enexo_138;
  reg reg_act_regs_data_0_3_2_enexo_4;
  reg reg_act_regs_data_1_3_2_enexo_4;
  reg reg_act_regs_data_3_3_2_enexo_4;
  reg reg_act_regs_data_2_3_2_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_139;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_139;
  reg reg_act_config_inst_counter_enexo_139;
  reg reg_act_regs_data_0_3_3_enexo_4;
  reg reg_act_regs_data_3_3_3_enexo_4;
  reg reg_act_regs_data_1_3_3_enexo_4;
  reg reg_act_regs_data_2_3_3_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_140;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_140;
  reg reg_act_config_inst_counter_enexo_140;
  reg reg_act_regs_data_0_3_1_enexo_4;
  reg reg_act_regs_data_3_3_1_enexo_4;
  reg reg_act_regs_data_1_3_1_enexo_4;
  reg reg_act_regs_data_2_3_1_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_141;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_141;
  reg reg_act_config_inst_counter_enexo_141;
  reg reg_act_regs_data_3_4_2_enexo_4;
  reg reg_act_regs_data_1_4_2_enexo_4;
  reg reg_act_regs_data_0_4_2_enexo_4;
  reg reg_act_regs_data_2_4_2_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_142;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_142;
  reg reg_act_config_inst_counter_enexo_142;
  reg reg_act_regs_data_0_4_3_enexo_4;
  reg reg_act_regs_data_1_4_3_enexo_4;
  reg reg_act_regs_data_3_4_3_enexo_4;
  reg reg_act_regs_data_2_4_3_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_143;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_143;
  reg reg_act_config_inst_counter_enexo_143;
  reg reg_act_regs_data_3_4_1_enexo_4;
  reg reg_act_regs_data_0_4_1_enexo_4;
  reg reg_act_regs_data_2_4_1_enexo_4;
  reg reg_act_regs_data_1_4_1_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_144;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_144;
  reg reg_act_config_inst_counter_enexo_144;
  reg reg_act_regs_data_2_5_2_enexo_4;
  reg reg_act_regs_data_1_5_2_enexo_4;
  reg reg_act_regs_data_3_5_2_enexo_4;
  reg reg_act_regs_data_0_5_2_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_145;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_145;
  reg reg_act_regs_data_0_5_3_enexo_4;
  reg reg_act_config_inst_counter_enexo_145;
  reg reg_act_regs_data_1_5_3_enexo_4;
  reg reg_act_regs_data_3_5_3_enexo_4;
  reg reg_act_regs_data_2_5_3_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_146;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_146;
  reg reg_act_config_inst_counter_enexo_146;
  reg reg_act_regs_data_3_5_1_enexo_4;
  reg reg_act_regs_data_0_5_1_enexo_4;
  reg reg_act_regs_data_1_5_1_enexo_4;
  reg reg_act_regs_data_2_5_1_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_147;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_147;
  reg reg_act_config_inst_counter_enexo_147;
  reg reg_act_regs_data_2_6_2_enexo_4;
  reg reg_act_regs_data_1_6_2_enexo_4;
  reg reg_act_regs_data_3_6_2_enexo_4;
  reg reg_act_regs_data_0_6_2_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_148;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_148;
  reg reg_act_config_inst_counter_enexo_148;
  reg reg_act_regs_data_2_6_3_enexo_4;
  reg reg_act_regs_data_3_6_3_enexo_4;
  reg reg_act_regs_data_0_6_3_enexo_4;
  reg reg_act_regs_data_1_6_3_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_149;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_149;
  reg reg_act_config_inst_counter_enexo_149;
  reg reg_act_regs_data_3_6_1_enexo_4;
  reg reg_act_regs_data_1_6_1_enexo_4;
  reg reg_act_regs_data_2_6_1_enexo_4;
  reg reg_act_regs_data_0_6_1_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_150;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_150;
  reg reg_act_config_inst_counter_enexo_150;
  reg reg_act_regs_data_0_7_2_enexo_4;
  reg reg_act_regs_data_2_7_2_enexo_4;
  reg reg_act_regs_data_3_7_2_enexo_4;
  reg reg_act_regs_data_1_7_2_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_151;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_151;
  reg reg_act_config_inst_counter_enexo_151;
  reg reg_act_regs_data_0_7_3_enexo_4;
  reg reg_act_regs_data_1_7_3_enexo_4;
  reg reg_act_regs_data_3_7_3_enexo_4;
  reg reg_act_regs_data_2_7_3_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_152;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_152;
  reg reg_act_config_inst_counter_enexo_152;
  reg reg_act_regs_data_3_7_1_enexo_4;
  reg reg_act_regs_data_1_7_1_enexo_4;
  reg reg_act_regs_data_0_7_1_enexo_4;
  reg reg_act_regs_data_2_7_1_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_153;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_153;
  reg reg_act_config_inst_counter_enexo_153;
  reg reg_act_regs_data_0_8_2_enexo_4;
  reg reg_act_regs_data_1_8_2_enexo_4;
  reg reg_act_regs_data_2_8_2_enexo_4;
  reg reg_act_regs_data_3_8_2_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_154;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_154;
  reg reg_act_config_inst_counter_enexo_154;
  reg reg_act_regs_data_0_8_3_enexo_4;
  reg reg_act_regs_data_2_8_3_enexo_4;
  reg reg_act_regs_data_1_8_3_enexo_4;
  reg reg_act_regs_data_3_8_3_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_155;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_155;
  reg reg_act_config_inst_counter_enexo_155;
  reg reg_act_regs_data_2_8_1_enexo_4;
  reg reg_act_regs_data_0_8_1_enexo_4;
  reg reg_act_regs_data_3_8_1_enexo_4;
  reg reg_act_regs_data_1_8_1_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_156;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_156;
  reg reg_act_config_inst_counter_enexo_156;
  reg reg_act_regs_data_0_9_2_enexo_4;
  reg reg_act_regs_data_2_9_2_enexo_4;
  reg reg_act_regs_data_1_9_2_enexo_4;
  reg reg_act_regs_data_3_9_2_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_157;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_157;
  reg reg_act_config_inst_counter_enexo_157;
  reg reg_act_regs_data_1_9_3_enexo_4;
  reg reg_act_regs_data_0_9_3_enexo_4;
  reg reg_act_regs_data_2_9_3_enexo_4;
  reg reg_act_regs_data_3_9_3_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_158;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_158;
  reg reg_act_config_inst_counter_enexo_158;
  reg reg_act_regs_data_1_9_1_enexo_4;
  reg reg_act_regs_data_3_9_1_enexo_4;
  reg reg_act_regs_data_0_9_1_enexo_4;
  reg reg_act_regs_data_2_9_1_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_159;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_159;
  reg reg_act_config_inst_counter_enexo_159;
  reg reg_act_regs_data_1_10_2_enexo_4;
  reg reg_act_regs_data_0_10_2_enexo_4;
  reg reg_act_regs_data_3_10_2_enexo_4;
  reg reg_act_regs_data_2_10_2_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_160;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_160;
  reg reg_act_config_inst_counter_enexo_160;
  reg reg_act_regs_data_3_10_3_enexo_4;
  reg reg_act_regs_data_0_10_3_enexo_4;
  reg reg_act_regs_data_2_10_3_enexo_4;
  reg reg_act_regs_data_1_10_3_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_161;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_161;
  reg reg_act_config_inst_counter_enexo_161;
  reg reg_act_regs_data_1_10_1_enexo_4;
  reg reg_act_regs_data_2_10_1_enexo_4;
  reg reg_act_regs_data_3_10_1_enexo_4;
  reg reg_act_regs_data_0_10_1_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_162;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_162;
  reg reg_act_config_inst_counter_enexo_162;
  reg reg_act_regs_data_2_11_2_enexo_4;
  reg reg_act_regs_data_0_11_2_enexo_4;
  reg reg_act_regs_data_3_11_2_enexo_4;
  reg reg_act_regs_data_1_11_2_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_163;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_163;
  reg reg_act_config_inst_counter_enexo_163;
  reg reg_act_regs_data_0_11_3_enexo_4;
  reg reg_act_regs_data_1_11_3_enexo_4;
  reg reg_act_regs_data_2_11_3_enexo_4;
  reg reg_act_regs_data_3_11_3_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_164;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_164;
  reg reg_act_config_inst_counter_enexo_164;
  reg reg_act_regs_data_2_11_1_enexo_4;
  reg reg_act_regs_data_3_11_1_enexo_4;
  reg reg_act_regs_data_0_11_1_enexo_4;
  reg reg_act_regs_data_1_11_1_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_165;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_165;
  reg reg_act_regs_data_2_12_2_enexo_4;
  reg reg_act_config_inst_counter_enexo_165;
  reg reg_act_regs_data_0_12_2_enexo_4;
  reg reg_act_regs_data_3_12_2_enexo_4;
  reg reg_act_regs_data_1_12_2_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_166;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_166;
  reg reg_act_config_inst_counter_enexo_166;
  reg reg_act_regs_data_0_12_3_enexo_4;
  reg reg_act_regs_data_2_12_3_enexo_4;
  reg reg_act_regs_data_3_12_3_enexo_4;
  reg reg_act_regs_data_1_12_3_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_167;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_167;
  reg reg_act_config_inst_counter_enexo_167;
  reg reg_act_regs_data_2_12_1_enexo_4;
  reg reg_act_regs_data_0_12_1_enexo_4;
  reg reg_act_regs_data_1_12_1_enexo_4;
  reg reg_act_regs_data_3_12_1_enexo_4;
  reg reg_act_regs_data_3_13_2_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_168;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_168;
  reg reg_act_regs_data_0_13_2_enexo_4;
  reg reg_act_config_inst_counter_enexo_168;
  reg reg_act_regs_data_1_13_2_enexo_4;
  reg reg_act_regs_data_2_13_2_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_169;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_169;
  reg reg_act_config_inst_counter_enexo_169;
  reg reg_act_regs_data_2_13_3_enexo_4;
  reg reg_act_regs_data_3_13_3_enexo_4;
  reg reg_act_regs_data_1_13_3_enexo_4;
  reg reg_act_regs_data_0_13_3_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_170;
  reg reg_act_regs_data_1_13_1_enexo_4;
  reg reg_act_regs_data_2_13_1_enexo_4;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_170;
  reg reg_act_config_inst_counter_enexo_170;
  reg reg_act_regs_data_0_13_1_enexo_4;
  reg reg_act_regs_data_3_13_1_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_171;
  reg reg_act_regs_data_0_14_2_enexo_4;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_171;
  reg reg_act_config_inst_counter_enexo_171;
  reg reg_act_regs_data_2_14_2_enexo_4;
  reg reg_act_regs_data_3_14_2_enexo_4;
  reg reg_act_regs_data_1_14_2_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_172;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_172;
  reg reg_act_config_inst_counter_enexo_172;
  reg reg_act_regs_data_0_14_3_enexo_4;
  reg reg_act_regs_data_2_14_3_enexo_4;
  reg reg_act_regs_data_3_14_3_enexo_4;
  reg reg_act_regs_data_1_14_3_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_173;
  reg reg_act_regs_data_1_14_1_enexo_4;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_173;
  reg reg_act_config_inst_counter_enexo_173;
  reg reg_act_regs_data_2_14_1_enexo_4;
  reg reg_act_regs_data_3_14_1_enexo_4;
  reg reg_act_regs_data_0_14_1_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_174;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_174;
  reg reg_act_config_inst_counter_enexo_174;
  reg reg_act_regs_data_3_15_2_enexo_4;
  reg reg_act_regs_data_2_15_2_enexo_4;
  reg reg_act_regs_data_0_15_2_enexo_4;
  reg reg_act_regs_data_1_15_2_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_175;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_175;
  reg reg_act_regs_data_2_15_3_enexo_4;
  reg reg_act_config_inst_counter_enexo_175;
  reg reg_act_regs_data_0_15_3_enexo_4;
  reg reg_act_regs_data_1_15_3_enexo_4;
  reg reg_act_regs_data_3_15_3_enexo_4;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_176;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_176;
  reg reg_act_config_inst_counter_enexo_176;
  reg reg_act_regs_data_0_15_1_enexo_4;
  reg reg_act_regs_data_1_15_1_enexo_4;
  reg reg_act_regs_data_2_15_1_enexo_4;
  reg reg_act_regs_data_3_15_1_enexo_4;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo;
  reg reg_act_regs_data_3_15_sva_dfm_2_30_26_enexo_1;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo_1;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo_1;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo_1;
  reg reg_act_regs_data_3_15_sva_dfm_2_25_22_enexo_1;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo_1;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo_1;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo_1;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo_1;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo_1;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo_1;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo_1;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo_1;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo_1;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo_1;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_1;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_1;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo_1;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo_1;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo_1;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo_2;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo_2;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo_2;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo_2;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo_2;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo_2;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo_2;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo_2;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo_2;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo_2;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo_2;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo_2;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo_2;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_2;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_2;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo_2;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo_2;
  reg reg_act_regs_data_3_15_sva_dfm_2_21_0_enexo_1;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo_2;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo_3;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo_3;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo_3;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo_3;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo_3;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo_3;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo_3;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo_3;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo_3;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo_3;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo_3;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo_3;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo_3;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_3;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_3;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo_3;
  reg reg_act_regs_data_3_14_sva_dfm_2_30_26_enexo_1;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo_3;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo_3;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo_4;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo_4;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo_4;
  reg reg_act_regs_data_3_14_sva_dfm_2_25_22_enexo_1;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo_4;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo_4;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo_4;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo_4;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo_4;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo_4;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo_4;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo_4;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo_4;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo_4;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_4;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_4;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo_4;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo_4;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo_4;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo_5;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo_5;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo_5;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo_5;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo_5;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo_5;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo_5;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo_5;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo_5;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo_5;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo_5;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo_5;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo_5;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_5;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_5;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo_5;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo_5;
  reg reg_act_regs_data_3_14_sva_dfm_2_21_0_enexo_1;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo_5;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo_6;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo_6;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo_6;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo_6;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo_6;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo_6;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo_6;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo_6;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo_6;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo_6;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo_6;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo_6;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo_6;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_6;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_6;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo_6;
  reg reg_act_regs_data_3_13_sva_dfm_2_30_26_enexo_1;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo_6;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo_6;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo_7;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo_7;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo_7;
  reg reg_act_regs_data_3_13_sva_dfm_2_25_22_enexo_1;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo_7;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo_7;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo_7;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo_7;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo_7;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo_7;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo_7;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo_7;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo_7;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo_7;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_7;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_7;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo_7;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo_7;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo_7;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo_8;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo_8;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo_8;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo_8;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo_8;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo_8;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo_8;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo_8;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo_8;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo_8;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo_8;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo_8;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo_8;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_8;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_8;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo_8;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo_8;
  reg reg_act_regs_data_3_13_sva_dfm_2_21_0_enexo_1;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo_8;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo_9;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo_9;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo_9;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo_9;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo_9;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo_9;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo_9;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo_9;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo_9;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo_9;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo_9;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo_9;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo_9;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_9;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_9;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo_9;
  reg reg_act_regs_data_3_12_sva_dfm_2_30_26_enexo_1;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo_9;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo_9;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo_10;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo_10;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo_10;
  reg reg_act_regs_data_3_12_sva_dfm_2_25_22_enexo_1;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo_10;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo_10;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo_10;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo_10;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo_10;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo_10;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo_10;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo_10;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo_10;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo_10;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_10;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_10;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo_10;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo_10;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo_10;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo_11;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo_11;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo_11;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo_11;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo_11;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo_11;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo_11;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo_11;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo_11;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo_11;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo_11;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo_11;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo_11;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_11;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_11;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo_11;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo_11;
  reg reg_act_regs_data_3_12_sva_dfm_2_21_0_enexo_1;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo_11;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo_12;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo_12;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo_12;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo_12;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo_12;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo_12;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo_12;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo_12;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo_12;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo_12;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo_12;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo_12;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo_12;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_12;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_12;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo_12;
  reg reg_act_regs_data_3_11_sva_dfm_2_30_26_enexo_1;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo_12;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo_12;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo_13;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo_13;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo_13;
  reg reg_act_regs_data_3_11_sva_dfm_2_25_22_enexo_1;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo_13;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo_13;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo_13;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo_13;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo_13;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo_13;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo_13;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo_13;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo_13;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo_13;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_13;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_13;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo_13;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo_13;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo_13;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo_14;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo_14;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo_14;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo_14;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo_14;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo_14;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo_14;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo_14;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo_14;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo_14;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo_14;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo_14;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo_14;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_14;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_14;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo_14;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo_14;
  reg reg_act_regs_data_3_11_sva_dfm_2_21_0_enexo_1;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo_14;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo_15;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo_15;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo_15;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo_15;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo_15;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo_15;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo_15;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo_15;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo_15;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo_15;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo_15;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo_15;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo_15;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_15;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_15;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo_15;
  reg reg_act_regs_data_3_10_sva_dfm_2_30_26_enexo_1;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo_15;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo_15;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo_16;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo_16;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo_16;
  reg reg_act_regs_data_3_10_sva_dfm_2_25_22_enexo_1;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo_16;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo_16;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo_16;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo_16;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo_16;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo_16;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo_16;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo_16;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo_16;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo_16;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_16;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_16;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo_16;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo_16;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo_16;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo_17;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo_17;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo_17;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo_17;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo_17;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo_17;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo_17;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo_17;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo_17;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo_17;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo_17;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo_17;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo_17;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_17;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_17;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo_17;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo_17;
  reg reg_act_regs_data_3_10_sva_dfm_2_21_0_enexo_1;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo_17;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo_18;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo_18;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo_18;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo_18;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo_18;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo_18;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo_18;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo_18;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo_18;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo_18;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo_18;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo_18;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo_18;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_18;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_18;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo_18;
  reg reg_act_regs_data_3_9_sva_dfm_2_30_26_enexo_1;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo_18;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo_18;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo_19;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo_19;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo_19;
  reg reg_act_regs_data_3_9_sva_dfm_2_25_22_enexo_1;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo_19;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo_19;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo_19;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo_19;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo_19;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo_19;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo_19;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo_19;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo_19;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo_19;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_19;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_19;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo_19;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo_19;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo_19;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo_20;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo_20;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo_20;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo_20;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo_20;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo_20;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo_20;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo_20;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo_20;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo_20;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo_20;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo_20;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo_20;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_20;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_20;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo_20;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo_20;
  reg reg_act_regs_data_3_9_sva_dfm_2_21_0_enexo_1;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo_20;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo_21;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo_21;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo_21;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo_21;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo_21;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo_21;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo_21;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo_21;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo_21;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo_21;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo_21;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo_21;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo_21;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_21;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_21;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo_21;
  reg reg_act_regs_data_3_8_sva_dfm_2_30_26_enexo_1;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo_21;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo_21;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo_22;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo_22;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo_22;
  reg reg_act_regs_data_3_8_sva_dfm_2_25_22_enexo_1;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo_22;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo_22;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo_22;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo_22;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo_22;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo_22;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo_22;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo_22;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo_22;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo_22;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_22;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_22;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo_22;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo_22;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo_22;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo_23;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo_23;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo_23;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo_23;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo_23;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo_23;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo_23;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo_23;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo_23;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo_23;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo_23;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo_23;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo_23;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_23;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_23;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo_23;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo_23;
  reg reg_act_regs_data_3_8_sva_dfm_2_21_0_enexo_1;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo_23;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo_24;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo_24;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo_24;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo_24;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo_24;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo_24;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo_24;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo_24;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo_24;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo_24;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo_24;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo_24;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo_24;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_24;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_24;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo_24;
  reg reg_act_regs_data_3_7_sva_dfm_2_30_26_enexo_1;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo_24;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo_24;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo_25;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo_25;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo_25;
  reg reg_act_regs_data_3_7_sva_dfm_2_25_22_enexo_1;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo_25;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo_25;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo_25;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo_25;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo_25;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo_25;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo_25;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo_25;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo_25;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo_25;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_25;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_25;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo_25;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo_25;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo_25;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo_26;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo_26;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo_26;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo_26;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo_26;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo_26;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo_26;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo_26;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo_26;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo_26;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo_26;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo_26;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo_26;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_26;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_26;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo_26;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo_26;
  reg reg_act_regs_data_3_7_sva_dfm_2_21_0_enexo_1;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo_26;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo_27;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo_27;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo_27;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo_27;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo_27;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo_27;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo_27;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo_27;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo_27;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo_27;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo_27;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo_27;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo_27;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_27;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_27;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo_27;
  reg reg_act_regs_data_3_6_sva_dfm_2_30_26_enexo_1;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo_27;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo_27;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo_28;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo_28;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo_28;
  reg reg_act_regs_data_3_6_sva_dfm_2_25_22_enexo_1;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo_28;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo_28;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo_28;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo_28;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo_28;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo_28;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo_28;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo_28;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo_28;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo_28;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_28;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_28;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo_28;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo_28;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo_28;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo_29;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo_29;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo_29;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo_29;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo_29;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo_29;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo_29;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo_29;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo_29;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo_29;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo_29;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo_29;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo_29;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_29;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_29;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo_29;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo_29;
  reg reg_act_regs_data_3_6_sva_dfm_2_21_0_enexo_1;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo_29;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo_30;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo_30;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo_30;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo_30;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo_30;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo_30;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo_30;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo_30;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo_30;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo_30;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo_30;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo_30;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo_30;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_30;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_30;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo_30;
  reg reg_act_regs_data_3_5_sva_dfm_2_30_26_enexo_1;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo_30;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo_30;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo_31;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo_31;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo_31;
  reg reg_act_regs_data_3_5_sva_dfm_2_25_22_enexo_1;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo_31;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo_31;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo_31;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo_31;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo_31;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo_31;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo_31;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo_31;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo_31;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo_31;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_31;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_31;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo_31;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo_31;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo_31;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo_32;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo_32;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo_32;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo_32;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo_32;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo_32;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo_32;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo_32;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo_32;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo_32;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo_32;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo_32;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo_32;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_32;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_32;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo_32;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo_32;
  reg reg_act_regs_data_3_5_sva_dfm_2_21_0_enexo_1;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo_32;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo_33;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo_33;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo_33;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo_33;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo_33;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo_33;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo_33;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo_33;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo_33;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo_33;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo_33;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo_33;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo_33;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_33;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_33;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo_33;
  reg reg_act_regs_data_3_4_sva_dfm_2_30_26_enexo_1;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo_33;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo_33;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo_34;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo_34;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo_34;
  reg reg_act_regs_data_3_4_sva_dfm_2_25_22_enexo_1;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo_34;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo_34;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo_34;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo_34;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo_34;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo_34;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo_34;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo_34;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo_34;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo_34;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_34;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_34;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo_34;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo_34;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo_34;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo_35;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo_35;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo_35;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo_35;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo_35;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo_35;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo_35;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo_35;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo_35;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo_35;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo_35;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo_35;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo_35;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_35;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_35;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo_35;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo_35;
  reg reg_act_regs_data_3_4_sva_dfm_2_21_0_enexo_1;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo_35;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo_36;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo_36;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo_36;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo_36;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo_36;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo_36;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo_36;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo_36;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo_36;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo_36;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo_36;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo_36;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo_36;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_36;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_36;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo_36;
  reg reg_act_regs_data_3_3_sva_dfm_2_30_26_enexo_1;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo_36;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo_36;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo_37;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo_37;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo_37;
  reg reg_act_regs_data_3_3_sva_dfm_2_25_22_enexo_1;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo_37;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo_37;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo_37;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo_37;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo_37;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo_37;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo_37;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo_37;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo_37;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo_37;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_37;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_37;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo_37;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo_37;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo_37;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo_38;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo_38;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo_38;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo_38;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo_38;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo_38;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo_38;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo_38;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo_38;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo_38;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo_38;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo_38;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo_38;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_38;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_38;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo_38;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo_38;
  reg reg_act_regs_data_3_3_sva_dfm_2_21_0_enexo_1;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo_38;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo_39;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo_39;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo_39;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo_39;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo_39;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo_39;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo_39;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo_39;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo_39;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo_39;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo_39;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo_39;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo_39;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_39;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_39;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo_39;
  reg reg_act_regs_data_3_2_sva_dfm_2_30_26_enexo_1;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo_39;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo_39;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo_40;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo_40;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo_40;
  reg reg_act_regs_data_3_2_sva_dfm_2_25_22_enexo_1;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo_40;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo_40;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo_40;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo_40;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo_40;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo_40;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo_40;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo_40;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo_40;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo_40;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_40;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_40;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo_40;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo_40;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo_40;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo_41;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo_41;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo_41;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo_41;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo_41;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo_41;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo_41;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo_41;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo_41;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo_41;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo_41;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo_41;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo_41;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_41;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_41;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo_41;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo_41;
  reg reg_act_regs_data_3_2_sva_dfm_2_21_0_enexo_1;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo_41;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo_42;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo_42;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo_42;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo_42;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo_42;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo_42;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo_42;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo_42;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo_42;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo_42;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo_42;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo_42;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo_42;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_42;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_42;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo_42;
  reg reg_act_regs_data_3_1_sva_dfm_2_30_26_enexo_1;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo_42;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo_42;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo_43;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo_43;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo_43;
  reg reg_act_regs_data_3_1_sva_dfm_2_25_22_enexo_1;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo_43;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo_43;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo_43;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo_43;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo_43;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo_43;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo_43;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo_43;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo_43;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo_43;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_43;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_43;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo_43;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo_43;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo_43;
  reg reg_act_port_read_out_data_0_5_sva_dfm_enexo_44;
  reg reg_act_port_read_out_data_0_6_sva_dfm_enexo_44;
  reg reg_act_port_read_out_data_0_13_sva_dfm_enexo_44;
  reg reg_act_port_read_out_data_0_10_sva_dfm_enexo_44;
  reg reg_act_port_read_out_data_0_11_sva_dfm_enexo_44;
  reg reg_act_port_read_out_data_0_15_sva_dfm_enexo_44;
  reg reg_act_port_read_out_data_0_7_sva_dfm_enexo_44;
  reg reg_act_port_read_out_data_0_8_sva_dfm_enexo_44;
  reg reg_act_port_read_out_data_0_0_sva_dfm_enexo_44;
  reg reg_act_port_read_out_data_0_12_sva_dfm_enexo_44;
  reg reg_act_port_read_out_data_0_3_sva_dfm_enexo_44;
  reg reg_act_port_read_out_data_0_9_sva_dfm_enexo_44;
  reg reg_act_port_read_out_data_0_1_sva_dfm_enexo_44;
  reg reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_44;
  reg reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_44;
  reg reg_act_port_read_out_data_0_14_sva_dfm_enexo_44;
  reg reg_act_port_read_out_data_0_4_sva_dfm_enexo_44;
  reg reg_act_regs_data_3_1_sva_dfm_2_21_0_enexo_1;
  reg reg_act_port_read_out_data_0_2_sva_dfm_enexo_44;
  reg reg_is_start_enexo_174;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_174;
  reg reg_act_regs_data_0_13_sva_8_30_26_enexo_1;
  reg reg_ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_1_30_26_enexo;
  reg reg_act_regs_data_0_13_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_174;
  reg reg_is_start_enexo_175;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_175;
  reg reg_ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_1_25_22_enexo;
  reg reg_act_regs_data_0_13_sva_8_25_22_enexo_1;
  reg reg_act_regs_data_0_13_sva_dfm_2_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_175;
  reg reg_is_start_enexo_176;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_176;
  reg reg_act_regs_data_0_13_sva_8_21_0_enexo_1;
  reg reg_Silu_for_16_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo;
  reg reg_act_regs_data_0_13_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_176;
  reg reg_is_start_enexo_177;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_177;
  reg reg_act_regs_data_0_12_sva_8_30_26_enexo_1;
  reg reg_ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_1_30_26_enexo;
  reg reg_act_regs_data_0_12_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_177;
  reg reg_is_start_enexo_178;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_178;
  reg reg_ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_1_25_22_enexo;
  reg reg_act_regs_data_0_12_sva_8_25_22_enexo_1;
  reg reg_act_regs_data_0_12_sva_dfm_2_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_178;
  reg reg_is_start_enexo_179;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_179;
  reg reg_act_regs_data_0_12_sva_8_21_0_enexo_1;
  reg reg_Silu_for_15_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo;
  reg reg_act_regs_data_0_12_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_179;
  reg reg_is_start_enexo_180;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_180;
  reg reg_act_regs_data_0_11_sva_8_30_26_enexo_1;
  reg reg_ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_1_30_26_enexo;
  reg reg_act_regs_data_0_11_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_180;
  reg reg_is_start_enexo_181;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_181;
  reg reg_ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_1_25_22_enexo;
  reg reg_act_regs_data_0_11_sva_8_25_22_enexo_1;
  reg reg_act_regs_data_0_11_sva_dfm_2_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_181;
  reg reg_is_start_enexo_182;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_182;
  reg reg_act_regs_data_0_11_sva_8_21_0_enexo_1;
  reg reg_act_regs_data_0_11_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_182;
  reg reg_Silu_for_14_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo;
  reg reg_is_start_enexo_183;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_183;
  reg reg_act_regs_data_0_10_sva_8_30_26_enexo_1;
  reg reg_ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_1_30_26_enexo;
  reg reg_act_regs_data_0_10_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_183;
  reg reg_is_start_enexo_184;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_184;
  reg reg_ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_1_25_22_enexo;
  reg reg_act_regs_data_0_10_sva_8_25_22_enexo_1;
  reg reg_act_regs_data_0_10_sva_dfm_2_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_184;
  reg reg_is_start_enexo_185;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_185;
  reg reg_act_regs_data_0_10_sva_8_21_0_enexo_1;
  reg reg_act_regs_data_0_10_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_185;
  reg reg_Silu_for_13_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo;
  reg reg_is_start_enexo_186;
  reg reg_act_regs_data_0_1_sva_8_30_26_enexo_1;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_186;
  reg reg_rva_out_reg_data_71_64_sva_dfm_6_1_enexo;
  reg reg_act_regs_data_0_1_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_186;
  reg reg_is_start_enexo_187;
  reg reg_act_regs_data_0_1_sva_8_25_22_enexo_1;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_187;
  reg reg_rva_out_reg_data_39_32_sva_dfm_6_1_enexo;
  reg reg_act_regs_data_0_1_sva_dfm_2_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_187;
  reg reg_is_start_enexo_188;
  reg reg_act_regs_data_0_1_sva_8_21_0_enexo_1;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_188;
  reg reg_act_regs_data_0_1_sva_dfm_2_21_0_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_188;
  reg reg_Silu_for_12_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo;
  reg reg_ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_1_30_26_enexo;
  reg reg_is_start_enexo_189;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_189;
  reg reg_act_regs_data_0_0_sva_8_30_26_enexo_1;
  reg reg_act_regs_data_0_0_sva_dfm_2_30_26_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_189;
  reg reg_is_start_enexo_190;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_190;
  reg reg_rva_out_reg_data_29_24_sva_dfm_6_1_enexo;
  reg reg_act_regs_data_0_0_sva_8_25_22_enexo_1;
  reg reg_act_regs_data_0_0_sva_dfm_2_25_22_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_190;
  reg reg_is_start_enexo_191;
  reg reg_act_config_is_zero_first_sva_dfm_4_enexo_191;
  reg reg_act_regs_data_0_0_sva_8_21_0_enexo_1;
  reg reg_act_regs_data_0_0_sva_dfm_2_21_0_enexo;
  reg reg_Silu_for_11_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo;
  reg reg_w_load_lpi_1_dfm_1_enexo_191;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_177;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_177;
  reg reg_act_config_inst_counter_enexo_177;
  reg reg_act_regs_data_3_0_2_enexo_5;
  reg reg_act_regs_data_0_0_2_enexo_5;
  reg reg_act_regs_data_1_0_2_enexo_5;
  reg reg_act_regs_data_2_0_2_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_178;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_178;
  reg reg_act_config_inst_counter_enexo_178;
  reg reg_act_regs_data_3_0_3_enexo_5;
  reg reg_act_regs_data_0_0_3_enexo_5;
  reg reg_act_regs_data_2_0_3_enexo_5;
  reg reg_act_regs_data_1_0_3_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_179;
  reg reg_act_regs_data_3_0_1_enexo_5;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_179;
  reg reg_act_config_inst_counter_enexo_179;
  reg reg_act_regs_data_0_0_1_enexo_5;
  reg reg_act_regs_data_2_0_1_enexo_5;
  reg reg_act_regs_data_1_0_1_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_180;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_180;
  reg reg_act_config_inst_counter_enexo_180;
  reg reg_act_regs_data_1_1_2_enexo_5;
  reg reg_act_regs_data_3_1_2_enexo_5;
  reg reg_act_regs_data_0_1_2_enexo_5;
  reg reg_act_regs_data_2_1_2_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_181;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_181;
  reg reg_act_config_inst_counter_enexo_181;
  reg reg_act_regs_data_0_1_3_enexo_5;
  reg reg_act_regs_data_3_1_3_enexo_5;
  reg reg_act_regs_data_1_1_3_enexo_5;
  reg reg_act_regs_data_2_1_3_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_182;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_182;
  reg reg_act_regs_data_2_1_1_enexo_5;
  reg reg_act_config_inst_counter_enexo_182;
  reg reg_act_regs_data_3_1_1_enexo_5;
  reg reg_act_regs_data_0_1_1_enexo_5;
  reg reg_act_regs_data_1_1_1_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_183;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_183;
  reg reg_act_config_inst_counter_enexo_183;
  reg reg_act_regs_data_0_2_2_enexo_5;
  reg reg_act_regs_data_1_2_2_enexo_5;
  reg reg_act_regs_data_3_2_2_enexo_5;
  reg reg_act_regs_data_2_2_2_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_184;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_184;
  reg reg_act_config_inst_counter_enexo_184;
  reg reg_act_regs_data_3_2_3_enexo_5;
  reg reg_act_regs_data_2_2_3_enexo_5;
  reg reg_act_regs_data_0_2_3_enexo_5;
  reg reg_act_regs_data_1_2_3_enexo_5;
  reg reg_act_regs_data_2_2_1_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_185;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_185;
  reg reg_act_config_inst_counter_enexo_185;
  reg reg_act_regs_data_3_2_1_enexo_5;
  reg reg_act_regs_data_1_2_1_enexo_5;
  reg reg_act_regs_data_0_2_1_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_186;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_186;
  reg reg_act_config_inst_counter_enexo_186;
  reg reg_act_regs_data_0_3_2_enexo_5;
  reg reg_act_regs_data_1_3_2_enexo_5;
  reg reg_act_regs_data_3_3_2_enexo_5;
  reg reg_act_regs_data_2_3_2_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_187;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_187;
  reg reg_act_config_inst_counter_enexo_187;
  reg reg_act_regs_data_0_3_3_enexo_5;
  reg reg_act_regs_data_3_3_3_enexo_5;
  reg reg_act_regs_data_1_3_3_enexo_5;
  reg reg_act_regs_data_2_3_3_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_188;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_188;
  reg reg_act_config_inst_counter_enexo_188;
  reg reg_act_regs_data_0_3_1_enexo_5;
  reg reg_act_regs_data_3_3_1_enexo_5;
  reg reg_act_regs_data_1_3_1_enexo_5;
  reg reg_act_regs_data_2_3_1_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_189;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_189;
  reg reg_act_config_inst_counter_enexo_189;
  reg reg_act_regs_data_3_4_2_enexo_5;
  reg reg_act_regs_data_1_4_2_enexo_5;
  reg reg_act_regs_data_0_4_2_enexo_5;
  reg reg_act_regs_data_2_4_2_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_190;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_190;
  reg reg_act_config_inst_counter_enexo_190;
  reg reg_act_regs_data_0_4_3_enexo_5;
  reg reg_act_regs_data_1_4_3_enexo_5;
  reg reg_act_regs_data_3_4_3_enexo_5;
  reg reg_act_regs_data_2_4_3_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_191;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_191;
  reg reg_act_config_inst_counter_enexo_191;
  reg reg_act_regs_data_3_4_1_enexo_5;
  reg reg_act_regs_data_0_4_1_enexo_5;
  reg reg_act_regs_data_2_4_1_enexo_5;
  reg reg_act_regs_data_1_4_1_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_192;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_192;
  reg reg_act_config_inst_counter_enexo_192;
  reg reg_act_regs_data_2_5_2_enexo_5;
  reg reg_act_regs_data_1_5_2_enexo_5;
  reg reg_act_regs_data_3_5_2_enexo_5;
  reg reg_act_regs_data_0_5_2_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_193;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_193;
  reg reg_act_regs_data_0_5_3_enexo_5;
  reg reg_act_config_inst_counter_enexo_193;
  reg reg_act_regs_data_1_5_3_enexo_5;
  reg reg_act_regs_data_3_5_3_enexo_5;
  reg reg_act_regs_data_2_5_3_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_194;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_194;
  reg reg_act_config_inst_counter_enexo_194;
  reg reg_act_regs_data_3_5_1_enexo_5;
  reg reg_act_regs_data_0_5_1_enexo_5;
  reg reg_act_regs_data_1_5_1_enexo_5;
  reg reg_act_regs_data_2_5_1_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_195;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_195;
  reg reg_act_config_inst_counter_enexo_195;
  reg reg_act_regs_data_2_6_2_enexo_5;
  reg reg_act_regs_data_1_6_2_enexo_5;
  reg reg_act_regs_data_3_6_2_enexo_5;
  reg reg_act_regs_data_0_6_2_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_196;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_196;
  reg reg_act_config_inst_counter_enexo_196;
  reg reg_act_regs_data_2_6_3_enexo_5;
  reg reg_act_regs_data_3_6_3_enexo_5;
  reg reg_act_regs_data_0_6_3_enexo_5;
  reg reg_act_regs_data_1_6_3_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_197;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_197;
  reg reg_act_config_inst_counter_enexo_197;
  reg reg_act_regs_data_3_6_1_enexo_5;
  reg reg_act_regs_data_1_6_1_enexo_5;
  reg reg_act_regs_data_2_6_1_enexo_5;
  reg reg_act_regs_data_0_6_1_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_198;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_198;
  reg reg_act_config_inst_counter_enexo_198;
  reg reg_act_regs_data_0_7_2_enexo_5;
  reg reg_act_regs_data_2_7_2_enexo_5;
  reg reg_act_regs_data_3_7_2_enexo_5;
  reg reg_act_regs_data_1_7_2_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_199;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_199;
  reg reg_act_config_inst_counter_enexo_199;
  reg reg_act_regs_data_0_7_3_enexo_5;
  reg reg_act_regs_data_1_7_3_enexo_5;
  reg reg_act_regs_data_3_7_3_enexo_5;
  reg reg_act_regs_data_2_7_3_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_200;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_200;
  reg reg_act_config_inst_counter_enexo_200;
  reg reg_act_regs_data_3_7_1_enexo_5;
  reg reg_act_regs_data_1_7_1_enexo_5;
  reg reg_act_regs_data_0_7_1_enexo_5;
  reg reg_act_regs_data_2_7_1_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_201;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_201;
  reg reg_act_config_inst_counter_enexo_201;
  reg reg_act_regs_data_0_8_2_enexo_5;
  reg reg_act_regs_data_1_8_2_enexo_5;
  reg reg_act_regs_data_2_8_2_enexo_5;
  reg reg_act_regs_data_3_8_2_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_202;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_202;
  reg reg_act_config_inst_counter_enexo_202;
  reg reg_act_regs_data_0_8_3_enexo_5;
  reg reg_act_regs_data_2_8_3_enexo_5;
  reg reg_act_regs_data_1_8_3_enexo_5;
  reg reg_act_regs_data_3_8_3_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_203;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_203;
  reg reg_act_config_inst_counter_enexo_203;
  reg reg_act_regs_data_2_8_1_enexo_5;
  reg reg_act_regs_data_0_8_1_enexo_5;
  reg reg_act_regs_data_3_8_1_enexo_5;
  reg reg_act_regs_data_1_8_1_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_204;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_204;
  reg reg_act_config_inst_counter_enexo_204;
  reg reg_act_regs_data_0_9_2_enexo_5;
  reg reg_act_regs_data_2_9_2_enexo_5;
  reg reg_act_regs_data_1_9_2_enexo_5;
  reg reg_act_regs_data_3_9_2_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_205;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_205;
  reg reg_act_config_inst_counter_enexo_205;
  reg reg_act_regs_data_1_9_3_enexo_5;
  reg reg_act_regs_data_0_9_3_enexo_5;
  reg reg_act_regs_data_2_9_3_enexo_5;
  reg reg_act_regs_data_3_9_3_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_206;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_206;
  reg reg_act_config_inst_counter_enexo_206;
  reg reg_act_regs_data_1_9_1_enexo_5;
  reg reg_act_regs_data_3_9_1_enexo_5;
  reg reg_act_regs_data_0_9_1_enexo_5;
  reg reg_act_regs_data_2_9_1_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_207;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_207;
  reg reg_act_config_inst_counter_enexo_207;
  reg reg_act_regs_data_1_10_2_enexo_5;
  reg reg_act_regs_data_0_10_2_enexo_5;
  reg reg_act_regs_data_3_10_2_enexo_5;
  reg reg_act_regs_data_2_10_2_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_208;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_208;
  reg reg_act_config_inst_counter_enexo_208;
  reg reg_act_regs_data_3_10_3_enexo_5;
  reg reg_act_regs_data_0_10_3_enexo_5;
  reg reg_act_regs_data_2_10_3_enexo_5;
  reg reg_act_regs_data_1_10_3_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_209;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_209;
  reg reg_act_config_inst_counter_enexo_209;
  reg reg_act_regs_data_1_10_1_enexo_5;
  reg reg_act_regs_data_2_10_1_enexo_5;
  reg reg_act_regs_data_3_10_1_enexo_5;
  reg reg_act_regs_data_0_10_1_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_210;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_210;
  reg reg_act_config_inst_counter_enexo_210;
  reg reg_act_regs_data_2_11_2_enexo_5;
  reg reg_act_regs_data_0_11_2_enexo_5;
  reg reg_act_regs_data_3_11_2_enexo_5;
  reg reg_act_regs_data_1_11_2_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_211;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_211;
  reg reg_act_config_inst_counter_enexo_211;
  reg reg_act_regs_data_0_11_3_enexo_5;
  reg reg_act_regs_data_1_11_3_enexo_5;
  reg reg_act_regs_data_2_11_3_enexo_5;
  reg reg_act_regs_data_3_11_3_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_212;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_212;
  reg reg_act_config_inst_counter_enexo_212;
  reg reg_act_regs_data_2_11_1_enexo_5;
  reg reg_act_regs_data_3_11_1_enexo_5;
  reg reg_act_regs_data_0_11_1_enexo_5;
  reg reg_act_regs_data_1_11_1_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_213;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_213;
  reg reg_act_regs_data_2_12_2_enexo_5;
  reg reg_act_config_inst_counter_enexo_213;
  reg reg_act_regs_data_0_12_2_enexo_5;
  reg reg_act_regs_data_3_12_2_enexo_5;
  reg reg_act_regs_data_1_12_2_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_214;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_214;
  reg reg_act_config_inst_counter_enexo_214;
  reg reg_act_regs_data_0_12_3_enexo_5;
  reg reg_act_regs_data_2_12_3_enexo_5;
  reg reg_act_regs_data_3_12_3_enexo_5;
  reg reg_act_regs_data_1_12_3_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_215;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_215;
  reg reg_act_config_inst_counter_enexo_215;
  reg reg_act_regs_data_2_12_1_enexo_5;
  reg reg_act_regs_data_0_12_1_enexo_5;
  reg reg_act_regs_data_1_12_1_enexo_5;
  reg reg_act_regs_data_3_12_1_enexo_5;
  reg reg_act_regs_data_3_13_2_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_216;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_216;
  reg reg_act_regs_data_0_13_2_enexo_5;
  reg reg_act_config_inst_counter_enexo_216;
  reg reg_act_regs_data_1_13_2_enexo_5;
  reg reg_act_regs_data_2_13_2_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_217;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_217;
  reg reg_act_config_inst_counter_enexo_217;
  reg reg_act_regs_data_2_13_3_enexo_5;
  reg reg_act_regs_data_3_13_3_enexo_5;
  reg reg_act_regs_data_1_13_3_enexo_5;
  reg reg_act_regs_data_0_13_3_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_218;
  reg reg_act_regs_data_1_13_1_enexo_5;
  reg reg_act_regs_data_2_13_1_enexo_5;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_218;
  reg reg_act_config_inst_counter_enexo_218;
  reg reg_act_regs_data_0_13_1_enexo_5;
  reg reg_act_regs_data_3_13_1_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_219;
  reg reg_act_regs_data_0_14_2_enexo_5;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_219;
  reg reg_act_config_inst_counter_enexo_219;
  reg reg_act_regs_data_2_14_2_enexo_5;
  reg reg_act_regs_data_3_14_2_enexo_5;
  reg reg_act_regs_data_1_14_2_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_220;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_220;
  reg reg_act_config_inst_counter_enexo_220;
  reg reg_act_regs_data_0_14_3_enexo_5;
  reg reg_act_regs_data_2_14_3_enexo_5;
  reg reg_act_regs_data_3_14_3_enexo_5;
  reg reg_act_regs_data_1_14_3_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_221;
  reg reg_act_regs_data_1_14_1_enexo_5;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_221;
  reg reg_act_config_inst_counter_enexo_221;
  reg reg_act_regs_data_2_14_1_enexo_5;
  reg reg_act_regs_data_3_14_1_enexo_5;
  reg reg_act_regs_data_0_14_1_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_222;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_222;
  reg reg_act_config_inst_counter_enexo_222;
  reg reg_act_regs_data_3_15_2_enexo_5;
  reg reg_act_regs_data_2_15_2_enexo_5;
  reg reg_act_regs_data_0_15_2_enexo_5;
  reg reg_act_regs_data_1_15_2_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_223;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_223;
  reg reg_act_regs_data_2_15_3_enexo_5;
  reg reg_act_config_inst_counter_enexo_223;
  reg reg_act_regs_data_0_15_3_enexo_5;
  reg reg_act_regs_data_1_15_3_enexo_5;
  reg reg_act_regs_data_3_15_3_enexo_5;
  reg reg_act_config_inst_regs_4_sva_dfm_5_enexo_224;
  reg reg_act_config_inst_regs_20_sva_dfm_6_enexo_224;
  reg reg_act_config_inst_counter_enexo_224;
  reg reg_act_regs_data_0_15_1_enexo_5;
  reg reg_act_regs_data_1_15_1_enexo_5;
  reg reg_act_regs_data_2_15_1_enexo_5;
  reg reg_act_regs_data_3_15_1_enexo_5;
  wire act_regs_data_and_2530_enex5;
  wire act_regs_data_and_2531_enex5;
  wire act_regs_data_and_2532_enex5;
  wire act_regs_data_and_2533_enex5;
  wire act_regs_data_and_2534_enex5;
  wire act_regs_data_and_2535_enex5;
  wire act_regs_data_and_2536_enex5;
  wire act_regs_data_and_2537_enex5;
  wire act_regs_data_and_2538_enex5;
  wire act_regs_data_and_2539_enex5;
  wire act_regs_data_and_2540_enex5;
  wire act_regs_data_and_2541_enex5;
  wire act_regs_data_and_2542_enex5;
  wire act_regs_data_and_2543_enex5;
  wire act_regs_data_and_2544_enex5;
  wire act_regs_data_and_2545_enex5;
  wire act_regs_data_and_2546_enex5;
  wire act_regs_data_and_2547_enex5;
  wire act_regs_data_and_2548_enex5;
  wire act_regs_data_and_2549_enex5;
  wire act_regs_data_and_2550_enex5;
  wire act_regs_data_and_2551_enex5;
  wire act_regs_data_and_2552_enex5;
  wire act_regs_data_and_2553_enex5;
  wire act_regs_data_and_2554_enex5;
  wire act_regs_data_and_2555_enex5;
  wire act_regs_data_and_2556_enex5;
  wire act_regs_data_and_2557_enex5;
  wire act_regs_data_and_2558_enex5;
  wire act_regs_data_and_2559_enex5;
  wire act_regs_data_and_2560_enex5;
  wire act_regs_data_and_2561_enex5;
  wire act_regs_data_and_2562_enex5;
  wire act_regs_data_and_2563_enex5;
  wire act_regs_data_and_2564_enex5;
  wire act_regs_data_and_2565_enex5;
  wire act_regs_data_and_2566_enex5;
  wire act_regs_data_and_2567_enex5;
  wire act_regs_data_and_2568_enex5;
  wire act_regs_data_and_2569_enex5;
  wire act_regs_data_and_2570_enex5;
  wire act_regs_data_and_2571_enex5;
  wire act_regs_data_and_2572_enex5;
  wire act_regs_data_and_2573_enex5;
  wire act_regs_data_and_2574_enex5;
  wire act_regs_data_and_2575_enex5;
  wire act_regs_data_and_2576_enex5;
  wire act_regs_data_and_2577_enex5;
  wire act_regs_data_and_2578_enex5;
  wire act_regs_data_and_2579_enex5;
  wire act_regs_data_and_2580_enex5;
  wire act_regs_data_and_2581_enex5;
  wire act_regs_data_and_2582_enex5;
  wire act_regs_data_and_2583_enex5;
  wire act_regs_data_and_2584_enex5;
  wire act_regs_data_and_2585_enex5;
  wire act_regs_data_and_2586_enex5;
  wire act_regs_data_and_2587_enex5;
  wire act_regs_data_and_2588_enex5;
  wire act_regs_data_and_2589_enex5;
  wire act_regs_data_and_2590_enex5;
  wire act_regs_data_and_2591_enex5;
  wire act_regs_data_and_2592_enex5;
  wire act_regs_data_and_2593_enex5;
  wire act_regs_data_and_2594_enex5;
  wire act_regs_data_and_2595_enex5;
  wire act_regs_data_and_2596_enex5;
  wire act_regs_data_and_2597_enex5;
  wire act_regs_data_and_2598_enex5;
  wire act_regs_data_and_2599_enex5;
  wire act_regs_data_and_2600_enex5;
  wire act_regs_data_and_2601_enex5;
  wire act_regs_data_and_2602_enex5;
  wire act_regs_data_and_2603_enex5;
  wire act_regs_data_and_2604_enex5;
  wire act_regs_data_and_2605_enex5;
  wire act_regs_data_and_2606_enex5;
  wire act_regs_data_and_2607_enex5;
  wire act_regs_data_and_2608_enex5;
  wire act_regs_data_and_2609_enex5;
  wire act_regs_data_and_2610_enex5;
  wire act_regs_data_and_2611_enex5;
  wire act_regs_data_and_2612_enex5;
  wire act_regs_data_and_2613_enex5;
  wire act_regs_data_and_2614_enex5;
  wire act_regs_data_and_2615_enex5;
  wire act_regs_data_and_2616_enex5;
  wire act_regs_data_and_2617_enex5;
  wire act_regs_data_and_2618_enex5;
  wire act_regs_data_and_2619_enex5;
  wire act_regs_data_and_2620_enex5;
  wire act_regs_data_and_2621_enex5;
  wire act_regs_data_and_2622_enex5;
  wire act_regs_data_and_2623_enex5;
  wire act_regs_data_and_2624_enex5;
  wire act_regs_data_and_2625_enex5;
  wire act_regs_data_and_2626_enex5;
  wire act_regs_data_and_2627_enex5;
  wire act_regs_data_and_2628_enex5;
  wire act_regs_data_and_2629_enex5;
  wire act_regs_data_and_2630_enex5;
  wire act_regs_data_and_2631_enex5;
  wire act_regs_data_and_2632_enex5;
  wire act_regs_data_and_2633_enex5;
  wire act_regs_data_and_2634_enex5;
  wire act_regs_data_and_2635_enex5;
  wire act_regs_data_and_2636_enex5;
  wire act_regs_data_and_2637_enex5;
  wire act_regs_data_and_2638_enex5;
  wire act_regs_data_and_2639_enex5;
  wire act_regs_data_and_2640_enex5;
  wire act_regs_data_and_2641_enex5;
  wire act_regs_data_and_2642_enex5;
  wire act_regs_data_and_2643_enex5;
  wire act_regs_data_and_2644_enex5;
  wire act_regs_data_and_2645_enex5;
  wire act_regs_data_and_2646_enex5;
  wire act_regs_data_and_2647_enex5;
  wire act_regs_data_and_2648_enex5;
  wire act_regs_data_and_2649_enex5;
  wire act_regs_data_and_2650_enex5;
  wire act_regs_data_and_2651_enex5;
  wire act_regs_data_and_2652_enex5;
  wire act_regs_data_and_2653_enex5;
  wire act_regs_data_and_2654_enex5;
  wire act_regs_data_and_2655_enex5;
  wire act_regs_data_and_2656_enex5;
  wire act_regs_data_and_2657_enex5;
  wire act_regs_data_and_2658_enex5;
  wire act_regs_data_and_2659_enex5;
  wire act_regs_data_and_2660_enex5;
  wire act_regs_data_and_2661_enex5;
  wire act_regs_data_and_2662_enex5;
  wire act_regs_data_and_2663_enex5;
  wire act_regs_data_and_2664_enex5;
  wire act_regs_data_and_2665_enex5;
  wire act_regs_data_and_2666_enex5;
  wire act_regs_data_and_2667_enex5;
  wire act_regs_data_and_2668_enex5;
  wire act_regs_data_and_2669_enex5;
  wire act_regs_data_and_2670_enex5;
  wire act_regs_data_and_2671_enex5;
  wire act_regs_data_and_2672_enex5;
  wire act_regs_data_and_2673_enex5;
  wire act_regs_data_and_2674_enex5;
  wire act_regs_data_and_2675_enex5;
  wire act_regs_data_and_2676_enex5;
  wire act_regs_data_and_2677_enex5;
  wire act_regs_data_and_2678_enex5;
  wire act_regs_data_and_2679_enex5;
  wire act_regs_data_and_2680_enex5;
  wire act_regs_data_and_2681_enex5;
  wire act_regs_data_and_2682_enex5;
  wire act_regs_data_and_2683_enex5;
  wire act_regs_data_and_2684_enex5;
  wire act_regs_data_and_2685_enex5;
  wire act_regs_data_and_2686_enex5;
  wire act_regs_data_and_2687_enex5;
  wire act_regs_data_and_2688_enex5;
  wire act_regs_data_and_2689_enex5;
  wire act_regs_data_and_2690_enex5;
  wire act_regs_data_and_2691_enex5;
  wire act_regs_data_and_2692_enex5;
  wire act_regs_data_and_2693_enex5;
  wire act_regs_data_and_2694_enex5;
  wire act_regs_data_and_2695_enex5;
  wire act_regs_data_and_2696_enex5;
  wire act_regs_data_and_2697_enex5;
  wire act_regs_data_and_2698_enex5;
  wire act_regs_data_and_2699_enex5;
  wire act_regs_data_and_2700_enex5;
  wire act_regs_data_and_2701_enex5;
  wire act_regs_data_and_2702_enex5;
  wire act_regs_data_and_2703_enex5;
  wire act_mem_banks_read_read_data_and_16_enex5;
  wire act_mem_banks_read_read_data_and_17_enex5;
  wire act_mem_banks_read_read_data_and_18_enex5;
  wire act_mem_banks_read_read_data_and_19_enex5;
  wire act_mem_banks_read_read_data_and_20_enex5;
  wire act_mem_banks_read_read_data_and_21_enex5;
  wire act_mem_banks_read_read_data_and_22_enex5;
  wire act_mem_banks_read_read_data_and_23_enex5;
  wire act_mem_banks_read_read_data_and_24_enex5;
  wire act_mem_banks_read_read_data_and_25_enex5;
  wire act_mem_banks_read_read_data_and_26_enex5;
  wire act_mem_banks_read_read_data_and_27_enex5;
  wire act_mem_banks_read_read_data_and_28_enex5;
  wire act_mem_banks_read_read_data_and_29_enex5;
  wire act_mem_banks_read_read_data_and_30_enex5;
  wire act_mem_banks_read_read_data_and_31_enex5;
  wire act_port_read_out_data_and_16_enex5;
  wire act_port_read_out_data_and_17_enex5;
  wire act_port_read_out_data_and_18_enex5;
  wire act_port_read_out_data_and_19_enex5;
  wire act_port_read_out_data_and_20_enex5;
  wire act_port_read_out_data_and_21_enex5;
  wire act_port_read_out_data_and_22_enex5;
  wire act_port_read_out_data_and_23_enex5;
  wire act_port_read_out_data_and_24_enex5;
  wire act_port_read_out_data_and_25_enex5;
  wire act_port_read_out_data_and_26_enex5;
  wire act_port_read_out_data_and_27_enex5;
  wire act_port_read_out_data_and_28_enex5;
  wire act_port_read_out_data_and_29_enex5;
  wire act_port_read_out_data_and_30_enex5;
  wire act_port_read_out_data_and_31_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_37_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_38_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_39_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_40_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_41_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_42_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_43_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_44_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_45_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_46_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_47_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_48_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_49_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_50_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_51_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_52_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_53_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_54_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_55_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_56_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_57_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_58_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_59_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_60_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_61_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_62_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_63_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_64_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_65_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_66_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_67_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_68_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_69_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_70_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_71_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_72_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_73_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_74_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_75_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_76_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_77_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_78_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_79_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_80_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_81_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_82_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_83_enex5;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_84_enex5;
  wire Tanh_for_y_and_31_enex5;
  wire Tanh_for_y_and_32_enex5;
  wire Tanh_for_y_and_33_enex5;
  wire Tanh_for_y_and_34_enex5;
  wire Tanh_for_y_and_35_enex5;
  wire Tanh_for_y_and_36_enex5;
  wire Tanh_for_y_and_37_enex5;
  wire Tanh_for_y_and_38_enex5;
  wire Tanh_for_y_and_39_enex5;
  wire Tanh_for_y_and_40_enex5;
  wire Tanh_for_y_and_41_enex5;
  wire Tanh_for_y_and_42_enex5;
  wire Tanh_for_y_and_43_enex5;
  wire Tanh_for_y_and_44_enex5;
  wire Tanh_for_y_and_45_enex5;
  wire Tanh_for_y_and_46_enex5;
  wire Tanh_for_y_and_47_enex5;
  wire Tanh_for_y_and_48_enex5;
  wire Tanh_for_y_and_49_enex5;
  wire Tanh_for_y_and_50_enex5;
  wire Tanh_for_y_and_51_enex5;
  wire Tanh_for_y_and_52_enex5;
  wire Tanh_for_y_and_53_enex5;
  wire Tanh_for_y_and_54_enex5;
  wire Tanh_for_y_and_55_enex5;
  wire Tanh_for_y_and_56_enex5;
  wire Tanh_for_y_and_57_enex5;
  wire Tanh_for_y_and_58_enex5;
  wire Tanh_for_y_and_59_enex5;
  wire Tanh_for_y_and_60_enex5;
  wire Tanh_for_y_and_61_enex5;
  wire Tanh_for_y_and_62_enex5;
  wire Relu_for_y_qelse_and_31_enex5;
  wire Relu_for_y_qelse_and_32_enex5;
  wire Relu_for_y_qelse_and_33_enex5;
  wire Relu_for_y_qelse_and_34_enex5;
  wire Relu_for_y_qelse_and_35_enex5;
  wire Relu_for_y_qelse_and_36_enex5;
  wire Relu_for_y_qelse_and_37_enex5;
  wire Relu_for_y_qelse_and_38_enex5;
  wire Relu_for_y_qelse_and_39_enex5;
  wire Relu_for_y_qelse_and_40_enex5;
  wire Relu_for_y_qelse_and_41_enex5;
  wire Relu_for_y_qelse_and_42_enex5;
  wire Relu_for_y_qelse_and_43_enex5;
  wire Relu_for_y_qelse_and_44_enex5;
  wire Relu_for_y_qelse_and_45_enex5;
  wire Relu_for_y_qelse_and_46_enex5;
  wire Relu_for_y_qelse_and_47_enex5;
  wire Relu_for_y_qelse_and_48_enex5;
  wire Relu_for_y_qelse_and_49_enex5;
  wire Relu_for_y_qelse_and_50_enex5;
  wire Relu_for_y_qelse_and_51_enex5;
  wire Relu_for_y_qelse_and_52_enex5;
  wire Relu_for_y_qelse_and_53_enex5;
  wire Relu_for_y_qelse_and_54_enex5;
  wire Relu_for_y_qelse_and_55_enex5;
  wire Relu_for_y_qelse_and_56_enex5;
  wire Relu_for_y_qelse_and_57_enex5;
  wire Relu_for_y_qelse_and_58_enex5;
  wire Relu_for_y_qelse_and_59_enex5;
  wire Relu_for_y_qelse_and_60_enex5;
  wire Relu_for_y_qelse_and_61_enex5;
  wire Relu_for_y_qelse_and_62_enex5;
  wire Relu_for_y_qelse_and_63_enex5;
  wire Relu_for_y_qelse_and_64_enex5;
  wire Relu_for_y_qelse_and_65_enex5;
  wire Relu_for_y_qelse_and_66_enex5;
  wire Relu_for_y_qelse_and_67_enex5;
  wire Relu_for_y_qelse_and_68_enex5;
  wire Relu_for_y_qelse_and_69_enex5;
  wire Relu_for_y_qelse_and_70_enex5;
  wire Relu_for_y_qelse_and_71_enex5;
  wire Relu_for_y_qelse_and_72_enex5;
  wire Relu_for_y_qelse_and_73_enex5;
  wire Relu_for_y_qelse_and_74_enex5;
  wire Relu_for_y_qelse_and_75_enex5;
  wire Relu_for_y_qelse_and_76_enex5;
  wire Relu_for_y_qelse_and_77_enex5;
  wire Relu_for_y_qelse_and_78_enex5;
  wire ActUnit_RunInst_curr_inst_and_enex5;
  wire ActUnit_RunInst_switch_lp_and_813_enex5;
  wire ActUnit_RunInst_switch_lp_and_814_enex5;
  wire ActUnit_RunInst_switch_lp_and_815_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_15_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_16_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_17_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_18_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_19_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_20_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_21_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_22_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_23_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_24_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_25_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_26_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_27_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_28_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_29_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_30_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_31_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_32_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_33_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_34_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_35_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_36_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_37_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_38_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_39_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_40_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_41_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_42_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_43_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_44_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_45_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_46_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_47_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_48_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_49_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_50_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_51_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_52_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_53_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_54_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_55_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_56_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_57_enex5;
  wire nv_scvector_cctor_nv_scvector_6_for_and_58_enex5;
  wire act_regs_data_and_2704_enex5;
  wire act_regs_data_and_2705_enex5;
  wire act_regs_data_and_2706_enex5;
  wire act_regs_data_and_2707_enex5;
  wire act_regs_data_and_2708_enex5;
  wire act_regs_data_and_2709_enex5;
  wire act_regs_data_and_2710_enex5;
  wire act_regs_data_and_2711_enex5;
  wire act_regs_data_and_2712_enex5;
  wire act_regs_data_and_2713_enex5;
  wire act_regs_data_and_2714_enex5;
  wire act_regs_data_and_2715_enex5;
  wire act_regs_data_and_2716_enex5;
  wire act_regs_data_and_2717_enex5;
  wire act_regs_data_and_2718_enex5;
  wire act_regs_data_and_2719_enex5;
  wire act_regs_data_and_2720_enex5;
  wire act_regs_data_and_2721_enex5;
  wire act_regs_data_and_2722_enex5;
  wire act_regs_data_and_2723_enex5;
  wire act_regs_data_and_2724_enex5;
  wire act_regs_data_and_2725_enex5;
  wire act_regs_data_and_2726_enex5;
  wire act_regs_data_and_2727_enex5;
  wire act_regs_data_and_2728_enex5;
  wire act_regs_data_and_2729_enex5;
  wire act_regs_data_and_2730_enex5;
  wire act_regs_data_and_2731_enex5;
  wire act_regs_data_and_2732_enex5;
  wire act_regs_data_and_2733_enex5;
  wire act_regs_data_and_2734_enex5;
  wire act_regs_data_and_2735_enex5;
  wire act_regs_data_and_2736_enex5;
  wire act_regs_data_and_2737_enex5;
  wire act_regs_data_and_2738_enex5;
  wire act_regs_data_and_2739_enex5;
  wire act_regs_data_and_2740_enex5;
  wire act_regs_data_and_2741_enex5;
  wire act_regs_data_and_2742_enex5;
  wire act_regs_data_and_2743_enex5;
  wire act_regs_data_and_2744_enex5;
  wire act_regs_data_and_2745_enex5;
  wire act_regs_data_and_2746_enex5;
  wire act_regs_data_and_2747_enex5;
  wire act_regs_data_and_2748_enex5;
  wire act_regs_data_and_2749_enex5;
  wire act_regs_data_and_2750_enex5;
  wire act_regs_data_and_2751_enex5;
  wire act_regs_data_and_2752_enex5;
  wire act_regs_data_and_2753_enex5;
  wire act_regs_data_and_2754_enex5;
  wire act_regs_data_and_2755_enex5;
  wire act_regs_data_and_2756_enex5;
  wire act_regs_data_and_2757_enex5;
  wire act_regs_data_and_2758_enex5;
  wire act_regs_data_and_2759_enex5;
  wire act_regs_data_and_2760_enex5;
  wire act_regs_data_and_2761_enex5;
  wire act_regs_data_and_2762_enex5;
  wire act_regs_data_and_2763_enex5;
  wire act_regs_data_and_2764_enex5;
  wire act_regs_data_and_2765_enex5;
  wire act_regs_data_and_2766_enex5;
  wire ActUnit_RunInst_switch_lp_and_816_enex5;
  wire ActUnit_RunInst_switch_lp_and_817_enex5;
  wire ActUnit_RunInst_switch_lp_and_818_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_15_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_16_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_17_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_18_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_19_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_20_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_21_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_22_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_23_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_24_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_25_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_26_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_27_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_28_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_29_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_30_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_31_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_32_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_33_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_34_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_35_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_36_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_37_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_38_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_39_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_40_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_41_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_42_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_43_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_44_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_45_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_46_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_47_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_48_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_49_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_50_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_51_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_52_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_53_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_54_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_55_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_56_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_57_enex5;
  wire nv_scvector_cctor_nv_scvector_5_for_and_58_enex5;
  wire is_start_and_tmp;
  wire and_2189_tmp;
  wire w_load_and_tmp;
  wire and_2187_tmp;
  wire and_2185_tmp;
  wire and_2183_tmp;
  wire and_2181_tmp;
  wire and_2179_tmp;
  wire and_2177_tmp;
  wire and_2175_tmp;
  wire and_2173_tmp;
  wire and_2171_tmp;
  wire and_2169_tmp;
  wire and_2167_tmp;
  wire and_2165_tmp;
  wire and_2163_tmp;
  wire and_2161_tmp;
  wire and_2159_tmp;
  wire and_2157_tmp;
  wire and_2155_tmp;
  wire and_2153_tmp;
  wire and_2151_tmp;
  wire and_2149_tmp;
  wire and_2147_tmp;
  wire and_2145_tmp;
  wire and_2143_tmp;
  wire and_2141_tmp;
  wire and_2139_tmp;
  wire and_2137_tmp;
  wire and_2135_tmp;
  wire and_2133_tmp;
  wire and_2131_tmp;
  wire and_2129_tmp;
  wire and_2127_tmp;
  wire and_2125_tmp;
  wire and_2123_tmp;
  wire and_2121_tmp;
  wire and_2119_tmp;
  wire and_2117_tmp;
  wire and_2115_tmp;
  wire and_2113_tmp;
  wire and_2111_tmp;
  wire and_2109_tmp;
  wire and_2107_tmp;
  wire and_2105_tmp;
  wire and_2103_tmp;
  wire and_2101_tmp;
  wire and_2099_tmp;
  wire and_2097_tmp;
  wire and_2095_tmp;
  wire and_2093_tmp;
  wire and_1891_tmp;
  wire and_1867_tmp;
  wire and_1933_tmp;
  wire and_2091_tmp;
  wire and_1889_tmp;
  wire and_1865_tmp;
  wire and_2081_tmp;
  wire and_2079_tmp;
  wire and_1877_tmp;
  wire and_2077_tmp;
  wire and_1903_tmp;
  wire and_1864_tmp;
  wire and_2075_tmp;
  wire and_1901_tmp;
  wire and_1879_tmp;
  wire and_2073_tmp;
  wire and_1899_tmp;
  wire and_1875_tmp;
  wire and_2071_tmp;
  wire and_1897_tmp;
  wire and_1873_tmp;
  wire and_2069_tmp;
  wire and_1895_tmp;
  wire and_1871_tmp;
  wire and_2067_tmp;
  wire and_1893_tmp;
  wire and_1869_tmp;
  wire act_config_inst_counter_and_tmp;
  wire ActUnit_PushOutput_if_for_i_and_tmp;
  wire ActUnit_RunLoad_if_a2_and_tmp;
  wire and_1927_tmp;
  wire and_2089_tmp;
  wire and_1887_tmp;
  wire and_2328_tmp;
  wire and_1921_tmp;
  wire and_2087_tmp;
  wire and_1885_tmp;
  wire and_2327_tmp;
  wire and_1915_tmp;
  wire and_2085_tmp;
  wire and_1883_tmp;
  wire and_2326_tmp;
  wire and_1909_tmp;
  wire and_2083_tmp;
  wire and_1881_tmp;
  wire and_2325_tmp;
  wire and_1803_tmp;
  wire and_2065_tmp;
  wire and_1801_tmp;
  wire and_2324_tmp;
  wire and_1808_tmp;
  wire and_2063_tmp;
  wire rva_out_reg_data_and_61_tmp;
  wire Silu_for_else_else_else_if_and_tmp;
  wire or_243_cse;
  wire Silu_for_else_if_Silu_for_else_if_or_itm;
  wire Silu_for_else_or_7_itm;
  wire Silu_for_else_or_6_itm;
  wire Silu_for_else_or_5_itm;
  wire Silu_for_else_or_4_itm;
  wire Silu_for_else_or_3_itm;
  wire Silu_for_else_or_2_itm;
  wire Silu_for_else_or_1_itm;
  wire Silu_for_else_or_itm;
  wire Silu_for_else_or_15_itm;
  wire Silu_for_else_or_14_itm;
  wire Silu_for_else_or_13_itm;
  wire Silu_for_else_or_12_itm;
  wire Silu_for_else_or_11_itm;
  wire Silu_for_else_or_10_itm;
  wire Silu_for_else_or_9_itm;
  wire Silu_for_else_or_8_itm;
  wire [24:0] Silu_for_1_else_else_else_if_acc_itm_25_1_1;
  wire [24:0] Silu_for_2_else_else_else_if_acc_itm_25_1_1;
  wire [24:0] Silu_for_3_else_else_else_if_acc_itm_25_1_1;
  wire [24:0] Silu_for_4_else_else_else_if_acc_itm_25_1_1;
  wire [24:0] Silu_for_5_else_else_else_if_acc_itm_25_1_1;
  wire [24:0] Silu_for_6_else_else_else_if_acc_itm_25_1_1;
  wire [24:0] Silu_for_7_else_else_else_if_acc_itm_25_1_1;
  wire [24:0] Silu_for_8_else_else_else_if_acc_itm_25_1_1;
  wire [24:0] Silu_for_9_else_else_else_if_acc_itm_25_1_1;
  wire [24:0] Silu_for_10_else_else_else_if_acc_itm_25_1_1;
  wire [24:0] Silu_for_11_else_else_else_if_acc_itm_25_1_1;
  wire [24:0] Silu_for_12_else_else_else_if_acc_itm_25_1_1;
  wire [24:0] Silu_for_13_else_else_else_if_acc_itm_25_1_1;
  wire [24:0] Silu_for_14_else_else_else_if_acc_itm_25_1_1;
  wire [24:0] Silu_for_15_else_else_else_if_acc_itm_25_1_1;
  wire [24:0] Silu_for_16_else_else_else_if_acc_itm_25_1_1;
  reg act_regs_data_0_0_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_0_0_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_0_1_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_0_1_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_0_2_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_0_2_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_0_3_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_0_3_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_0_4_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_0_4_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_0_5_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_0_5_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_0_6_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_0_6_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_0_7_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_0_7_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_0_8_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_0_8_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_0_9_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_0_9_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_0_10_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_0_10_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_0_11_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_0_11_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_0_12_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_0_12_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_0_13_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_0_13_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_0_14_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_0_14_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_0_15_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_0_15_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_1_0_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_1_0_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_1_1_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_1_1_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_1_2_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_1_2_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_1_3_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_1_3_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_1_4_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_1_4_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_1_5_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_1_5_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_1_6_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_1_6_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_1_7_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_1_7_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_1_8_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_1_8_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_1_9_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_1_9_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_1_10_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_1_10_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_1_11_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_1_11_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_1_12_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_1_12_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_1_13_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_1_13_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_1_14_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_1_14_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_1_15_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_1_15_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_2_0_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_2_0_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_2_1_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_2_1_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_2_2_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_2_2_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_2_3_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_2_3_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_2_4_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_2_4_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_2_5_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_2_5_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_2_6_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_2_6_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_2_7_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_2_7_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_2_8_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_2_8_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_2_9_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_2_9_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_2_10_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_2_10_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_2_11_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_2_11_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_2_12_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_2_12_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_2_13_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_2_13_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_2_14_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_2_14_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_2_15_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_2_15_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_3_0_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_3_0_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_3_1_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_3_1_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_3_2_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_3_2_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_3_3_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_3_3_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_3_4_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_3_4_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_3_5_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_3_5_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_3_6_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_3_6_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_3_7_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_3_7_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_3_8_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_3_8_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_3_9_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_3_9_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_3_10_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_3_10_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_3_11_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_3_11_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_3_12_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_3_12_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_3_13_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_3_13_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_3_14_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_3_14_sva_dfm_2_25_22_rsp_1;
  reg act_regs_data_3_15_sva_dfm_2_25_22_rsp_0;
  reg [2:0] act_regs_data_3_15_sva_dfm_2_25_22_rsp_1;
  reg reg_act_regs_data_0_13_ftd_2_3;
  reg [2:0] reg_act_regs_data_0_13_ftd_2_2_0;
  reg reg_act_regs_data_0_12_ftd_2_3;
  reg [2:0] reg_act_regs_data_0_12_ftd_2_2_0;
  reg reg_act_regs_data_0_11_ftd_2_3;
  reg [2:0] reg_act_regs_data_0_11_ftd_2_2_0;
  reg reg_act_regs_data_0_10_ftd_2_3;
  reg [2:0] reg_act_regs_data_0_10_ftd_2_2_0;
  reg reg_act_regs_data_0_1_ftd_2_3;
  reg [2:0] reg_act_regs_data_0_1_ftd_2_2_0;
  reg reg_act_regs_data_0_0_ftd_2_3;
  reg [2:0] reg_act_regs_data_0_0_ftd_2_2_0;
  wire [3:0] Silu_for_2_else_else_else_else_if_acc_sdt;
  wire [4:0] nl_Silu_for_2_else_else_else_else_if_acc_sdt;
  reg ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_1_25;
  reg [2:0] ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_1_24_22;
  wire [3:0] Silu_for_1_else_else_else_else_if_acc_sdt;
  wire [4:0] nl_Silu_for_1_else_else_else_else_if_acc_sdt;
  reg ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_1_25;
  reg [2:0] ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_1_24_22;
  wire [3:0] Silu_for_16_else_else_else_else_if_acc_sdt;
  wire [4:0] nl_Silu_for_16_else_else_else_else_if_acc_sdt;
  reg ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_1_25;
  reg [2:0] ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_1_24_22;
  wire [3:0] Silu_for_15_else_else_else_else_if_acc_sdt;
  wire [4:0] nl_Silu_for_15_else_else_else_else_if_acc_sdt;
  reg ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_1_25;
  reg [2:0] ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_1_24_22;
  wire [3:0] Silu_for_14_else_else_else_else_if_acc_sdt;
  wire [4:0] nl_Silu_for_14_else_else_else_else_if_acc_sdt;
  reg ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_1_25;
  reg [2:0] ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_1_24_22;
  reg ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_1_25;
  reg [2:0] ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_1_24_22;
  wire [3:0] Silu_for_9_else_else_else_else_if_acc_sdt;
  wire [4:0] nl_Silu_for_9_else_else_else_else_if_acc_sdt;
  reg ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_1_25;
  reg [2:0] ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_1_24_22;
  wire [3:0] Silu_for_8_else_else_else_else_if_acc_sdt;
  wire [4:0] nl_Silu_for_8_else_else_else_else_if_acc_sdt;
  reg ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_1_25;
  reg [2:0] ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_1_24_22;
  wire [3:0] Silu_for_7_else_else_else_else_if_acc_sdt;
  wire [4:0] nl_Silu_for_7_else_else_else_else_if_acc_sdt;
  reg ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_1_25;
  reg [2:0] ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_1_24_22;
  wire [3:0] Silu_for_6_else_else_else_else_if_acc_sdt;
  wire [4:0] nl_Silu_for_6_else_else_else_else_if_acc_sdt;
  reg ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_1_25;
  reg [2:0] ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_1_24_22;
  wire [3:0] Silu_for_5_else_else_else_else_if_acc_sdt;
  wire [4:0] nl_Silu_for_5_else_else_else_else_if_acc_sdt;
  reg ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_1_25;
  reg [2:0] ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_1_24_22;
  wire [3:0] Silu_for_4_else_else_else_else_if_acc_sdt;
  wire [4:0] nl_Silu_for_4_else_else_else_else_if_acc_sdt;
  reg ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_1_25;
  reg [2:0] ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_1_24_22;
  wire [3:0] Silu_for_3_else_else_else_else_if_acc_sdt;
  wire [4:0] nl_Silu_for_3_else_else_else_else_if_acc_sdt;
  reg ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_1_25;
  reg [2:0] ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_1_24_22;
  wire [3:0] Silu_for_13_else_else_else_else_if_acc_sdt;
  wire [4:0] nl_Silu_for_13_else_else_else_else_if_acc_sdt;
  wire and_1715_ssc;
  reg rva_out_reg_data_39_32_sva_dfm_6_3;
  reg [2:0] rva_out_reg_data_39_32_sva_dfm_6_2_0;
  wire [3:0] Silu_for_12_else_else_else_else_if_acc_sdt;
  wire [4:0] nl_Silu_for_12_else_else_else_else_if_acc_sdt;
  reg rva_out_reg_data_29_24_sva_dfm_6_3;
  reg [2:0] rva_out_reg_data_29_24_sva_dfm_6_2_0;
  reg Silu_for_y_1_lpi_1_dfm_4_25;
  reg [2:0] Silu_for_y_1_lpi_1_dfm_4_24_22;
  reg Silu_for_y_2_lpi_1_dfm_4_25;
  reg [2:0] Silu_for_y_2_lpi_1_dfm_4_24_22;
  reg Silu_for_y_3_lpi_1_dfm_4_25;
  reg [2:0] Silu_for_y_3_lpi_1_dfm_4_24_22;
  reg Silu_for_y_4_lpi_1_dfm_4_25;
  reg [2:0] Silu_for_y_4_lpi_1_dfm_4_24_22;
  reg Silu_for_y_5_lpi_1_dfm_4_25;
  reg [2:0] Silu_for_y_5_lpi_1_dfm_4_24_22;
  reg Silu_for_y_6_lpi_1_dfm_4_25;
  reg [2:0] Silu_for_y_6_lpi_1_dfm_4_24_22;
  reg Silu_for_y_7_lpi_1_dfm_4_25;
  reg [2:0] Silu_for_y_7_lpi_1_dfm_4_24_22;
  reg Silu_for_y_8_lpi_1_dfm_4_25;
  reg [2:0] Silu_for_y_8_lpi_1_dfm_4_24_22;
  reg act_regs_data_1_15_sva_8_25;
  reg [2:0] act_regs_data_1_15_sva_8_24_22;
  reg act_regs_data_2_0_sva_8_25;
  reg [2:0] act_regs_data_2_0_sva_8_24_22;
  reg act_regs_data_1_14_sva_8_25;
  reg [2:0] act_regs_data_1_14_sva_8_24_22;
  reg act_regs_data_2_1_sva_8_25;
  reg [2:0] act_regs_data_2_1_sva_8_24_22;
  reg act_regs_data_1_13_sva_8_25;
  reg [2:0] act_regs_data_1_13_sva_8_24_22;
  reg act_regs_data_2_2_sva_8_25;
  reg [2:0] act_regs_data_2_2_sva_8_24_22;
  reg act_regs_data_1_12_sva_8_25;
  reg [2:0] act_regs_data_1_12_sva_8_24_22;
  reg act_regs_data_2_3_sva_8_25;
  reg [2:0] act_regs_data_2_3_sva_8_24_22;
  reg act_regs_data_1_11_sva_8_25;
  reg [2:0] act_regs_data_1_11_sva_8_24_22;
  reg act_regs_data_2_4_sva_8_25;
  reg [2:0] act_regs_data_2_4_sva_8_24_22;
  reg act_regs_data_1_10_sva_8_25;
  reg [2:0] act_regs_data_1_10_sva_8_24_22;
  reg act_regs_data_2_5_sva_8_25;
  reg [2:0] act_regs_data_2_5_sva_8_24_22;
  reg act_regs_data_1_9_sva_8_25;
  reg [2:0] act_regs_data_1_9_sva_8_24_22;
  reg act_regs_data_2_6_sva_8_25;
  reg [2:0] act_regs_data_2_6_sva_8_24_22;
  reg act_regs_data_1_8_sva_8_25;
  reg [2:0] act_regs_data_1_8_sva_8_24_22;
  reg act_regs_data_2_7_sva_8_25;
  reg [2:0] act_regs_data_2_7_sva_8_24_22;
  reg act_regs_data_1_7_sva_8_25;
  reg [2:0] act_regs_data_1_7_sva_8_24_22;
  reg act_regs_data_2_8_sva_8_25;
  reg [2:0] act_regs_data_2_8_sva_8_24_22;
  reg act_regs_data_1_6_sva_8_25;
  reg [2:0] act_regs_data_1_6_sva_8_24_22;
  reg act_regs_data_2_9_sva_8_25;
  reg [2:0] act_regs_data_2_9_sva_8_24_22;
  reg act_regs_data_1_5_sva_8_25;
  reg [2:0] act_regs_data_1_5_sva_8_24_22;
  reg act_regs_data_2_10_sva_8_25;
  reg [2:0] act_regs_data_2_10_sva_8_24_22;
  reg act_regs_data_1_4_sva_8_25;
  reg [2:0] act_regs_data_1_4_sva_8_24_22;
  reg act_regs_data_2_11_sva_8_25;
  reg [2:0] act_regs_data_2_11_sva_8_24_22;
  reg act_regs_data_1_3_sva_8_25;
  reg [2:0] act_regs_data_1_3_sva_8_24_22;
  reg act_regs_data_2_12_sva_8_25;
  reg [2:0] act_regs_data_2_12_sva_8_24_22;
  reg act_regs_data_1_2_sva_8_25;
  reg [2:0] act_regs_data_1_2_sva_8_24_22;
  reg act_regs_data_2_13_sva_8_25;
  reg [2:0] act_regs_data_2_13_sva_8_24_22;
  reg act_regs_data_1_1_sva_8_25;
  reg [2:0] act_regs_data_1_1_sva_8_24_22;
  reg act_regs_data_2_14_sva_8_25;
  reg [2:0] act_regs_data_2_14_sva_8_24_22;
  reg act_regs_data_1_0_sva_8_25;
  reg [2:0] act_regs_data_1_0_sva_8_24_22;
  reg act_regs_data_2_15_sva_8_25;
  reg [2:0] act_regs_data_2_15_sva_8_24_22;
  reg act_regs_data_0_15_sva_8_25;
  reg [2:0] act_regs_data_0_15_sva_8_24_22;
  reg act_regs_data_3_0_sva_8_25;
  reg [2:0] act_regs_data_3_0_sva_8_24_22;
  reg act_regs_data_0_14_sva_8_25;
  reg [2:0] act_regs_data_0_14_sva_8_24_22;
  reg act_regs_data_3_1_sva_8_25;
  reg [2:0] act_regs_data_3_1_sva_8_24_22;
  reg act_regs_data_0_13_sva_8_25;
  reg [2:0] act_regs_data_0_13_sva_8_24_22;
  reg act_regs_data_3_2_sva_8_25;
  reg [2:0] act_regs_data_3_2_sva_8_24_22;
  reg act_regs_data_0_12_sva_8_25;
  reg [2:0] act_regs_data_0_12_sva_8_24_22;
  reg act_regs_data_3_3_sva_8_25;
  reg [2:0] act_regs_data_3_3_sva_8_24_22;
  reg act_regs_data_0_11_sva_8_25;
  reg [2:0] act_regs_data_0_11_sva_8_24_22;
  reg act_regs_data_3_4_sva_8_25;
  reg [2:0] act_regs_data_3_4_sva_8_24_22;
  reg act_regs_data_0_10_sva_8_25;
  reg [2:0] act_regs_data_0_10_sva_8_24_22;
  reg act_regs_data_3_5_sva_8_25;
  reg [2:0] act_regs_data_3_5_sva_8_24_22;
  reg act_regs_data_0_9_sva_8_25;
  reg [2:0] act_regs_data_0_9_sva_8_24_22;
  reg act_regs_data_3_6_sva_8_25;
  reg [2:0] act_regs_data_3_6_sva_8_24_22;
  reg act_regs_data_0_8_sva_8_25;
  reg [2:0] act_regs_data_0_8_sva_8_24_22;
  reg act_regs_data_3_7_sva_8_25;
  reg [2:0] act_regs_data_3_7_sva_8_24_22;
  reg act_regs_data_0_7_sva_8_25;
  reg [2:0] act_regs_data_0_7_sva_8_24_22;
  reg act_regs_data_3_8_sva_8_25;
  reg [2:0] act_regs_data_3_8_sva_8_24_22;
  reg act_regs_data_0_6_sva_8_25;
  reg [2:0] act_regs_data_0_6_sva_8_24_22;
  reg act_regs_data_3_9_sva_8_25;
  reg [2:0] act_regs_data_3_9_sva_8_24_22;
  reg act_regs_data_0_5_sva_8_25;
  reg [2:0] act_regs_data_0_5_sva_8_24_22;
  reg act_regs_data_3_10_sva_8_25;
  reg [2:0] act_regs_data_3_10_sva_8_24_22;
  reg act_regs_data_0_4_sva_8_25;
  reg [2:0] act_regs_data_0_4_sva_8_24_22;
  reg act_regs_data_3_11_sva_8_25;
  reg [2:0] act_regs_data_3_11_sva_8_24_22;
  reg act_regs_data_0_3_sva_8_25;
  reg [2:0] act_regs_data_0_3_sva_8_24_22;
  reg act_regs_data_3_12_sva_8_25;
  reg [2:0] act_regs_data_3_12_sva_8_24_22;
  reg act_regs_data_0_2_sva_8_25;
  reg [2:0] act_regs_data_0_2_sva_8_24_22;
  reg act_regs_data_3_13_sva_8_25;
  reg [2:0] act_regs_data_3_13_sva_8_24_22;
  reg act_regs_data_0_1_sva_8_25;
  reg [2:0] act_regs_data_0_1_sva_8_24_22;
  reg act_regs_data_3_14_sva_8_25;
  reg [2:0] act_regs_data_3_14_sva_8_24_22;
  reg act_regs_data_0_0_sva_8_25;
  reg [2:0] act_regs_data_0_0_sva_8_24_22;
  reg act_regs_data_3_15_sva_8_25;
  reg [2:0] act_regs_data_3_15_sva_8_24_22;
  wire Silu_for_y_lpi_1_dfm_4_25;
  wire [2:0] Silu_for_y_lpi_1_dfm_4_24_22;
  wire Silu_for_y_15_lpi_1_dfm_4_25;
  wire [2:0] Silu_for_y_15_lpi_1_dfm_4_24_22;
  wire Silu_for_y_14_lpi_1_dfm_4_25;
  wire [2:0] Silu_for_y_14_lpi_1_dfm_4_24_22;
  wire Silu_for_y_13_lpi_1_dfm_4_25;
  wire [2:0] Silu_for_y_13_lpi_1_dfm_4_24_22;
  wire Silu_for_y_12_lpi_1_dfm_4_25;
  wire [2:0] Silu_for_y_12_lpi_1_dfm_4_24_22;
  wire Silu_for_y_11_lpi_1_dfm_4_25;
  wire [2:0] Silu_for_y_11_lpi_1_dfm_4_24_22;
  wire Silu_for_y_10_lpi_1_dfm_4_25;
  wire [2:0] Silu_for_y_10_lpi_1_dfm_4_24_22;
  wire Silu_for_y_9_lpi_1_dfm_4_25;
  wire [2:0] Silu_for_y_9_lpi_1_dfm_4_24_22;
  reg act_regs_data_1_15_sva_25;
  reg [2:0] act_regs_data_1_15_sva_24_22;
  reg act_regs_data_2_0_sva_25;
  reg [2:0] act_regs_data_2_0_sva_24_22;
  reg act_regs_data_1_14_sva_25;
  reg [2:0] act_regs_data_1_14_sva_24_22;
  reg act_regs_data_2_1_sva_25;
  reg [2:0] act_regs_data_2_1_sva_24_22;
  reg act_regs_data_1_13_sva_25;
  reg [2:0] act_regs_data_1_13_sva_24_22;
  reg act_regs_data_2_2_sva_25;
  reg [2:0] act_regs_data_2_2_sva_24_22;
  reg act_regs_data_1_12_sva_25;
  reg [2:0] act_regs_data_1_12_sva_24_22;
  reg act_regs_data_2_3_sva_25;
  reg [2:0] act_regs_data_2_3_sva_24_22;
  reg act_regs_data_1_11_sva_25;
  reg [2:0] act_regs_data_1_11_sva_24_22;
  reg act_regs_data_2_4_sva_25;
  reg [2:0] act_regs_data_2_4_sva_24_22;
  reg act_regs_data_1_10_sva_25;
  reg [2:0] act_regs_data_1_10_sva_24_22;
  reg act_regs_data_2_5_sva_25;
  reg [2:0] act_regs_data_2_5_sva_24_22;
  reg act_regs_data_1_9_sva_25;
  reg [2:0] act_regs_data_1_9_sva_24_22;
  reg act_regs_data_2_6_sva_25;
  reg [2:0] act_regs_data_2_6_sva_24_22;
  reg act_regs_data_1_8_sva_25;
  reg [2:0] act_regs_data_1_8_sva_24_22;
  reg act_regs_data_2_7_sva_25;
  reg [2:0] act_regs_data_2_7_sva_24_22;
  reg act_regs_data_1_7_sva_25;
  reg [2:0] act_regs_data_1_7_sva_24_22;
  reg act_regs_data_2_8_sva_25;
  reg [2:0] act_regs_data_2_8_sva_24_22;
  reg act_regs_data_1_6_sva_25;
  reg [2:0] act_regs_data_1_6_sva_24_22;
  reg act_regs_data_2_9_sva_25;
  reg [2:0] act_regs_data_2_9_sva_24_22;
  reg act_regs_data_1_5_sva_25;
  reg [2:0] act_regs_data_1_5_sva_24_22;
  reg act_regs_data_2_10_sva_25;
  reg [2:0] act_regs_data_2_10_sva_24_22;
  reg act_regs_data_1_4_sva_25;
  reg [2:0] act_regs_data_1_4_sva_24_22;
  reg act_regs_data_2_11_sva_25;
  reg [2:0] act_regs_data_2_11_sva_24_22;
  reg act_regs_data_1_3_sva_25;
  reg [2:0] act_regs_data_1_3_sva_24_22;
  reg act_regs_data_2_12_sva_25;
  reg [2:0] act_regs_data_2_12_sva_24_22;
  reg act_regs_data_1_2_sva_25;
  reg [2:0] act_regs_data_1_2_sva_24_22;
  reg act_regs_data_2_13_sva_25;
  reg [2:0] act_regs_data_2_13_sva_24_22;
  reg act_regs_data_1_1_sva_25;
  reg [2:0] act_regs_data_1_1_sva_24_22;
  reg act_regs_data_2_14_sva_25;
  reg [2:0] act_regs_data_2_14_sva_24_22;
  reg act_regs_data_1_0_sva_25;
  reg [2:0] act_regs_data_1_0_sva_24_22;
  reg act_regs_data_2_15_sva_25;
  reg [2:0] act_regs_data_2_15_sva_24_22;
  reg act_regs_data_0_15_sva_25;
  reg [2:0] act_regs_data_0_15_sva_24_22;
  reg act_regs_data_3_0_sva_25;
  reg [2:0] act_regs_data_3_0_sva_24_22;
  reg act_regs_data_0_14_sva_25;
  reg [2:0] act_regs_data_0_14_sva_24_22;
  reg act_regs_data_3_1_sva_25;
  reg [2:0] act_regs_data_3_1_sva_24_22;
  reg act_regs_data_3_2_sva_25;
  reg [2:0] act_regs_data_3_2_sva_24_22;
  reg act_regs_data_3_3_sva_25;
  reg [2:0] act_regs_data_3_3_sva_24_22;
  reg act_regs_data_3_4_sva_25;
  reg [2:0] act_regs_data_3_4_sva_24_22;
  reg act_regs_data_3_5_sva_25;
  reg [2:0] act_regs_data_3_5_sva_24_22;
  reg act_regs_data_0_9_sva_25;
  reg [2:0] act_regs_data_0_9_sva_24_22;
  reg act_regs_data_3_6_sva_25;
  reg [2:0] act_regs_data_3_6_sva_24_22;
  reg act_regs_data_0_8_sva_25;
  reg [2:0] act_regs_data_0_8_sva_24_22;
  reg act_regs_data_3_7_sva_25;
  reg [2:0] act_regs_data_3_7_sva_24_22;
  reg act_regs_data_0_7_sva_25;
  reg [2:0] act_regs_data_0_7_sva_24_22;
  reg act_regs_data_3_8_sva_25;
  reg [2:0] act_regs_data_3_8_sva_24_22;
  reg act_regs_data_0_6_sva_25;
  reg [2:0] act_regs_data_0_6_sva_24_22;
  reg act_regs_data_3_9_sva_25;
  reg [2:0] act_regs_data_3_9_sva_24_22;
  reg act_regs_data_0_5_sva_25;
  reg [2:0] act_regs_data_0_5_sva_24_22;
  reg act_regs_data_3_10_sva_25;
  reg [2:0] act_regs_data_3_10_sva_24_22;
  reg act_regs_data_0_4_sva_25;
  reg [2:0] act_regs_data_0_4_sva_24_22;
  reg act_regs_data_3_11_sva_25;
  reg [2:0] act_regs_data_3_11_sva_24_22;
  reg act_regs_data_0_3_sva_25;
  reg [2:0] act_regs_data_0_3_sva_24_22;
  reg act_regs_data_3_12_sva_25;
  reg [2:0] act_regs_data_3_12_sva_24_22;
  reg act_regs_data_0_2_sva_25;
  reg [2:0] act_regs_data_0_2_sva_24_22;
  reg act_regs_data_3_13_sva_25;
  reg [2:0] act_regs_data_3_13_sva_24_22;
  reg act_regs_data_3_14_sva_25;
  reg [2:0] act_regs_data_3_14_sva_24_22;
  reg act_regs_data_3_15_sva_25;
  reg [2:0] act_regs_data_3_15_sva_24_22;
  wire ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_25_22_mx0w2_3;
  wire [2:0] ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_25_22_mx0w2_2_0;
  wire nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
  wire [2:0] nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
  wire nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
  wire [2:0] nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
  wire nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
  wire [2:0] nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
  wire nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
  wire [2:0] nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
  wire nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
  wire [2:0] nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
  wire nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
  wire [2:0] nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
  wire nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
  wire [2:0] nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
  wire nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
  wire [2:0] nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
  wire nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
  wire [2:0] nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
  wire nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
  wire [2:0] nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
  wire nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
  wire [2:0] nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
  wire nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
  wire [2:0] nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
  wire nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
  wire [2:0] nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
  wire nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
  wire [2:0] nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
  wire nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
  wire [2:0] nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
  wire nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
  wire [2:0] nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
  wire ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_25;
  wire [2:0] ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_24_22;
  reg rva_out_reg_data_39_32_sva_dfm_3_3;
  reg [2:0] rva_out_reg_data_39_32_sva_dfm_3_2_0;
  reg rva_out_reg_data_29_24_sva_dfm_3_3;
  reg [2:0] rva_out_reg_data_29_24_sva_dfm_3_2_0;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25;
  reg [2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25;
  reg [2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25;
  reg [2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25;
  reg [2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25;
  reg [2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25;
  reg [2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25;
  reg [2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25;
  reg [2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25;
  reg [2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25;
  reg [2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25;
  reg [2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25;
  reg [2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25;
  reg [2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25;
  reg [2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25;
  reg [2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22;
  reg nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25;
  reg [2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22;
  reg reg_ActUnit_RunInst_case_15_nv_scvector_cctor_data_0_ftd_rsp_0;
  reg [2:0] reg_ActUnit_RunInst_case_15_nv_scvector_cctor_data_0_ftd_rsp_1;
  reg reg_nv_scvector_cctor_nv_scvector_6_for_2_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0;
  reg [2:0] reg_nv_scvector_cctor_nv_scvector_6_for_2_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1;
  reg reg_nv_scvector_cctor_nv_scvector_6_for_3_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0;
  reg [2:0] reg_nv_scvector_cctor_nv_scvector_6_for_3_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1;
  reg reg_nv_scvector_cctor_nv_scvector_6_for_4_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0;
  reg [2:0] reg_nv_scvector_cctor_nv_scvector_6_for_4_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1;
  reg reg_nv_scvector_cctor_nv_scvector_6_for_5_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0;
  reg [2:0] reg_nv_scvector_cctor_nv_scvector_6_for_5_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1;
  reg reg_nv_scvector_cctor_nv_scvector_6_for_6_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0;
  reg [2:0] reg_nv_scvector_cctor_nv_scvector_6_for_6_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1;
  reg reg_nv_scvector_cctor_nv_scvector_6_for_7_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0;
  reg [2:0] reg_nv_scvector_cctor_nv_scvector_6_for_7_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1;
  reg reg_nv_scvector_cctor_nv_scvector_6_for_8_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0;
  reg [2:0] reg_nv_scvector_cctor_nv_scvector_6_for_8_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1;
  reg reg_nv_scvector_cctor_nv_scvector_6_for_9_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0;
  reg [2:0] reg_nv_scvector_cctor_nv_scvector_6_for_9_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1;
  reg reg_nv_scvector_cctor_nv_scvector_6_for_10_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0;
  reg [2:0] reg_nv_scvector_cctor_nv_scvector_6_for_10_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1;
  reg reg_nv_scvector_cctor_nv_scvector_6_for_11_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0;
  reg [2:0] reg_nv_scvector_cctor_nv_scvector_6_for_11_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1;
  reg reg_nv_scvector_cctor_nv_scvector_6_for_12_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0;
  reg [2:0] reg_nv_scvector_cctor_nv_scvector_6_for_12_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1;
  reg reg_nv_scvector_cctor_nv_scvector_6_for_13_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0;
  reg [2:0] reg_nv_scvector_cctor_nv_scvector_6_for_13_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1;
  reg reg_nv_scvector_cctor_nv_scvector_6_for_14_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0;
  reg [2:0] reg_nv_scvector_cctor_nv_scvector_6_for_14_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1;
  reg reg_nv_scvector_cctor_nv_scvector_6_for_15_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0;
  reg [2:0] reg_nv_scvector_cctor_nv_scvector_6_for_15_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1;
  reg reg_nv_scvector_cctor_nv_scvector_6_for_16_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0;
  reg [2:0] reg_nv_scvector_cctor_nv_scvector_6_for_16_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1;
  reg reg_ActUnit_RunInst_case_14_nv_scvector_cctor_data_0_1_ftd_rsp_0;
  reg [2:0] reg_ActUnit_RunInst_case_14_nv_scvector_cctor_data_0_1_ftd_rsp_1;
  reg reg_nv_scvector_cctor_nv_scvector_5_for_2_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0;
  reg [2:0] reg_nv_scvector_cctor_nv_scvector_5_for_2_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1;
  reg reg_nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0;
  reg [2:0] reg_nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1;
  reg reg_nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0;
  reg [2:0] reg_nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1;
  reg reg_nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0;
  reg [2:0] reg_nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1;
  reg reg_nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0;
  reg [2:0] reg_nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1;
  reg reg_nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0;
  reg [2:0] reg_nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1;
  reg reg_nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0;
  reg [2:0] reg_nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1;
  reg reg_nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0;
  reg [2:0] reg_nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1;
  reg reg_nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0;
  reg [2:0] reg_nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1;
  reg reg_nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0;
  reg [2:0] reg_nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1;
  reg reg_nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0;
  reg [2:0] reg_nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1;
  reg reg_nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0;
  reg [2:0] reg_nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1;
  reg reg_nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0;
  reg [2:0] reg_nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1;
  reg reg_nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0;
  reg [2:0] reg_nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1;
  reg reg_nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0;
  reg [2:0] reg_nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1;
  reg reg_Tanh_for_y_25_0_lpi_1_dfm_1_ftd;
  reg [2:0] reg_Tanh_for_y_25_0_lpi_1_dfm_1_ftd_1;
  reg reg_Tanh_for_y_25_0_15_lpi_1_dfm_1_ftd;
  reg [2:0] reg_Tanh_for_y_25_0_15_lpi_1_dfm_1_ftd_1;
  reg reg_Tanh_for_y_25_0_14_lpi_1_dfm_1_ftd;
  reg [2:0] reg_Tanh_for_y_25_0_14_lpi_1_dfm_1_ftd_1;
  reg reg_Tanh_for_y_25_0_13_lpi_1_dfm_1_ftd;
  reg [2:0] reg_Tanh_for_y_25_0_13_lpi_1_dfm_1_ftd_1;
  reg reg_Tanh_for_y_25_0_12_lpi_1_dfm_1_ftd;
  reg [2:0] reg_Tanh_for_y_25_0_12_lpi_1_dfm_1_ftd_1;
  reg reg_Tanh_for_y_25_0_11_lpi_1_dfm_1_ftd;
  reg [2:0] reg_Tanh_for_y_25_0_11_lpi_1_dfm_1_ftd_1;
  reg reg_Tanh_for_y_25_0_10_lpi_1_dfm_1_ftd;
  reg [2:0] reg_Tanh_for_y_25_0_10_lpi_1_dfm_1_ftd_1;
  reg reg_Tanh_for_y_25_0_9_lpi_1_dfm_1_ftd;
  reg [2:0] reg_Tanh_for_y_25_0_9_lpi_1_dfm_1_ftd_1;
  reg reg_Tanh_for_y_25_0_8_lpi_1_dfm_1_ftd;
  reg [2:0] reg_Tanh_for_y_25_0_8_lpi_1_dfm_1_ftd_1;
  reg reg_Tanh_for_y_25_0_7_lpi_1_dfm_1_ftd;
  reg [2:0] reg_Tanh_for_y_25_0_7_lpi_1_dfm_1_ftd_1;
  reg reg_Tanh_for_y_25_0_6_lpi_1_dfm_1_ftd;
  reg [2:0] reg_Tanh_for_y_25_0_6_lpi_1_dfm_1_ftd_1;
  reg reg_Tanh_for_y_25_0_5_lpi_1_dfm_1_ftd;
  reg [2:0] reg_Tanh_for_y_25_0_5_lpi_1_dfm_1_ftd_1;
  reg reg_Tanh_for_y_25_0_4_lpi_1_dfm_1_ftd;
  reg [2:0] reg_Tanh_for_y_25_0_4_lpi_1_dfm_1_ftd_1;
  reg reg_Tanh_for_y_25_0_3_lpi_1_dfm_1_ftd;
  reg [2:0] reg_Tanh_for_y_25_0_3_lpi_1_dfm_1_ftd_1;
  reg reg_Tanh_for_y_25_0_2_lpi_1_dfm_1_ftd;
  reg [2:0] reg_Tanh_for_y_25_0_2_lpi_1_dfm_1_ftd_1;
  reg reg_Tanh_for_y_25_0_1_lpi_1_dfm_1_ftd;
  reg [2:0] reg_Tanh_for_y_25_0_1_lpi_1_dfm_1_ftd_1;
  reg reg_act_write_data_data_0_15_2_ftd;
  reg [2:0] reg_act_write_data_data_0_15_2_ftd_1;
  reg reg_act_write_data_data_0_0_2_ftd;
  reg [2:0] reg_act_write_data_data_0_0_2_ftd_1;
  wire [3:0] Silu_for_11_else_else_else_else_if_acc_sdt;
  wire [4:0] nl_Silu_for_11_else_else_else_else_if_acc_sdt;
  wire act_config_output_counter_and_3_ssc;
  wire act_config_output_counter_and_2_ssc;
  reg act_config_output_counter_sva_3;
  reg [2:0] act_config_output_counter_sva_2_0;
  reg Relu_for_y_qr_30_0_1_lpi_1_dfm_25;
  reg [2:0] Relu_for_y_qr_30_0_1_lpi_1_dfm_24_22;
  reg Relu_for_y_qr_30_0_2_lpi_1_dfm_25;
  reg [2:0] Relu_for_y_qr_30_0_2_lpi_1_dfm_24_22;
  reg Relu_for_y_qr_30_0_3_lpi_1_dfm_25;
  reg [2:0] Relu_for_y_qr_30_0_3_lpi_1_dfm_24_22;
  reg Relu_for_y_qr_30_0_4_lpi_1_dfm_25;
  reg [2:0] Relu_for_y_qr_30_0_4_lpi_1_dfm_24_22;
  reg Relu_for_y_qr_30_0_5_lpi_1_dfm_25;
  reg [2:0] Relu_for_y_qr_30_0_5_lpi_1_dfm_24_22;
  reg Relu_for_y_qr_30_0_6_lpi_1_dfm_25;
  reg [2:0] Relu_for_y_qr_30_0_6_lpi_1_dfm_24_22;
  reg Relu_for_y_qr_30_0_7_lpi_1_dfm_25;
  reg [2:0] Relu_for_y_qr_30_0_7_lpi_1_dfm_24_22;
  reg Relu_for_y_qr_30_0_8_lpi_1_dfm_25;
  reg [2:0] Relu_for_y_qr_30_0_8_lpi_1_dfm_24_22;
  reg Relu_for_y_qr_30_0_9_lpi_1_dfm_25;
  reg [2:0] Relu_for_y_qr_30_0_9_lpi_1_dfm_24_22;
  reg Relu_for_y_qr_30_0_10_lpi_1_dfm_25;
  reg [2:0] Relu_for_y_qr_30_0_10_lpi_1_dfm_24_22;
  reg Relu_for_y_qr_30_0_11_lpi_1_dfm_25;
  reg [2:0] Relu_for_y_qr_30_0_11_lpi_1_dfm_24_22;
  reg Relu_for_y_qr_30_0_12_lpi_1_dfm_25;
  reg [2:0] Relu_for_y_qr_30_0_12_lpi_1_dfm_24_22;
  reg Relu_for_y_qr_30_0_13_lpi_1_dfm_25;
  reg [2:0] Relu_for_y_qr_30_0_13_lpi_1_dfm_24_22;
  reg Relu_for_y_qr_30_0_14_lpi_1_dfm_25;
  reg [2:0] Relu_for_y_qr_30_0_14_lpi_1_dfm_24_22;
  reg Relu_for_y_qr_30_0_15_lpi_1_dfm_25;
  reg [2:0] Relu_for_y_qr_30_0_15_lpi_1_dfm_24_22;
  reg Relu_for_y_qr_30_0_lpi_1_dfm_25;
  reg [2:0] Relu_for_y_qr_30_0_lpi_1_dfm_24_22;
  reg act_write_data_data_0_7_sva_25;
  reg [2:0] act_write_data_data_0_7_sva_24_22;
  reg act_write_data_data_0_8_sva_25;
  reg [2:0] act_write_data_data_0_8_sva_24_22;
  reg act_write_data_data_0_6_sva_25;
  reg [2:0] act_write_data_data_0_6_sva_24_22;
  reg act_write_data_data_0_9_sva_25;
  reg [2:0] act_write_data_data_0_9_sva_24_22;
  reg act_write_data_data_0_5_sva_25;
  reg [2:0] act_write_data_data_0_5_sva_24_22;
  reg act_write_data_data_0_10_sva_25;
  reg [2:0] act_write_data_data_0_10_sva_24_22;
  reg act_write_data_data_0_4_sva_25;
  reg [2:0] act_write_data_data_0_4_sva_24_22;
  reg act_write_data_data_0_11_sva_25;
  reg [2:0] act_write_data_data_0_11_sva_24_22;
  reg act_write_data_data_0_3_sva_25;
  reg [2:0] act_write_data_data_0_3_sva_24_22;
  reg act_write_data_data_0_12_sva_25;
  reg [2:0] act_write_data_data_0_12_sva_24_22;
  reg act_write_data_data_0_2_sva_25;
  reg [2:0] act_write_data_data_0_2_sva_24_22;
  reg act_write_data_data_0_13_sva_25;
  reg [2:0] act_write_data_data_0_13_sva_24_22;
  reg act_write_data_data_0_1_sva_25;
  reg [2:0] act_write_data_data_0_1_sva_24_22;
  reg act_write_data_data_0_14_sva_25;
  reg [2:0] act_write_data_data_0_14_sva_24_22;
  reg reg_act_config_output_counter_sva_dfm_3_ftd_1_3;
  reg [2:0] reg_act_config_output_counter_sva_dfm_3_ftd_1_2_0;

  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb;
  wire pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_prb_1;
  wire pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_1;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_1;
  wire pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_1;
  wire mux_330_nl;
  wire or_866_nl;
  wire mux_340_nl;
  wire mux_339_nl;
  wire mux_338_nl;
  wire mux_337_nl;
  wire or_872_nl;
  wire or_871_nl;
  wire mux_336_nl;
  wire mux_335_nl;
  wire nor_143_nl;
  wire nor_142_nl;
  wire mux_350_nl;
  wire mux_349_nl;
  wire mux_348_nl;
  wire mux_347_nl;
  wire or_877_nl;
  wire or_876_nl;
  wire mux_346_nl;
  wire mux_345_nl;
  wire nor_147_nl;
  wire nor_146_nl;
  wire mux_360_nl;
  wire mux_359_nl;
  wire mux_358_nl;
  wire mux_357_nl;
  wire or_882_nl;
  wire or_881_nl;
  wire mux_356_nl;
  wire mux_355_nl;
  wire nor_151_nl;
  wire nor_150_nl;
  wire mux_370_nl;
  wire mux_369_nl;
  wire mux_368_nl;
  wire mux_367_nl;
  wire or_887_nl;
  wire or_886_nl;
  wire mux_366_nl;
  wire mux_365_nl;
  wire nor_155_nl;
  wire nor_154_nl;
  wire mux_380_nl;
  wire mux_379_nl;
  wire mux_378_nl;
  wire mux_377_nl;
  wire or_892_nl;
  wire or_891_nl;
  wire mux_376_nl;
  wire mux_375_nl;
  wire nor_159_nl;
  wire nor_158_nl;
  wire mux_390_nl;
  wire mux_389_nl;
  wire mux_388_nl;
  wire mux_387_nl;
  wire or_897_nl;
  wire or_896_nl;
  wire mux_386_nl;
  wire mux_385_nl;
  wire nor_163_nl;
  wire nor_162_nl;
  wire mux_400_nl;
  wire mux_399_nl;
  wire mux_398_nl;
  wire mux_397_nl;
  wire or_902_nl;
  wire or_901_nl;
  wire mux_396_nl;
  wire mux_395_nl;
  wire nor_167_nl;
  wire nor_166_nl;
  wire mux_410_nl;
  wire mux_409_nl;
  wire mux_408_nl;
  wire mux_407_nl;
  wire or_907_nl;
  wire or_906_nl;
  wire mux_406_nl;
  wire mux_405_nl;
  wire nor_171_nl;
  wire nor_170_nl;
  wire mux_412_nl;
  wire and_1658_nl;
  wire nor_431_nl;
  wire mux_413_nl;
  wire and_1661_nl;
  wire nor_432_nl;
  wire mux_414_nl;
  wire and_1664_nl;
  wire nor_433_nl;
  wire mux_415_nl;
  wire and_1667_nl;
  wire nor_434_nl;
  wire mux_416_nl;
  wire and_1670_nl;
  wire nor_435_nl;
  wire mux_417_nl;
  wire and_1673_nl;
  wire nor_436_nl;
  wire mux_418_nl;
  wire and_1676_nl;
  wire nor_437_nl;
  wire mux_419_nl;
  wire and_1679_nl;
  wire nor_438_nl;
  wire mux_420_nl;
  wire and_1682_nl;
  wire nor_439_nl;
  wire mux_421_nl;
  wire and_1685_nl;
  wire nor_440_nl;
  wire mux_422_nl;
  wire and_1688_nl;
  wire nor_441_nl;
  wire mux_423_nl;
  wire and_1691_nl;
  wire nor_442_nl;
  wire mux_424_nl;
  wire and_1694_nl;
  wire nor_443_nl;
  wire mux_425_nl;
  wire and_1697_nl;
  wire nor_444_nl;
  wire mux_426_nl;
  wire and_1701_nl;
  wire nor_445_nl;
  wire mux_427_nl;
  wire and_1704_nl;
  wire nor_446_nl;
  wire and_1122_nl;
  wire mux_103_nl;
  wire mux_102_nl;
  wire nor_223_nl;
  wire or_359_nl;
  wire nor_42_nl;
  wire while_else_1_while_else_1_nand_1_nl;
  wire mux_320_nl;
  wire mux_319_nl;
  wire and_1521_nl;
  wire mux_318_nl;
  wire or_695_nl;
  wire mux_317_nl;
  wire mux_316_nl;
  wire or_656_nl;
  wire mux_315_nl;
  wire mux_314_nl;
  wire or_692_nl;
  wire[4:0] and_1716_nl;
  wire[4:0] mux1h_1_nl;
  wire[4:0] Silu_for_Silu_for_and_22_nl;
  wire[4:0] Silu_for_else_Silu_for_else_mux1h_2_nl;
  wire Silu_for_else_nor_5_nl;
  wire not_2610_nl;
  wire[3:0] act_config_InstIncr_if_act_config_InstIncr_if_and_1_nl;
  wire act_config_InstIncr_if_not_9_nl;
  wire act_config_InstIncr_if_act_config_InstIncr_if_and_2_nl;
  wire[2:0] act_config_InstIncr_if_act_config_InstIncr_if_and_3_nl;
  wire act_config_InstIncr_if_not_10_nl;
  wire[4:0] act_config_InstIncr_act_config_InstIncr_and_1_nl;
  wire[4:0] operator_5_false_acc_nl;
  wire[5:0] nl_operator_5_false_acc_nl;
  wire act_config_InstIncr_if_not_7_nl;
  wire and_1276_nl;
  wire mux_622_nl;
  wire and_2331_nl;
  wire mux_621_nl;
  wire mux_620_nl;
  wire mux_619_nl;
  wire mux_618_nl;
  wire mux_617_nl;
  wire nor_1408_nl;
  wire nor_1409_nl;
  wire mux_616_nl;
  wire nor_1410_nl;
  wire nor_1411_nl;
  wire mux_615_nl;
  wire mux_614_nl;
  wire nor_1412_nl;
  wire nor_1413_nl;
  wire mux_613_nl;
  wire nor_1414_nl;
  wire nor_1415_nl;
  wire mux_612_nl;
  wire mux_611_nl;
  wire mux_610_nl;
  wire nor_1416_nl;
  wire nor_1417_nl;
  wire mux_609_nl;
  wire nor_1418_nl;
  wire nor_1419_nl;
  wire mux_608_nl;
  wire mux_607_nl;
  wire nor_1420_nl;
  wire nor_1421_nl;
  wire mux_606_nl;
  wire nor_1422_nl;
  wire nor_1423_nl;
  wire mux_605_nl;
  wire mux_604_nl;
  wire mux_603_nl;
  wire mux_602_nl;
  wire nor_1424_nl;
  wire nor_1425_nl;
  wire mux_601_nl;
  wire nor_1426_nl;
  wire nor_1427_nl;
  wire mux_600_nl;
  wire mux_599_nl;
  wire nor_1428_nl;
  wire nor_1429_nl;
  wire mux_598_nl;
  wire nor_1430_nl;
  wire nor_1431_nl;
  wire mux_597_nl;
  wire mux_596_nl;
  wire mux_595_nl;
  wire nor_1432_nl;
  wire nor_1433_nl;
  wire mux_594_nl;
  wire nor_1434_nl;
  wire nor_1435_nl;
  wire mux_593_nl;
  wire mux_592_nl;
  wire nor_1436_nl;
  wire nor_1437_nl;
  wire mux_591_nl;
  wire nor_1438_nl;
  wire nor_1439_nl;
  wire nor_1440_nl;
  wire mux_439_nl;
  wire[4:0] Silu_for_Silu_for_and_19_nl;
  wire[4:0] Silu_for_else_Silu_for_else_mux1h_1_nl;
  wire Silu_for_else_nor_3_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_121_nl;
  wire mux_631_nl;
  wire mux_630_nl;
  wire nor_1442_nl;
  wire mux_629_nl;
  wire and_2332_nl;
  wire nor_1443_nl;
  wire nor_1444_nl;
  wire or_1582_nl;
  wire[31:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_13_nl;
  wire[31:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_12_nl;
  wire[31:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_11_nl;
  wire[31:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_10_nl;
  wire[31:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_9_nl;
  wire[31:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_8_nl;
  wire[31:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_7_nl;
  wire[31:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_6_nl;
  wire[31:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_5_nl;
  wire[31:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_4_nl;
  wire[31:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_3_nl;
  wire[31:0] ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_nl;
  wire mux_442_nl;
  wire mux_441_nl;
  wire mux_440_nl;
  wire or_1306_nl;
  wire and_1647_nl;
  wire[1:0] and_1721_nl;
  wire[1:0] mux_572_nl;
  wire not_2612_nl;
  wire[7:0] and_1723_nl;
  wire[7:0] mux_573_nl;
  wire not_2614_nl;
  wire[7:0] and_1725_nl;
  wire[7:0] mux_574_nl;
  wire not_2616_nl;
  wire[7:0] and_1727_nl;
  wire[7:0] mux_575_nl;
  wire not_2618_nl;
  wire[7:0] and_1729_nl;
  wire[7:0] mux_576_nl;
  wire not_2620_nl;
  wire[7:0] and_1731_nl;
  wire[7:0] mux_577_nl;
  wire not_2622_nl;
  wire[7:0] and_1733_nl;
  wire[7:0] mux_578_nl;
  wire not_2624_nl;
  wire[7:0] and_1735_nl;
  wire[7:0] mux_579_nl;
  wire not_2626_nl;
  wire[7:0] and_1737_nl;
  wire[7:0] mux_580_nl;
  wire not_2628_nl;
  wire[7:0] and_1739_nl;
  wire[7:0] mux_581_nl;
  wire not_2630_nl;
  wire[7:0] and_1741_nl;
  wire[7:0] mux_582_nl;
  wire not_2632_nl;
  wire[6:0] and_1743_nl;
  wire[6:0] mux_583_nl;
  wire not_2634_nl;
  wire[6:0] and_1745_nl;
  wire[6:0] mux_584_nl;
  wire not_2636_nl;
  wire[2:0] and_1747_nl;
  wire[2:0] mux_585_nl;
  wire not_2638_nl;
  wire ActUnit_RunInst_switch_lp_mux_3_nl;
  wire ActUnit_RunInst_switch_lp_mux_4_nl;
  wire ActUnit_RunInst_switch_lp_mux_6_nl;
  wire ActUnit_RunInst_switch_lp_mux_8_nl;
  wire ActUnit_RunInst_switch_lp_mux_10_nl;
  wire ActUnit_RunInst_switch_lp_mux_12_nl;
  wire ActUnit_RunInst_switch_lp_mux_14_nl;
  wire ActUnit_RunInst_switch_lp_mux_16_nl;
  wire mux_443_nl;
  wire mux_444_nl;
  wire Tanh_for_or_2_nl;
  wire Tanh_for_nor_1_nl;
  wire Tanh_for_or_3_nl;
  wire Tanh_for_nor_2_nl;
  wire Tanh_for_or_4_nl;
  wire Tanh_for_nor_3_nl;
  wire Tanh_for_or_5_nl;
  wire Tanh_for_nor_4_nl;
  wire Tanh_for_or_6_nl;
  wire Tanh_for_nor_5_nl;
  wire Tanh_for_or_7_nl;
  wire Tanh_for_nor_6_nl;
  wire Tanh_for_or_8_nl;
  wire Tanh_for_nor_7_nl;
  wire Tanh_for_or_9_nl;
  wire Tanh_for_nor_8_nl;
  wire Tanh_for_or_10_nl;
  wire Tanh_for_nor_9_nl;
  wire Tanh_for_or_11_nl;
  wire Tanh_for_nor_10_nl;
  wire Tanh_for_or_12_nl;
  wire Tanh_for_nor_11_nl;
  wire Tanh_for_or_13_nl;
  wire Tanh_for_nor_12_nl;
  wire Tanh_for_or_14_nl;
  wire Tanh_for_nor_13_nl;
  wire Tanh_for_or_15_nl;
  wire Tanh_for_nor_14_nl;
  wire Tanh_for_or_16_nl;
  wire Tanh_for_nor_15_nl;
  wire Tanh_for_or_17_nl;
  wire Tanh_for_nor_16_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_43_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_59_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_14_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_41_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_58_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_13_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_39_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_57_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_12_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_37_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_56_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_11_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_35_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_55_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_10_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_33_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_54_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_9_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_31_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_53_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_8_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_29_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_52_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_7_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_27_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_51_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_6_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_25_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_50_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_5_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_23_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_49_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_4_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_21_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_48_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_3_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_19_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_47_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_2_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_17_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_46_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_1_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_15_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_45_nl;
  wire nv_scvector_cctor_nv_scvector_4_for_not_nl;
  wire ActUnit_RunInst_switch_lp_not_10_nl;
  wire ActUnit_RunInst_switch_lp_not_12_nl;
  wire ActUnit_RunInst_switch_lp_not_1_nl;
  wire[4:0] ActUnit_RunInst_case_2_for_ActUnit_RunInst_case_2_for_and_1_nl;
  wire ActUnit_RunInst_case_2_for_ActUnit_RunInst_case_2_for_and_2_nl;
  wire[2:0] ActUnit_RunInst_case_2_for_ActUnit_RunInst_case_2_for_and_4_nl;
  wire[21:0] ActUnit_RunInst_case_2_for_ActUnit_RunInst_case_2_for_and_3_nl;
  wire mux_665_nl;
  wire[4:0] act_write_data_data_act_write_data_data_act_write_data_data_mux_nl;
  wire not_3249_nl;
  wire act_write_data_data_act_write_data_data_act_write_data_data_mux_1_nl;
  wire[2:0] act_write_data_data_act_write_data_data_act_write_data_data_mux_42_nl;
  wire not_8967_nl;
  wire[21:0] act_write_data_data_act_write_data_data_act_write_data_data_mux_2_nl;
  wire not_2573_nl;
  wire mux_669_nl;
  wire mux_668_nl;
  wire or_1678_nl;
  wire[4:0] act_write_data_data_act_write_data_data_act_write_data_data_mux_3_nl;
  wire not_3247_nl;
  wire act_write_data_data_act_write_data_data_act_write_data_data_mux_4_nl;
  wire[2:0] act_write_data_data_act_write_data_data_act_write_data_data_mux_43_nl;
  wire not_8966_nl;
  wire[21:0] act_write_data_data_act_write_data_data_act_write_data_data_mux_5_nl;
  wire not_2571_nl;
  wire mux_675_nl;
  wire mux_674_nl;
  wire or_1690_nl;
  wire[4:0] act_write_data_data_act_write_data_data_act_write_data_data_mux_6_nl;
  wire not_3245_nl;
  wire act_write_data_data_act_write_data_data_act_write_data_data_mux_7_nl;
  wire[2:0] act_write_data_data_act_write_data_data_act_write_data_data_mux_44_nl;
  wire not_8965_nl;
  wire[21:0] act_write_data_data_act_write_data_data_act_write_data_data_mux_8_nl;
  wire not_2569_nl;
  wire mux_680_nl;
  wire[4:0] act_write_data_data_act_write_data_data_act_write_data_data_mux_9_nl;
  wire not_3243_nl;
  wire act_write_data_data_act_write_data_data_act_write_data_data_mux_10_nl;
  wire[2:0] act_write_data_data_act_write_data_data_act_write_data_data_mux_45_nl;
  wire not_8964_nl;
  wire[21:0] act_write_data_data_act_write_data_data_act_write_data_data_mux_11_nl;
  wire not_2567_nl;
  wire mux_683_nl;
  wire[4:0] act_write_data_data_act_write_data_data_act_write_data_data_mux_12_nl;
  wire not_3241_nl;
  wire act_write_data_data_act_write_data_data_act_write_data_data_mux_13_nl;
  wire[2:0] act_write_data_data_act_write_data_data_act_write_data_data_mux_46_nl;
  wire not_8963_nl;
  wire[21:0] act_write_data_data_act_write_data_data_act_write_data_data_mux_14_nl;
  wire not_2565_nl;
  wire mux_687_nl;
  wire mux_1529_nl;
  wire[4:0] act_write_data_data_act_write_data_data_act_write_data_data_mux_15_nl;
  wire not_3239_nl;
  wire act_write_data_data_act_write_data_data_act_write_data_data_mux_16_nl;
  wire[2:0] act_write_data_data_act_write_data_data_act_write_data_data_mux_47_nl;
  wire not_8962_nl;
  wire[21:0] act_write_data_data_act_write_data_data_act_write_data_data_mux_17_nl;
  wire not_2563_nl;
  wire mux_693_nl;
  wire mux_686_nl;
  wire[4:0] act_write_data_data_act_write_data_data_act_write_data_data_mux_18_nl;
  wire not_3237_nl;
  wire act_write_data_data_act_write_data_data_act_write_data_data_mux_19_nl;
  wire[2:0] act_write_data_data_act_write_data_data_act_write_data_data_mux_48_nl;
  wire not_8961_nl;
  wire[21:0] act_write_data_data_act_write_data_data_act_write_data_data_mux_20_nl;
  wire not_2561_nl;
  wire mux_698_nl;
  wire[4:0] act_write_data_data_act_write_data_data_act_write_data_data_mux_21_nl;
  wire not_3235_nl;
  wire act_write_data_data_act_write_data_data_act_write_data_data_mux_22_nl;
  wire[2:0] act_write_data_data_act_write_data_data_act_write_data_data_mux_49_nl;
  wire not_8960_nl;
  wire[21:0] act_write_data_data_act_write_data_data_act_write_data_data_mux_23_nl;
  wire not_2559_nl;
  wire mux_701_nl;
  wire[4:0] act_write_data_data_act_write_data_data_act_write_data_data_mux_24_nl;
  wire not_3233_nl;
  wire act_write_data_data_act_write_data_data_act_write_data_data_mux_25_nl;
  wire[2:0] act_write_data_data_act_write_data_data_act_write_data_data_mux_50_nl;
  wire not_8959_nl;
  wire[21:0] act_write_data_data_act_write_data_data_act_write_data_data_mux_26_nl;
  wire not_2557_nl;
  wire mux_705_nl;
  wire mux_704_nl;
  wire or_1774_nl;
  wire[4:0] act_write_data_data_act_write_data_data_act_write_data_data_mux_27_nl;
  wire not_3231_nl;
  wire act_write_data_data_act_write_data_data_act_write_data_data_mux_28_nl;
  wire[2:0] act_write_data_data_act_write_data_data_act_write_data_data_mux_51_nl;
  wire not_8958_nl;
  wire[21:0] act_write_data_data_act_write_data_data_act_write_data_data_mux_29_nl;
  wire not_2555_nl;
  wire mux_711_nl;
  wire mux_710_nl;
  wire or_1786_nl;
  wire[4:0] act_write_data_data_act_write_data_data_act_write_data_data_mux_30_nl;
  wire not_3229_nl;
  wire act_write_data_data_act_write_data_data_act_write_data_data_mux_31_nl;
  wire[2:0] act_write_data_data_act_write_data_data_act_write_data_data_mux_52_nl;
  wire not_8957_nl;
  wire[21:0] act_write_data_data_act_write_data_data_act_write_data_data_mux_32_nl;
  wire not_2553_nl;
  wire mux_716_nl;
  wire[4:0] act_write_data_data_act_write_data_data_act_write_data_data_mux_33_nl;
  wire not_3227_nl;
  wire act_write_data_data_act_write_data_data_act_write_data_data_mux_34_nl;
  wire[2:0] act_write_data_data_act_write_data_data_act_write_data_data_mux_53_nl;
  wire not_8956_nl;
  wire[21:0] act_write_data_data_act_write_data_data_act_write_data_data_mux_35_nl;
  wire not_2551_nl;
  wire mux_719_nl;
  wire[4:0] act_write_data_data_act_write_data_data_act_write_data_data_mux_36_nl;
  wire not_3225_nl;
  wire act_write_data_data_act_write_data_data_act_write_data_data_mux_37_nl;
  wire[2:0] act_write_data_data_act_write_data_data_act_write_data_data_mux_54_nl;
  wire not_8955_nl;
  wire[21:0] act_write_data_data_act_write_data_data_act_write_data_data_mux_38_nl;
  wire not_2549_nl;
  wire mux_723_nl;
  wire mux_722_nl;
  wire[4:0] act_write_data_data_act_write_data_data_act_write_data_data_mux_39_nl;
  wire not_3223_nl;
  wire act_write_data_data_act_write_data_data_act_write_data_data_mux_40_nl;
  wire[2:0] act_write_data_data_act_write_data_data_act_write_data_data_mux_55_nl;
  wire not_8954_nl;
  wire[21:0] act_write_data_data_act_write_data_data_act_write_data_data_mux_41_nl;
  wire not_2547_nl;
  wire ActUnit_CheckStart_if_ActUnit_CheckStart_if_and_nl;
  wire ActUnit_RunInst_switch_lp_or_1_nl;
  wire mux_445_nl;
  wire ActUnit_PushOutput_if_for_i_not_nl;
  wire[4:0] Silu_for_Silu_for_and_16_nl;
  wire[4:0] Silu_for_else_Silu_for_else_mux1h_nl;
  wire Silu_for_else_nor_1_nl;
  wire ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_5_nl;
  wire ActUnit_DecodeAxiRead_else_mux_1_nl;
  wire ActUnit_DecodeAxi_mux_93_nl;
  wire ActUnit_DecodeAxi_if_mux_91_nl;
  wire ActUnit_DecodeAxiRead_mux_33_nl;
  wire act_config_ActConfigRead_mux_19_nl;
  wire act_config_ActConfigRead_else_mux_19_nl;
  wire act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_24_nl;
  wire ActUnit_DecodeAxi_mux_94_nl;
  wire ActUnit_DecodeAxi_if_mux_89_nl;
  wire ActUnit_DecodeAxiRead_mux_31_nl;
  wire act_config_ActConfigRead_mux_17_nl;
  wire act_config_ActConfigRead_else_mux_17_nl;
  wire act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_18_nl;
  wire[4:0] act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_22_nl;
  wire ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_7_nl;
  wire ActUnit_DecodeAxiRead_else_mux_3_nl;
  wire mux_433_nl;
  wire[25:0] Silu_for_1_else_else_else_if_acc_nl;
  wire[26:0] nl_Silu_for_1_else_else_else_if_acc_nl;
  wire[21:0] and_1749_nl;
  wire[21:0] mux_1495_nl;
  wire not_2640_nl;
  wire[25:0] Silu_for_2_else_else_else_if_acc_nl;
  wire[26:0] nl_Silu_for_2_else_else_else_if_acc_nl;
  wire[21:0] and_1752_nl;
  wire[21:0] mux1h_3_nl;
  wire and_1452_nl;
  wire not_2642_nl;
  wire[25:0] Silu_for_3_else_else_else_if_acc_nl;
  wire[26:0] nl_Silu_for_3_else_else_else_if_acc_nl;
  wire[21:0] and_1756_nl;
  wire[21:0] mux_1496_nl;
  wire not_2644_nl;
  wire[25:0] Silu_for_4_else_else_else_if_acc_nl;
  wire[26:0] nl_Silu_for_4_else_else_else_if_acc_nl;
  wire[21:0] and_1759_nl;
  wire[21:0] mux_1497_nl;
  wire not_2646_nl;
  wire[25:0] Silu_for_5_else_else_else_if_acc_nl;
  wire[26:0] nl_Silu_for_5_else_else_else_if_acc_nl;
  wire[21:0] and_1762_nl;
  wire[21:0] mux_1498_nl;
  wire not_2648_nl;
  wire[25:0] Silu_for_6_else_else_else_if_acc_nl;
  wire[26:0] nl_Silu_for_6_else_else_else_if_acc_nl;
  wire[21:0] and_1765_nl;
  wire[21:0] mux_1499_nl;
  wire not_2650_nl;
  wire[25:0] Silu_for_7_else_else_else_if_acc_nl;
  wire[26:0] nl_Silu_for_7_else_else_else_if_acc_nl;
  wire[21:0] and_1768_nl;
  wire[21:0] mux_1500_nl;
  wire not_2652_nl;
  wire[25:0] Silu_for_8_else_else_else_if_acc_nl;
  wire[26:0] nl_Silu_for_8_else_else_else_if_acc_nl;
  wire[21:0] and_1771_nl;
  wire[21:0] mux_1501_nl;
  wire not_2654_nl;
  wire[25:0] Silu_for_9_else_else_else_if_acc_nl;
  wire[26:0] nl_Silu_for_9_else_else_else_if_acc_nl;
  wire[21:0] and_1774_nl;
  wire[21:0] mux_1502_nl;
  wire not_2656_nl;
  wire mux_125_nl;
  wire and_1577_nl;
  wire mux_126_nl;
  wire and_1578_nl;
  wire mux_127_nl;
  wire and_1579_nl;
  wire mux_128_nl;
  wire and_1580_nl;
  wire mux_129_nl;
  wire and_1581_nl;
  wire mux_130_nl;
  wire and_1582_nl;
  wire mux_131_nl;
  wire and_1583_nl;
  wire mux_132_nl;
  wire and_1584_nl;
  wire mux_133_nl;
  wire and_1585_nl;
  wire mux_134_nl;
  wire and_1586_nl;
  wire mux_135_nl;
  wire and_1587_nl;
  wire mux_136_nl;
  wire and_1588_nl;
  wire mux_137_nl;
  wire and_1589_nl;
  wire mux_138_nl;
  wire and_1590_nl;
  wire mux_139_nl;
  wire and_1591_nl;
  wire mux_140_nl;
  wire and_1592_nl;
  wire mux_141_nl;
  wire and_1593_nl;
  wire mux_142_nl;
  wire and_1594_nl;
  wire mux_143_nl;
  wire and_1595_nl;
  wire mux_144_nl;
  wire and_1596_nl;
  wire mux_145_nl;
  wire and_1597_nl;
  wire mux_146_nl;
  wire and_1598_nl;
  wire mux_147_nl;
  wire and_1599_nl;
  wire mux_148_nl;
  wire and_1600_nl;
  wire mux_149_nl;
  wire and_1601_nl;
  wire mux_150_nl;
  wire and_1602_nl;
  wire mux_151_nl;
  wire and_1603_nl;
  wire mux_152_nl;
  wire and_1604_nl;
  wire mux_153_nl;
  wire and_1605_nl;
  wire mux_154_nl;
  wire and_1606_nl;
  wire mux_155_nl;
  wire and_1607_nl;
  wire mux_156_nl;
  wire and_1608_nl;
  wire[1:0] ActUnit_DecodeAxiWrite_if_mux_5_nl;
  wire[1:0] ActUnit_DecodeAxiWrite_if_mux_7_nl;
  wire[1:0] ActUnit_DecodeAxiWrite_if_mux_9_nl;
  wire[1:0] ActUnit_DecodeAxiWrite_if_mux_11_nl;
  wire[1:0] ActUnit_DecodeAxiWrite_if_mux_13_nl;
  wire[1:0] ActUnit_DecodeAxiWrite_if_mux_15_nl;
  wire[1:0] ActUnit_DecodeAxiWrite_if_mux_17_nl;
  wire[1:0] ActUnit_DecodeAxiWrite_if_mux_19_nl;
  wire[1:0] ActUnit_DecodeAxiWrite_if_mux_21_nl;
  wire[1:0] ActUnit_DecodeAxiWrite_if_mux_23_nl;
  wire[1:0] ActUnit_DecodeAxiWrite_if_mux_25_nl;
  wire[1:0] ActUnit_DecodeAxiWrite_if_mux_27_nl;
  wire[1:0] ActUnit_DecodeAxiWrite_if_mux_29_nl;
  wire[1:0] ActUnit_DecodeAxiWrite_if_mux_31_nl;
  wire[1:0] ActUnit_DecodeAxiWrite_if_mux_33_nl;
  wire[1:0] ActUnit_DecodeAxiWrite_if_mux_35_nl;
  wire act_regs_data_mux_320_nl;
  wire act_regs_data_or_64_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_231_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_229_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_230_nl;
  wire act_regs_data_mux_324_nl;
  wire act_regs_data_or_65_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_291_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_4_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_289_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_290_nl;
  wire act_regs_data_mux_328_nl;
  wire act_regs_data_or_66_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_279_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_8_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_277_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_278_nl;
  wire act_regs_data_mux_332_nl;
  wire act_regs_data_or_67_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_267_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_12_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_265_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_266_nl;
  wire act_regs_data_mux_336_nl;
  wire act_regs_data_or_68_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_255_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_16_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_253_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_254_nl;
  wire act_regs_data_mux_340_nl;
  wire act_regs_data_or_69_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_243_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_20_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_241_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_242_nl;
  wire act_regs_data_mux_344_nl;
  wire act_regs_data_or_70_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_132_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_24_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_130_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_131_nl;
  wire act_regs_data_mux_348_nl;
  wire act_regs_data_or_71_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_219_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_28_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_217_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_218_nl;
  wire act_regs_data_mux_352_nl;
  wire act_regs_data_or_72_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_204_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_32_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_202_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_203_nl;
  wire act_regs_data_mux_356_nl;
  wire act_regs_data_or_73_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_192_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_36_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_190_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_191_nl;
  wire act_regs_data_mux_360_nl;
  wire act_regs_data_or_74_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_180_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_40_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_178_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_179_nl;
  wire act_regs_data_mux_364_nl;
  wire act_regs_data_or_75_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_168_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_44_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_166_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_167_nl;
  wire act_regs_data_mux_368_nl;
  wire act_regs_data_or_76_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_156_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_48_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_154_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_155_nl;
  wire act_regs_data_mux_372_nl;
  wire act_regs_data_or_77_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_144_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_52_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_142_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_143_nl;
  wire act_regs_data_mux_376_nl;
  wire act_regs_data_or_78_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_303_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_56_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_301_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_302_nl;
  wire act_regs_data_mux_380_nl;
  wire act_regs_data_or_79_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_120_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_60_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_118_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_119_nl;
  wire act_regs_data_mux_384_nl;
  wire act_regs_data_or_80_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_225_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_64_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_223_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_224_nl;
  wire act_regs_data_mux_388_nl;
  wire act_regs_data_or_81_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_285_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_68_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_283_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_284_nl;
  wire act_regs_data_mux_392_nl;
  wire act_regs_data_or_82_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_273_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_72_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_271_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_272_nl;
  wire act_regs_data_mux_396_nl;
  wire act_regs_data_or_83_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_261_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_76_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_259_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_260_nl;
  wire act_regs_data_mux_400_nl;
  wire act_regs_data_or_84_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_249_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_80_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_247_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_248_nl;
  wire act_regs_data_mux_404_nl;
  wire act_regs_data_or_85_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_237_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_84_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_235_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_236_nl;
  wire act_regs_data_mux_408_nl;
  wire act_regs_data_or_86_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_126_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_88_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_124_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_125_nl;
  wire act_regs_data_mux_412_nl;
  wire act_regs_data_or_87_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_213_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_92_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_211_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_212_nl;
  wire act_regs_data_mux_416_nl;
  wire act_regs_data_or_88_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_198_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_96_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_196_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_197_nl;
  wire act_regs_data_mux_420_nl;
  wire act_regs_data_or_89_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_186_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_100_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_184_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_185_nl;
  wire act_regs_data_mux_424_nl;
  wire act_regs_data_or_90_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_174_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_104_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_172_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_173_nl;
  wire act_regs_data_mux_428_nl;
  wire act_regs_data_or_91_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_162_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_108_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_160_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_161_nl;
  wire act_regs_data_mux_432_nl;
  wire act_regs_data_or_92_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_150_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_112_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_148_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_149_nl;
  wire act_regs_data_mux_436_nl;
  wire act_regs_data_or_93_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_138_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_116_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_136_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_137_nl;
  wire act_regs_data_mux_440_nl;
  wire act_regs_data_or_94_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_297_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_120_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_295_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_296_nl;
  wire act_regs_data_mux_444_nl;
  wire act_regs_data_or_95_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_114_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_124_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_112_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_113_nl;
  wire act_regs_data_mux_448_nl;
  wire act_regs_data_or_96_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_222_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_128_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_220_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_221_nl;
  wire act_regs_data_mux_452_nl;
  wire act_regs_data_or_97_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_282_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_132_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_280_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_281_nl;
  wire act_regs_data_mux_456_nl;
  wire act_regs_data_or_98_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_270_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_136_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_268_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_269_nl;
  wire act_regs_data_mux_460_nl;
  wire act_regs_data_or_99_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_258_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_140_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_256_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_257_nl;
  wire act_regs_data_mux_464_nl;
  wire act_regs_data_or_100_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_246_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_144_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_244_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_245_nl;
  wire act_regs_data_mux_468_nl;
  wire act_regs_data_or_101_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_234_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_148_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_232_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_233_nl;
  wire act_regs_data_mux_472_nl;
  wire act_regs_data_or_102_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_129_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_152_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_127_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_128_nl;
  wire act_regs_data_mux_476_nl;
  wire act_regs_data_or_103_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_210_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_156_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_208_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_209_nl;
  wire act_regs_data_mux_480_nl;
  wire act_regs_data_or_104_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_201_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_160_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_199_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_200_nl;
  wire act_regs_data_mux_484_nl;
  wire act_regs_data_or_105_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_189_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_164_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_187_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_188_nl;
  wire act_regs_data_mux_488_nl;
  wire act_regs_data_or_106_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_177_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_168_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_175_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_176_nl;
  wire act_regs_data_mux_492_nl;
  wire act_regs_data_or_107_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_165_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_172_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_163_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_164_nl;
  wire act_regs_data_mux_496_nl;
  wire act_regs_data_or_108_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_153_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_176_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_151_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_152_nl;
  wire act_regs_data_mux_500_nl;
  wire act_regs_data_or_109_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_141_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_180_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_139_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_140_nl;
  wire act_regs_data_mux_504_nl;
  wire act_regs_data_or_110_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_294_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_184_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_292_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_293_nl;
  wire act_regs_data_mux_508_nl;
  wire act_regs_data_or_111_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_117_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_188_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_115_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_116_nl;
  wire act_regs_data_mux_512_nl;
  wire act_regs_data_or_112_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_228_nl;
  wire ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_192_nl;
  wire[4:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_226_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_227_nl;
  wire ActUnit_DecodeAxiWrite_mux_4_nl;
  wire act_config_ActConfigWrite_mux_1_nl;
  wire while_and_64_nl;
  wire mux_451_nl;
  wire or_1426_nl;
  wire and_2363_nl;
  wire or_1866_nl;
  wire mux_18_nl;
  wire mux_17_nl;
  wire and_nl;
  wire mux_16_nl;
  wire nor_nl;
  wire Silu_for_else_mux_32_nl;
  wire[1:0] Silu_for_else_Silu_for_else_mux1h_39_nl;
  wire[19:0] Silu_for_else_Silu_for_else_mux1h_48_nl;
  wire Silu_for_else_mux_33_nl;
  wire[1:0] Silu_for_else_Silu_for_else_mux1h_38_nl;
  wire[19:0] Silu_for_else_Silu_for_else_mux1h_50_nl;
  wire Silu_for_else_mux_34_nl;
  wire[1:0] Silu_for_else_Silu_for_else_mux1h_37_nl;
  wire[19:0] Silu_for_else_Silu_for_else_mux1h_52_nl;
  wire Silu_for_else_mux_35_nl;
  wire[1:0] Silu_for_else_Silu_for_else_mux1h_36_nl;
  wire[19:0] Silu_for_else_Silu_for_else_mux1h_54_nl;
  wire Silu_for_else_mux_36_nl;
  wire[1:0] Silu_for_else_Silu_for_else_mux1h_35_nl;
  wire[19:0] Silu_for_else_Silu_for_else_mux1h_56_nl;
  wire Silu_for_else_mux_37_nl;
  wire[1:0] Silu_for_else_Silu_for_else_mux1h_34_nl;
  wire[19:0] Silu_for_else_Silu_for_else_mux1h_58_nl;
  wire Silu_for_else_mux_38_nl;
  wire[1:0] Silu_for_else_Silu_for_else_mux1h_33_nl;
  wire[19:0] Silu_for_else_Silu_for_else_mux1h_60_nl;
  wire Silu_for_else_mux_39_nl;
  wire[1:0] Silu_for_else_Silu_for_else_mux1h_32_nl;
  wire[19:0] Silu_for_else_Silu_for_else_mux1h_62_nl;
  wire[4:0] ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_70_nl;
  wire[4:0] Silu_for_Silu_for_and_25_nl;
  wire[4:0] Silu_for_else_Silu_for_else_mux1h_3_nl;
  wire Silu_for_else_nor_7_nl;
  wire not_8877_nl;
  wire[4:0] ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_75_nl;
  wire[4:0] Silu_for_Silu_for_and_28_nl;
  wire[4:0] Silu_for_else_Silu_for_else_mux1h_4_nl;
  wire Silu_for_else_nor_9_nl;
  wire not_8878_nl;
  wire[4:0] ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_80_nl;
  wire[4:0] Silu_for_Silu_for_and_31_nl;
  wire[4:0] Silu_for_else_Silu_for_else_mux1h_5_nl;
  wire Silu_for_else_nor_11_nl;
  wire not_8879_nl;
  wire[4:0] ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_85_nl;
  wire[4:0] Silu_for_Silu_for_and_34_nl;
  wire[4:0] Silu_for_else_Silu_for_else_mux1h_6_nl;
  wire Silu_for_else_nor_13_nl;
  wire not_8880_nl;
  wire[4:0] ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_90_nl;
  wire[4:0] Silu_for_Silu_for_and_37_nl;
  wire[4:0] Silu_for_else_Silu_for_else_mux1h_7_nl;
  wire Silu_for_else_nor_15_nl;
  wire not_8881_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_123_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_mux_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_288_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_mux_1_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_135_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_mux_2_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_276_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_mux_3_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_300_nl;
  wire[4:0] ActUnit_PushOutput_if_output_port_reg_data_data_mux_4_nl;
  wire not_8882_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_mux_5_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_264_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_mux_6_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_147_nl;
  wire[4:0] ActUnit_PushOutput_if_output_port_reg_data_data_mux_7_nl;
  wire not_8883_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_mux_8_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_252_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_mux_9_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_159_nl;
  wire[4:0] ActUnit_PushOutput_if_output_port_reg_data_data_mux_10_nl;
  wire not_8884_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_mux_11_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_240_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_mux_12_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_171_nl;
  wire[4:0] ActUnit_PushOutput_if_output_port_reg_data_data_mux_13_nl;
  wire not_8885_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_mux_14_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_216_nl;
  wire[4:0] ActUnit_PushOutput_if_output_port_reg_data_data_mux_15_nl;
  wire not_8886_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_mux_16_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_183_nl;
  wire[4:0] ActUnit_PushOutput_if_output_port_reg_data_data_mux_17_nl;
  wire not_8888_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_mux_18_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_207_nl;
  wire[4:0] ActUnit_PushOutput_if_output_port_reg_data_data_mux_19_nl;
  wire not_8889_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_mux_20_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_195_nl;
  wire[4:0] ActUnit_PushOutput_if_output_port_reg_data_data_mux_21_nl;
  wire not_8890_nl;
  wire while_and_213_nl;
  wire while_while_mux1h_150_nl;
  wire while_and_214_nl;
  wire while_while_mux1h_153_nl;
  wire while_and_215_nl;
  wire while_while_mux1h_156_nl;
  wire while_and_216_nl;
  wire while_while_mux1h_159_nl;
  wire while_and_217_nl;
  wire while_while_mux1h_162_nl;
  wire while_and_218_nl;
  wire while_while_mux1h_165_nl;
  wire while_and_219_nl;
  wire while_while_mux1h_168_nl;
  wire while_and_220_nl;
  wire while_while_mux1h_171_nl;
  wire while_and_221_nl;
  wire while_while_mux1h_174_nl;
  wire while_and_222_nl;
  wire while_while_mux1h_177_nl;
  wire while_and_223_nl;
  wire while_while_mux1h_180_nl;
  wire while_and_224_nl;
  wire while_while_mux1h_183_nl;
  wire while_and_225_nl;
  wire while_while_mux1h_186_nl;
  wire while_and_226_nl;
  wire while_while_mux1h_189_nl;
  wire while_and_227_nl;
  wire while_while_mux1h_192_nl;
  wire while_and_228_nl;
  wire while_while_mux1h_195_nl;
  wire while_and_229_nl;
  wire while_while_mux1h_198_nl;
  wire while_and_230_nl;
  wire while_while_mux1h_201_nl;
  wire while_and_231_nl;
  wire while_while_mux1h_204_nl;
  wire while_and_232_nl;
  wire while_while_mux1h_207_nl;
  wire while_and_233_nl;
  wire while_while_mux1h_210_nl;
  wire while_and_234_nl;
  wire while_while_mux1h_213_nl;
  wire while_and_235_nl;
  wire while_while_mux1h_216_nl;
  wire while_and_236_nl;
  wire while_while_mux1h_219_nl;
  wire while_and_237_nl;
  wire while_while_mux1h_222_nl;
  wire while_and_238_nl;
  wire while_while_mux1h_225_nl;
  wire while_and_239_nl;
  wire while_while_mux1h_228_nl;
  wire while_and_240_nl;
  wire while_while_mux1h_231_nl;
  wire while_and_241_nl;
  wire while_while_mux1h_234_nl;
  wire while_and_242_nl;
  wire while_while_mux1h_237_nl;
  wire while_and_243_nl;
  wire while_while_mux1h_240_nl;
  wire while_and_244_nl;
  wire while_while_mux1h_243_nl;
  wire while_and_245_nl;
  wire while_while_mux1h_246_nl;
  wire while_and_246_nl;
  wire while_while_mux1h_249_nl;
  wire while_and_247_nl;
  wire while_while_mux1h_252_nl;
  wire while_and_248_nl;
  wire while_while_mux1h_255_nl;
  wire while_and_249_nl;
  wire while_while_mux1h_258_nl;
  wire while_and_250_nl;
  wire while_while_mux1h_261_nl;
  wire while_and_251_nl;
  wire while_while_mux1h_264_nl;
  wire while_and_252_nl;
  wire while_while_mux1h_267_nl;
  wire while_and_253_nl;
  wire while_while_mux1h_270_nl;
  wire while_and_254_nl;
  wire while_while_mux1h_273_nl;
  wire while_and_255_nl;
  wire while_while_mux1h_276_nl;
  wire while_and_256_nl;
  wire while_while_mux1h_279_nl;
  wire while_and_257_nl;
  wire while_while_mux1h_282_nl;
  wire while_and_258_nl;
  wire while_while_mux1h_285_nl;
  wire while_and_259_nl;
  wire while_while_mux1h_288_nl;
  wire while_and_260_nl;
  wire while_while_mux1h_291_nl;
  wire while_and_261_nl;
  wire while_while_mux1h_294_nl;
  wire while_and_262_nl;
  wire while_while_mux1h_297_nl;
  wire while_and_263_nl;
  wire while_while_mux1h_300_nl;
  wire while_and_264_nl;
  wire while_while_mux1h_303_nl;
  wire while_and_265_nl;
  wire while_while_mux1h_306_nl;
  wire while_and_266_nl;
  wire while_while_mux1h_309_nl;
  wire while_and_267_nl;
  wire while_while_mux1h_312_nl;
  wire while_and_268_nl;
  wire while_while_mux1h_315_nl;
  wire while_and_269_nl;
  wire while_while_mux1h_318_nl;
  wire while_and_270_nl;
  wire while_while_mux1h_321_nl;
  wire while_and_271_nl;
  wire while_while_mux1h_324_nl;
  wire while_and_272_nl;
  wire while_while_mux1h_327_nl;
  wire while_and_273_nl;
  wire while_while_mux1h_330_nl;
  wire while_and_274_nl;
  wire while_while_mux1h_333_nl;
  wire while_and_275_nl;
  wire while_while_mux1h_336_nl;
  wire while_and_276_nl;
  wire while_while_mux1h_339_nl;
  wire and_2391_nl;
  wire mux_770_nl;
  wire mux_772_nl;
  wire mux_775_nl;
  wire mux_778_nl;
  wire mux_781_nl;
  wire mux_784_nl;
  wire mux_787_nl;
  wire mux_790_nl;
  wire mux_793_nl;
  wire mux_797_nl;
  wire mux_796_nl;
  wire mux_801_nl;
  wire mux_800_nl;
  wire mux_805_nl;
  wire mux_804_nl;
  wire mux_809_nl;
  wire mux_808_nl;
  wire mux_813_nl;
  wire mux_812_nl;
  wire mux_817_nl;
  wire mux_816_nl;
  wire mux_821_nl;
  wire mux_820_nl;
  wire mux_825_nl;
  wire mux_824_nl;
  wire and_2427_nl;
  wire mux_826_nl;
  wire mux_828_nl;
  wire mux_831_nl;
  wire mux_834_nl;
  wire mux_837_nl;
  wire mux_840_nl;
  wire mux_843_nl;
  wire mux_846_nl;
  wire mux_849_nl;
  wire mux_853_nl;
  wire mux_852_nl;
  wire mux_857_nl;
  wire mux_856_nl;
  wire mux_861_nl;
  wire mux_860_nl;
  wire mux_865_nl;
  wire mux_864_nl;
  wire mux_869_nl;
  wire mux_868_nl;
  wire mux_873_nl;
  wire mux_872_nl;
  wire mux_877_nl;
  wire mux_876_nl;
  wire mux_881_nl;
  wire mux_880_nl;
  wire and_2463_nl;
  wire mux_882_nl;
  wire mux_884_nl;
  wire mux_887_nl;
  wire mux_890_nl;
  wire mux_893_nl;
  wire mux_896_nl;
  wire mux_899_nl;
  wire mux_902_nl;
  wire mux_905_nl;
  wire mux_909_nl;
  wire mux_908_nl;
  wire mux_913_nl;
  wire mux_912_nl;
  wire mux_917_nl;
  wire mux_916_nl;
  wire mux_921_nl;
  wire mux_920_nl;
  wire mux_925_nl;
  wire mux_924_nl;
  wire mux_929_nl;
  wire mux_928_nl;
  wire mux_933_nl;
  wire mux_932_nl;
  wire mux_937_nl;
  wire mux_936_nl;
  wire and_2499_nl;
  wire mux_938_nl;
  wire mux_940_nl;
  wire mux_943_nl;
  wire mux_946_nl;
  wire mux_949_nl;
  wire mux_952_nl;
  wire mux_955_nl;
  wire mux_958_nl;
  wire mux_961_nl;
  wire mux_965_nl;
  wire mux_964_nl;
  wire mux_969_nl;
  wire mux_968_nl;
  wire mux_973_nl;
  wire mux_972_nl;
  wire mux_977_nl;
  wire mux_976_nl;
  wire mux_981_nl;
  wire mux_980_nl;
  wire mux_985_nl;
  wire mux_984_nl;
  wire mux_989_nl;
  wire mux_988_nl;
  wire mux_993_nl;
  wire mux_992_nl;
  wire and_2535_nl;
  wire mux_994_nl;
  wire and_2571_nl;
  wire mux_1051_nl;
  wire and_2607_nl;
  wire mux_1122_nl;
  wire and_2643_nl;
  wire mux_1179_nl;
  wire act_config_InstIncr_mux_2_nl;
  wire act_config_InstIncr_if_act_config_InstIncr_if_and_nl;
  wire ActUnit_RunInst_switch_lp_nor_nl;
  wire[4:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_6_nl;
  wire[4:0] ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_and_18_nl;
  wire ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_nl;
  wire ActUnit_DecodeAxiWrite_else_not_17_nl;
  wire[31:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_8_nl;
  wire[31:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_9_nl;
  wire[31:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_10_nl;
  wire[31:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_11_nl;
  wire[31:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_12_nl;
  wire[31:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_13_nl;
  wire[31:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_14_nl;
  wire[31:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_15_nl;
  wire[31:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_16_nl;
  wire[31:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_17_nl;
  wire[31:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_18_nl;
  wire[31:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_19_nl;
  wire[31:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_20_nl;
  wire[31:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_21_nl;
  wire[31:0] ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_22_nl;
  wire while_mux_32_nl;
  wire[4:0] while_mux_427_nl;
  wire while_mux_428_nl;
  wire[2:0] while_mux_430_nl;
  wire[21:0] while_mux_429_nl;
  wire while_while_nand_nl;
  wire Silu_for_else_mux_40_nl;
  wire[1:0] Silu_for_else_Silu_for_else_mux1h_47_nl;
  wire[19:0] Silu_for_else_Silu_for_else_mux1h_64_nl;
  wire[4:0] Silu_for_else_Silu_for_else_mux1h_15_nl;
  wire Silu_for_else_nor_31_nl;
  wire Silu_for_else_mux_41_nl;
  wire[1:0] Silu_for_else_Silu_for_else_mux1h_46_nl;
  wire[19:0] Silu_for_else_Silu_for_else_mux1h_66_nl;
  wire[4:0] Silu_for_else_Silu_for_else_mux1h_14_nl;
  wire Silu_for_else_nor_29_nl;
  wire Silu_for_else_mux_42_nl;
  wire[1:0] Silu_for_else_Silu_for_else_mux1h_45_nl;
  wire[19:0] Silu_for_else_Silu_for_else_mux1h_68_nl;
  wire[4:0] Silu_for_else_Silu_for_else_mux1h_13_nl;
  wire Silu_for_else_nor_27_nl;
  wire Silu_for_else_mux_43_nl;
  wire[1:0] Silu_for_else_Silu_for_else_mux1h_44_nl;
  wire[19:0] Silu_for_else_Silu_for_else_mux1h_70_nl;
  wire[4:0] Silu_for_else_Silu_for_else_mux1h_12_nl;
  wire Silu_for_else_nor_25_nl;
  wire Silu_for_else_mux_44_nl;
  wire[1:0] Silu_for_else_Silu_for_else_mux1h_43_nl;
  wire[19:0] Silu_for_else_Silu_for_else_mux1h_72_nl;
  wire[4:0] Silu_for_else_Silu_for_else_mux1h_11_nl;
  wire Silu_for_else_nor_23_nl;
  wire Silu_for_else_mux_45_nl;
  wire[1:0] Silu_for_else_Silu_for_else_mux1h_42_nl;
  wire[19:0] Silu_for_else_Silu_for_else_mux1h_74_nl;
  wire[4:0] Silu_for_else_Silu_for_else_mux1h_10_nl;
  wire Silu_for_else_nor_21_nl;
  wire Silu_for_else_mux_46_nl;
  wire[1:0] Silu_for_else_Silu_for_else_mux1h_41_nl;
  wire[19:0] Silu_for_else_Silu_for_else_mux1h_76_nl;
  wire[4:0] Silu_for_else_Silu_for_else_mux1h_9_nl;
  wire Silu_for_else_nor_19_nl;
  wire Silu_for_else_mux_47_nl;
  wire[1:0] Silu_for_else_Silu_for_else_mux1h_40_nl;
  wire[19:0] Silu_for_else_Silu_for_else_mux1h_78_nl;
  wire[4:0] Silu_for_else_Silu_for_else_mux1h_8_nl;
  wire Silu_for_else_nor_17_nl;
  wire Gelu_for_else_Gelu_for_else_mux1h_15_nl;
  wire[21:0] Gelu_for_else_Gelu_for_else_mux1h_47_nl;
  wire Gelu_for_else_or_nl;
  wire[4:0] Gelu_for_else_Gelu_for_else_mux1h_31_nl;
  wire Gelu_for_else_Gelu_for_else_mux1h_63_nl;
  wire[2:0] Gelu_for_else_Gelu_for_else_mux1h_79_nl;
  wire Gelu_for_else_Gelu_for_else_mux1h_14_nl;
  wire[21:0] Gelu_for_else_Gelu_for_else_mux1h_46_nl;
  wire Gelu_for_else_or_1_nl;
  wire[4:0] Gelu_for_else_Gelu_for_else_mux1h_30_nl;
  wire Gelu_for_else_Gelu_for_else_mux1h_62_nl;
  wire[2:0] Gelu_for_else_Gelu_for_else_mux1h_78_nl;
  wire Gelu_for_else_Gelu_for_else_mux1h_13_nl;
  wire[21:0] Gelu_for_else_Gelu_for_else_mux1h_45_nl;
  wire Gelu_for_else_or_2_nl;
  wire[4:0] Gelu_for_else_Gelu_for_else_mux1h_29_nl;
  wire Gelu_for_else_Gelu_for_else_mux1h_61_nl;
  wire[2:0] Gelu_for_else_Gelu_for_else_mux1h_77_nl;
  wire Gelu_for_else_Gelu_for_else_mux1h_12_nl;
  wire[21:0] Gelu_for_else_Gelu_for_else_mux1h_44_nl;
  wire Gelu_for_else_or_3_nl;
  wire[4:0] Gelu_for_else_Gelu_for_else_mux1h_28_nl;
  wire Gelu_for_else_Gelu_for_else_mux1h_60_nl;
  wire[2:0] Gelu_for_else_Gelu_for_else_mux1h_76_nl;
  wire Gelu_for_else_Gelu_for_else_mux1h_11_nl;
  wire[21:0] Gelu_for_else_Gelu_for_else_mux1h_43_nl;
  wire Gelu_for_else_or_4_nl;
  wire[4:0] Gelu_for_else_Gelu_for_else_mux1h_27_nl;
  wire Gelu_for_else_Gelu_for_else_mux1h_59_nl;
  wire[2:0] Gelu_for_else_Gelu_for_else_mux1h_75_nl;
  wire Gelu_for_else_Gelu_for_else_mux1h_10_nl;
  wire[21:0] Gelu_for_else_Gelu_for_else_mux1h_42_nl;
  wire Gelu_for_else_or_5_nl;
  wire[4:0] Gelu_for_else_Gelu_for_else_mux1h_26_nl;
  wire Gelu_for_else_Gelu_for_else_mux1h_58_nl;
  wire[2:0] Gelu_for_else_Gelu_for_else_mux1h_74_nl;
  wire Gelu_for_else_Gelu_for_else_mux1h_9_nl;
  wire[21:0] Gelu_for_else_Gelu_for_else_mux1h_41_nl;
  wire Gelu_for_else_or_6_nl;
  wire[4:0] Gelu_for_else_Gelu_for_else_mux1h_25_nl;
  wire Gelu_for_else_Gelu_for_else_mux1h_57_nl;
  wire[2:0] Gelu_for_else_Gelu_for_else_mux1h_73_nl;
  wire Gelu_for_else_Gelu_for_else_mux1h_8_nl;
  wire[21:0] Gelu_for_else_Gelu_for_else_mux1h_40_nl;
  wire Gelu_for_else_or_7_nl;
  wire[4:0] Gelu_for_else_Gelu_for_else_mux1h_24_nl;
  wire Gelu_for_else_Gelu_for_else_mux1h_56_nl;
  wire[2:0] Gelu_for_else_Gelu_for_else_mux1h_72_nl;
  wire Gelu_for_else_Gelu_for_else_mux1h_7_nl;
  wire[21:0] Gelu_for_else_Gelu_for_else_mux1h_39_nl;
  wire Gelu_for_else_or_8_nl;
  wire[4:0] Gelu_for_else_Gelu_for_else_mux1h_23_nl;
  wire Gelu_for_else_Gelu_for_else_mux1h_55_nl;
  wire[2:0] Gelu_for_else_Gelu_for_else_mux1h_71_nl;
  wire Gelu_for_else_Gelu_for_else_mux1h_6_nl;
  wire[21:0] Gelu_for_else_Gelu_for_else_mux1h_38_nl;
  wire Gelu_for_else_or_9_nl;
  wire[4:0] Gelu_for_else_Gelu_for_else_mux1h_22_nl;
  wire Gelu_for_else_Gelu_for_else_mux1h_54_nl;
  wire[2:0] Gelu_for_else_Gelu_for_else_mux1h_70_nl;
  wire Gelu_for_else_Gelu_for_else_mux1h_5_nl;
  wire[21:0] Gelu_for_else_Gelu_for_else_mux1h_37_nl;
  wire Gelu_for_else_or_10_nl;
  wire[4:0] Gelu_for_else_Gelu_for_else_mux1h_21_nl;
  wire Gelu_for_else_Gelu_for_else_mux1h_53_nl;
  wire[2:0] Gelu_for_else_Gelu_for_else_mux1h_69_nl;
  wire Gelu_for_else_Gelu_for_else_mux1h_4_nl;
  wire[21:0] Gelu_for_else_Gelu_for_else_mux1h_36_nl;
  wire Gelu_for_else_or_11_nl;
  wire[4:0] Gelu_for_else_Gelu_for_else_mux1h_20_nl;
  wire Gelu_for_else_Gelu_for_else_mux1h_52_nl;
  wire[2:0] Gelu_for_else_Gelu_for_else_mux1h_68_nl;
  wire Gelu_for_else_Gelu_for_else_mux1h_3_nl;
  wire[21:0] Gelu_for_else_Gelu_for_else_mux1h_35_nl;
  wire Gelu_for_else_or_12_nl;
  wire[4:0] Gelu_for_else_Gelu_for_else_mux1h_19_nl;
  wire Gelu_for_else_Gelu_for_else_mux1h_51_nl;
  wire[2:0] Gelu_for_else_Gelu_for_else_mux1h_67_nl;
  wire Gelu_for_else_Gelu_for_else_mux1h_2_nl;
  wire[21:0] Gelu_for_else_Gelu_for_else_mux1h_34_nl;
  wire Gelu_for_else_or_13_nl;
  wire[4:0] Gelu_for_else_Gelu_for_else_mux1h_18_nl;
  wire Gelu_for_else_Gelu_for_else_mux1h_50_nl;
  wire[2:0] Gelu_for_else_Gelu_for_else_mux1h_66_nl;
  wire Gelu_for_else_Gelu_for_else_mux1h_1_nl;
  wire[21:0] Gelu_for_else_Gelu_for_else_mux1h_33_nl;
  wire Gelu_for_else_or_14_nl;
  wire[4:0] Gelu_for_else_Gelu_for_else_mux1h_17_nl;
  wire Gelu_for_else_Gelu_for_else_mux1h_49_nl;
  wire[2:0] Gelu_for_else_Gelu_for_else_mux1h_65_nl;
  wire Gelu_for_else_Gelu_for_else_mux1h_nl;
  wire[21:0] Gelu_for_else_Gelu_for_else_mux1h_32_nl;
  wire Gelu_for_else_or_15_nl;
  wire[4:0] Gelu_for_else_Gelu_for_else_mux1h_16_nl;
  wire Gelu_for_else_Gelu_for_else_mux1h_48_nl;
  wire[2:0] Gelu_for_else_Gelu_for_else_mux1h_64_nl;
  wire[4:0] ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_and_1_nl;
  wire mux_101_nl;
  wire nor_221_nl;
  wire or_356_nl;
  wire mux_114_nl;
  wire nor_224_nl;
  wire or_870_nl;
  wire or_869_nl;
  wire mux_332_nl;
  wire nand_22_nl;
  wire or_875_nl;
  wire or_874_nl;
  wire mux_342_nl;
  wire nand_24_nl;
  wire or_880_nl;
  wire or_879_nl;
  wire mux_352_nl;
  wire nand_26_nl;
  wire or_885_nl;
  wire or_884_nl;
  wire mux_362_nl;
  wire nand_28_nl;
  wire or_890_nl;
  wire or_889_nl;
  wire mux_372_nl;
  wire nand_30_nl;
  wire or_895_nl;
  wire or_894_nl;
  wire mux_382_nl;
  wire nand_32_nl;
  wire or_900_nl;
  wire or_899_nl;
  wire mux_392_nl;
  wire nand_34_nl;
  wire or_905_nl;
  wire or_904_nl;
  wire mux_402_nl;
  wire nand_36_nl;
  wire mux_428_nl;
  wire mux_434_nl;
  wire nand_252_nl;
  wire nand_39_nl;
  wire mux_435_nl;
  wire mux_446_nl;
  wire nor_451_nl;
  wire mux_1474_nl;
  wire nor_1650_nl;
  wire or_3343_nl;
  wire[25:0] Silu_for_10_else_else_else_if_acc_nl;
  wire[26:0] nl_Silu_for_10_else_else_else_if_acc_nl;
  wire[25:0] Silu_for_11_else_else_else_if_acc_nl;
  wire[26:0] nl_Silu_for_11_else_else_else_if_acc_nl;
  wire[21:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_122_nl;
  wire[25:0] Silu_for_12_else_else_else_if_acc_nl;
  wire[26:0] nl_Silu_for_12_else_else_else_if_acc_nl;
  wire[21:0] and_1777_nl;
  wire[21:0] mux1h_11_nl;
  wire not_2658_nl;
  wire[25:0] Silu_for_13_else_else_else_if_acc_nl;
  wire[26:0] nl_Silu_for_13_else_else_else_if_acc_nl;
  wire[21:0] and_1782_nl;
  wire[21:0] mux1h_12_nl;
  wire and_1442_nl;
  wire not_2660_nl;
  wire[25:0] Silu_for_14_else_else_else_if_acc_nl;
  wire[26:0] nl_Silu_for_14_else_else_else_if_acc_nl;
  wire[21:0] and_1786_nl;
  wire[21:0] mux1h_13_nl;
  wire and_1445_nl;
  wire not_2662_nl;
  wire[25:0] Silu_for_15_else_else_else_if_acc_nl;
  wire[26:0] nl_Silu_for_15_else_else_else_if_acc_nl;
  wire[21:0] and_1790_nl;
  wire[21:0] mux1h_14_nl;
  wire and_1448_nl;
  wire not_2664_nl;
  wire[25:0] Silu_for_16_else_else_else_if_acc_nl;
  wire[26:0] nl_Silu_for_16_else_else_else_if_acc_nl;
  wire[21:0] and_1794_nl;
  wire[21:0] mux1h_15_nl;
  wire and_1450_nl;
  wire not_2666_nl;
  wire mux_459_nl;
  wire nor_471_nl;
  wire nor_472_nl;
  wire mux_1050_nl;
  wire or_2499_nl;
  wire mux_1178_nl;
  wire or_2739_nl;
  wire mux_1249_nl;
  wire mux_1248_nl;
  wire mux_1244_nl;
  wire mux_1243_nl;
  wire mux_1239_nl;
  wire mux_1238_nl;
  wire mux_1234_nl;
  wire mux_1233_nl;
  wire mux_1229_nl;
  wire mux_1228_nl;
  wire mux_1224_nl;
  wire mux_1223_nl;
  wire mux_1219_nl;
  wire mux_1218_nl;
  wire mux_1214_nl;
  wire mux_1213_nl;
  wire mux_1209_nl;
  wire mux_1205_nl;
  wire mux_1201_nl;
  wire mux_1197_nl;
  wire mux_1193_nl;
  wire mux_1189_nl;
  wire mux_1185_nl;
  wire mux_1181_nl;
  wire mux_1177_nl;
  wire mux_1176_nl;
  wire mux_1173_nl;
  wire mux_1172_nl;
  wire mux_1169_nl;
  wire mux_1168_nl;
  wire mux_1165_nl;
  wire mux_1164_nl;
  wire mux_1161_nl;
  wire mux_1160_nl;
  wire mux_1157_nl;
  wire mux_1156_nl;
  wire mux_1153_nl;
  wire mux_1152_nl;
  wire mux_1149_nl;
  wire mux_1148_nl;
  wire mux_1145_nl;
  wire mux_1142_nl;
  wire mux_1139_nl;
  wire mux_1136_nl;
  wire mux_1133_nl;
  wire mux_1130_nl;
  wire mux_1127_nl;
  wire mux_1124_nl;
  wire mux_1121_nl;
  wire mux_1120_nl;
  wire mux_1116_nl;
  wire mux_1115_nl;
  wire mux_1111_nl;
  wire mux_1110_nl;
  wire mux_1106_nl;
  wire mux_1105_nl;
  wire mux_1101_nl;
  wire mux_1100_nl;
  wire mux_1096_nl;
  wire mux_1095_nl;
  wire mux_1091_nl;
  wire mux_1090_nl;
  wire mux_1086_nl;
  wire mux_1085_nl;
  wire mux_1081_nl;
  wire mux_1077_nl;
  wire mux_1073_nl;
  wire mux_1069_nl;
  wire mux_1065_nl;
  wire mux_1061_nl;
  wire mux_1057_nl;
  wire mux_1053_nl;
  wire mux_1049_nl;
  wire mux_1048_nl;
  wire mux_757_nl;
  wire mux_732_nl;
  wire mux_731_nl;
  wire nand_532_nl;
  wire mux_1045_nl;
  wire mux_1044_nl;
  wire mux_755_nl;
  wire mux_730_nl;
  wire or_1838_nl;
  wire mux_1025_nl;
  wire mux_1024_nl;
  wire mux_1021_nl;
  wire mux_1020_nl;
  wire mux_742_nl;
  wire mux_741_nl;
  wire nand_538_nl;
  wire mux_1017_nl;
  wire mux_769_nl;
  wire mux_729_nl;
  wire mux_728_nl;
  wire nand_530_nl;
  wire mux_1014_nl;
  wire mux_767_nl;
  wire and_2387_nl;
  wire mux_745_nl;
  wire mux_744_nl;
  wire mux_743_nl;
  wire and_1878_nl;
  wire mux_1011_nl;
  wire mux_765_nl;
  wire mux_740_nl;
  wire mux_739_nl;
  wire nand_537_nl;
  wire mux_1008_nl;
  wire mux_763_nl;
  wire nor_511_nl;
  wire mux_738_nl;
  wire mux_737_nl;
  wire nand_536_nl;
  wire mux_1005_nl;
  wire mux_761_nl;
  wire mux_736_nl;
  wire mux_735_nl;
  wire nand_535_nl;
  wire mux_1002_nl;
  wire mux_759_nl;
  wire nor_506_nl;
  wire mux_734_nl;
  wire mux_733_nl;
  wire nand_534_nl;
  wire mux_447_nl;
  wire or_943_nl;
  wire mux_1041_nl;
  wire mux_1040_nl;
  wire mux_753_nl;
  wire mux_1494_nl;
  wire mux_1493_nl;
  wire and_2822_nl;
  wire mux_1492_nl;
  wire mux_1491_nl;
  wire or_3389_nl;
  wire mux_1037_nl;
  wire mux_1036_nl;
  wire mux_751_nl;
  wire mux_1490_nl;
  wire mux_1489_nl;
  wire nor_1665_nl;
  wire mux_1488_nl;
  wire mux_1487_nl;
  wire or_3380_nl;
  wire mux_1033_nl;
  wire mux_1032_nl;
  wire mux_749_nl;
  wire mux_1486_nl;
  wire mux_1485_nl;
  wire nor_1661_nl;
  wire mux_1484_nl;
  wire mux_1483_nl;
  wire or_3370_nl;
  wire mux_1029_nl;
  wire mux_1028_nl;
  wire mux_747_nl;
  wire mux_1482_nl;
  wire mux_1481_nl;
  wire nor_1657_nl;
  wire mux_1480_nl;
  wire mux_1479_nl;
  wire or_3360_nl;
  wire mux_590_nl;
  wire and_2329_nl;
  wire mux_999_nl;
  wire mux_589_nl;
  wire mux_588_nl;
  wire nor_1404_nl;
  wire mux_1478_nl;
  wire mux_1477_nl;
  wire nor_1653_nl;
  wire mux_1476_nl;
  wire mux_1475_nl;
  wire or_3350_nl;
  wire mux_628_nl;
  wire mux_627_nl;
  wire mux_626_nl;
  wire mux_625_nl;
  wire mux_624_nl;
  wire mux_623_nl;
  wire mux_996_nl;
  wire mux_454_nl;
  wire mux_453_nl;
  wire or_1429_nl;
  wire mux_452_nl;
  wire or_1428_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_6_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_304_nl;
  wire and_1711_nl;
  wire mux1h_nl;
  wire[2:0] and_3505_nl;
  wire[2:0] mux1h_16_nl;
  wire not_8904_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_69_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_338_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_104_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_336_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_97_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_334_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_90_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_332_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_83_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_330_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_76_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_328_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_12_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_326_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_62_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_324_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_54_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_322_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_47_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_320_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_40_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_318_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_33_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_316_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_26_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_314_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_19_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_312_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_111_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_310_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_5_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_308_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_67_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_306_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_102_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_305_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_95_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_307_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_88_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_309_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_81_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_311_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_74_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_313_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_10_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_315_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_60_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_317_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_52_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_319_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_45_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_321_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_38_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_323_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_31_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_325_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_24_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_327_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_17_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_329_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_109_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_331_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_3_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_333_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_66_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_335_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_101_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_337_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_94_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_339_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_87_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_340_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_80_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_341_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_73_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_342_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_11_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_343_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_59_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_344_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_53_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_345_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_46_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_346_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_39_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_347_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_32_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_348_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_25_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_349_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_18_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_350_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_108_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_351_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_4_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_352_nl;
  wire nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_68_nl;
  wire[2:0] nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_353_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_9_nl;
  wire[2:0] ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_191_nl;
  wire not_8895_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_14_nl;
  wire[2:0] ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_190_nl;
  wire not_8894_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_19_nl;
  wire[2:0] ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_189_nl;
  wire not_8893_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_24_nl;
  wire[2:0] ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_188_nl;
  wire not_8892_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_29_nl;
  wire[2:0] ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_187_nl;
  wire not_8891_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_34_nl;
  wire[2:0] ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_198_nl;
  wire not_8903_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_39_nl;
  wire[2:0] ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_197_nl;
  wire not_8902_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_44_nl;
  wire[2:0] ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_196_nl;
  wire not_8901_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_49_nl;
  wire[2:0] ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_195_nl;
  wire not_8900_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_54_nl;
  wire[2:0] ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_194_nl;
  wire not_8899_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_59_nl;
  wire[2:0] ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_193_nl;
  wire not_8898_nl;
  wire ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_64_nl;
  wire[2:0] ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_192_nl;
  wire not_8897_nl;
  wire Silu_for_else_Silu_for_else_mux1h_23_nl;
  wire[2:0] Silu_for_else_Silu_for_else_mux1h_49_nl;
  wire Silu_for_else_Silu_for_else_mux1h_22_nl;
  wire[2:0] Silu_for_else_Silu_for_else_mux1h_51_nl;
  wire Silu_for_else_Silu_for_else_mux1h_21_nl;
  wire[2:0] Silu_for_else_Silu_for_else_mux1h_53_nl;
  wire Silu_for_else_Silu_for_else_mux1h_20_nl;
  wire[2:0] Silu_for_else_Silu_for_else_mux1h_55_nl;
  wire Silu_for_else_Silu_for_else_mux1h_19_nl;
  wire[2:0] Silu_for_else_Silu_for_else_mux1h_57_nl;
  wire Silu_for_else_Silu_for_else_mux1h_18_nl;
  wire[2:0] Silu_for_else_Silu_for_else_mux1h_59_nl;
  wire Silu_for_else_Silu_for_else_mux1h_17_nl;
  wire[2:0] Silu_for_else_Silu_for_else_mux1h_61_nl;
  wire Silu_for_else_Silu_for_else_mux1h_16_nl;
  wire[2:0] Silu_for_else_Silu_for_else_mux1h_63_nl;
  wire ActUnit_PushOutput_if_for_i_mux_nl;
  wire[2:0] ActUnit_PushOutput_if_for_i_mux_1_nl;
  wire not_8896_nl;
  wire Silu_for_else_Silu_for_else_mux1h_31_nl;
  wire[2:0] Silu_for_else_Silu_for_else_mux1h_65_nl;
  wire Silu_for_else_Silu_for_else_mux1h_30_nl;
  wire[2:0] Silu_for_else_Silu_for_else_mux1h_67_nl;
  wire Silu_for_else_Silu_for_else_mux1h_29_nl;
  wire[2:0] Silu_for_else_Silu_for_else_mux1h_69_nl;
  wire Silu_for_else_Silu_for_else_mux1h_28_nl;
  wire[2:0] Silu_for_else_Silu_for_else_mux1h_71_nl;
  wire Silu_for_else_Silu_for_else_mux1h_27_nl;
  wire[2:0] Silu_for_else_Silu_for_else_mux1h_73_nl;
  wire Silu_for_else_Silu_for_else_mux1h_26_nl;
  wire[2:0] Silu_for_else_Silu_for_else_mux1h_75_nl;
  wire Silu_for_else_Silu_for_else_mux1h_25_nl;
  wire[2:0] Silu_for_else_Silu_for_else_mux1h_77_nl;
  wire Silu_for_else_Silu_for_else_mux1h_24_nl;
  wire[2:0] Silu_for_else_Silu_for_else_mux1h_79_nl;
  wire[3:0] Silu_for_else_else_else_else_if_mux_nl;

  // Interconnect Declarations for Component Instantiations 
  wire[1:0] mux_535_nl;
  wire[2:0] mux_536_nl;
  wire[1:0] mux_537_nl;
  wire [24:0] nl_Gelu_for_1_else_else_else_if_mul_cmp_a;
  assign mux_535_nl = MUX_v_2_2_2(2'b10, 2'b01, operator_32_8_true_AC_TRN_AC_WRAP_6_less_15_tmp);
  assign mux_536_nl = MUX_v_3_2_2(3'b100, 3'b011, operator_32_8_true_AC_TRN_AC_WRAP_6_less_15_tmp);
  assign mux_537_nl = MUX_v_2_2_2(2'b01, 2'b10, operator_32_8_true_AC_TRN_AC_WRAP_6_less_15_tmp);
  assign nl_Gelu_for_1_else_else_else_if_mul_cmp_a = {mux_15_rmff , 2'b01 , mux_535_nl
      , 1'b0 , (signext_4_3(mux_536_nl)) , 3'b110 , mux_537_nl , 1'b1 , ({{1{mux_15_rmff[2]}},
      mux_15_rmff}) , 3'b001};
  wire Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_nl;
  wire [25:0] nl_Gelu_for_1_else_else_else_if_mul_cmp_b;
  assign Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_nl = reg_ActUnit_RunInst_case_15_nv_scvector_cctor_data_0_ftd_rsp_0
      & operator_32_8_true_AC_TRN_AC_WRAP_6_less_15_tmp;
  assign nl_Gelu_for_1_else_else_else_if_mul_cmp_b = {Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_nl
      , reg_ActUnit_RunInst_case_15_nv_scvector_cctor_data_0_ftd_rsp_1 , reg_ActUnit_RunInst_case_15_nv_scvector_cctor_data_0_ftd_1};
  wire[1:0] mux_531_nl;
  wire[2:0] mux_532_nl;
  wire[1:0] mux_533_nl;
  wire [24:0] nl_Gelu_for_1_else_else_else_if_mul_cmp_1_a;
  assign mux_531_nl = MUX_v_2_2_2(2'b10, 2'b01, operator_32_8_true_AC_TRN_AC_WRAP_6_less_tmp);
  assign mux_532_nl = MUX_v_3_2_2(3'b100, 3'b011, operator_32_8_true_AC_TRN_AC_WRAP_6_less_tmp);
  assign mux_533_nl = MUX_v_2_2_2(2'b01, 2'b10, operator_32_8_true_AC_TRN_AC_WRAP_6_less_tmp);
  assign nl_Gelu_for_1_else_else_else_if_mul_cmp_1_a = {mux_14_rmff , 2'b01 , mux_531_nl
      , 1'b0 , (signext_4_3(mux_532_nl)) , 3'b110 , mux_533_nl , 1'b1 , ({{1{mux_14_rmff[2]}},
      mux_14_rmff}) , 3'b001};
  wire Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_1_nl;
  wire [25:0] nl_Gelu_for_1_else_else_else_if_mul_cmp_1_b;
  assign Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_1_nl = reg_nv_scvector_cctor_nv_scvector_6_for_16_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      & operator_32_8_true_AC_TRN_AC_WRAP_6_less_tmp;
  assign nl_Gelu_for_1_else_else_else_if_mul_cmp_1_b = {Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_1_nl
      , reg_nv_scvector_cctor_nv_scvector_6_for_16_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_16_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1};
  wire[1:0] mux_527_nl;
  wire[2:0] mux_528_nl;
  wire[1:0] mux_529_nl;
  wire [24:0] nl_Gelu_for_1_else_else_else_if_mul_cmp_2_a;
  assign mux_527_nl = MUX_v_2_2_2(2'b10, 2'b01, operator_32_8_true_AC_TRN_AC_WRAP_6_less_1_tmp);
  assign mux_528_nl = MUX_v_3_2_2(3'b100, 3'b011, operator_32_8_true_AC_TRN_AC_WRAP_6_less_1_tmp);
  assign mux_529_nl = MUX_v_2_2_2(2'b01, 2'b10, operator_32_8_true_AC_TRN_AC_WRAP_6_less_1_tmp);
  assign nl_Gelu_for_1_else_else_else_if_mul_cmp_2_a = {mux_13_rmff , 2'b01 , mux_527_nl
      , 1'b0 , (signext_4_3(mux_528_nl)) , 3'b110 , mux_529_nl , 1'b1 , ({{1{mux_13_rmff[2]}},
      mux_13_rmff}) , 3'b001};
  wire Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_2_nl;
  wire [25:0] nl_Gelu_for_1_else_else_else_if_mul_cmp_2_b;
  assign Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_2_nl = reg_nv_scvector_cctor_nv_scvector_6_for_15_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      & operator_32_8_true_AC_TRN_AC_WRAP_6_less_1_tmp;
  assign nl_Gelu_for_1_else_else_else_if_mul_cmp_2_b = {Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_2_nl
      , reg_nv_scvector_cctor_nv_scvector_6_for_15_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_15_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1};
  wire[1:0] mux_523_nl;
  wire[2:0] mux_524_nl;
  wire[1:0] mux_525_nl;
  wire [24:0] nl_Gelu_for_1_else_else_else_if_mul_cmp_3_a;
  assign mux_523_nl = MUX_v_2_2_2(2'b10, 2'b01, operator_32_8_true_AC_TRN_AC_WRAP_6_less_2_tmp);
  assign mux_524_nl = MUX_v_3_2_2(3'b100, 3'b011, operator_32_8_true_AC_TRN_AC_WRAP_6_less_2_tmp);
  assign mux_525_nl = MUX_v_2_2_2(2'b01, 2'b10, operator_32_8_true_AC_TRN_AC_WRAP_6_less_2_tmp);
  assign nl_Gelu_for_1_else_else_else_if_mul_cmp_3_a = {mux_12_rmff , 2'b01 , mux_523_nl
      , 1'b0 , (signext_4_3(mux_524_nl)) , 3'b110 , mux_525_nl , 1'b1 , ({{1{mux_12_rmff[2]}},
      mux_12_rmff}) , 3'b001};
  wire Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_3_nl;
  wire [25:0] nl_Gelu_for_1_else_else_else_if_mul_cmp_3_b;
  assign Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_3_nl = reg_nv_scvector_cctor_nv_scvector_6_for_14_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      & operator_32_8_true_AC_TRN_AC_WRAP_6_less_2_tmp;
  assign nl_Gelu_for_1_else_else_else_if_mul_cmp_3_b = {Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_3_nl
      , reg_nv_scvector_cctor_nv_scvector_6_for_14_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_14_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1};
  wire[1:0] mux_519_nl;
  wire[2:0] mux_520_nl;
  wire[1:0] mux_521_nl;
  wire [24:0] nl_Gelu_for_1_else_else_else_if_mul_cmp_4_a;
  assign mux_519_nl = MUX_v_2_2_2(2'b10, 2'b01, operator_32_8_true_AC_TRN_AC_WRAP_6_less_3_tmp);
  assign mux_520_nl = MUX_v_3_2_2(3'b100, 3'b011, operator_32_8_true_AC_TRN_AC_WRAP_6_less_3_tmp);
  assign mux_521_nl = MUX_v_2_2_2(2'b01, 2'b10, operator_32_8_true_AC_TRN_AC_WRAP_6_less_3_tmp);
  assign nl_Gelu_for_1_else_else_else_if_mul_cmp_4_a = {mux_11_rmff , 2'b01 , mux_519_nl
      , 1'b0 , (signext_4_3(mux_520_nl)) , 3'b110 , mux_521_nl , 1'b1 , ({{1{mux_11_rmff[2]}},
      mux_11_rmff}) , 3'b001};
  wire Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_4_nl;
  wire [25:0] nl_Gelu_for_1_else_else_else_if_mul_cmp_4_b;
  assign Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_4_nl = reg_nv_scvector_cctor_nv_scvector_6_for_13_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      & operator_32_8_true_AC_TRN_AC_WRAP_6_less_3_tmp;
  assign nl_Gelu_for_1_else_else_else_if_mul_cmp_4_b = {Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_4_nl
      , reg_nv_scvector_cctor_nv_scvector_6_for_13_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_13_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1};
  wire[1:0] mux_515_nl;
  wire[2:0] mux_516_nl;
  wire[1:0] mux_517_nl;
  wire [24:0] nl_Gelu_for_1_else_else_else_if_mul_cmp_5_a;
  assign mux_515_nl = MUX_v_2_2_2(2'b10, 2'b01, operator_32_8_true_AC_TRN_AC_WRAP_6_less_4_tmp);
  assign mux_516_nl = MUX_v_3_2_2(3'b100, 3'b011, operator_32_8_true_AC_TRN_AC_WRAP_6_less_4_tmp);
  assign mux_517_nl = MUX_v_2_2_2(2'b01, 2'b10, operator_32_8_true_AC_TRN_AC_WRAP_6_less_4_tmp);
  assign nl_Gelu_for_1_else_else_else_if_mul_cmp_5_a = {mux_10_rmff , 2'b01 , mux_515_nl
      , 1'b0 , (signext_4_3(mux_516_nl)) , 3'b110 , mux_517_nl , 1'b1 , ({{1{mux_10_rmff[2]}},
      mux_10_rmff}) , 3'b001};
  wire Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_5_nl;
  wire [25:0] nl_Gelu_for_1_else_else_else_if_mul_cmp_5_b;
  assign Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_5_nl = reg_nv_scvector_cctor_nv_scvector_6_for_12_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      & operator_32_8_true_AC_TRN_AC_WRAP_6_less_4_tmp;
  assign nl_Gelu_for_1_else_else_else_if_mul_cmp_5_b = {Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_5_nl
      , reg_nv_scvector_cctor_nv_scvector_6_for_12_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_12_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1};
  wire[1:0] mux_511_nl;
  wire[2:0] mux_512_nl;
  wire[1:0] mux_513_nl;
  wire [24:0] nl_Gelu_for_1_else_else_else_if_mul_cmp_6_a;
  assign mux_511_nl = MUX_v_2_2_2(2'b10, 2'b01, operator_32_8_true_AC_TRN_AC_WRAP_6_less_5_tmp);
  assign mux_512_nl = MUX_v_3_2_2(3'b100, 3'b011, operator_32_8_true_AC_TRN_AC_WRAP_6_less_5_tmp);
  assign mux_513_nl = MUX_v_2_2_2(2'b01, 2'b10, operator_32_8_true_AC_TRN_AC_WRAP_6_less_5_tmp);
  assign nl_Gelu_for_1_else_else_else_if_mul_cmp_6_a = {mux_9_rmff , 2'b01 , mux_511_nl
      , 1'b0 , (signext_4_3(mux_512_nl)) , 3'b110 , mux_513_nl , 1'b1 , ({{1{mux_9_rmff[2]}},
      mux_9_rmff}) , 3'b001};
  wire Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_6_nl;
  wire [25:0] nl_Gelu_for_1_else_else_else_if_mul_cmp_6_b;
  assign Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_6_nl = reg_nv_scvector_cctor_nv_scvector_6_for_11_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      & operator_32_8_true_AC_TRN_AC_WRAP_6_less_5_tmp;
  assign nl_Gelu_for_1_else_else_else_if_mul_cmp_6_b = {Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_6_nl
      , reg_nv_scvector_cctor_nv_scvector_6_for_11_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_11_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1};
  wire[1:0] mux_507_nl;
  wire[2:0] mux_508_nl;
  wire[1:0] mux_509_nl;
  wire [24:0] nl_Gelu_for_1_else_else_else_if_mul_cmp_7_a;
  assign mux_507_nl = MUX_v_2_2_2(2'b10, 2'b01, operator_32_8_true_AC_TRN_AC_WRAP_6_less_6_tmp);
  assign mux_508_nl = MUX_v_3_2_2(3'b100, 3'b011, operator_32_8_true_AC_TRN_AC_WRAP_6_less_6_tmp);
  assign mux_509_nl = MUX_v_2_2_2(2'b01, 2'b10, operator_32_8_true_AC_TRN_AC_WRAP_6_less_6_tmp);
  assign nl_Gelu_for_1_else_else_else_if_mul_cmp_7_a = {mux_8_rmff , 2'b01 , mux_507_nl
      , 1'b0 , (signext_4_3(mux_508_nl)) , 3'b110 , mux_509_nl , 1'b1 , ({{1{mux_8_rmff[2]}},
      mux_8_rmff}) , 3'b001};
  wire Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_7_nl;
  wire [25:0] nl_Gelu_for_1_else_else_else_if_mul_cmp_7_b;
  assign Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_7_nl = reg_nv_scvector_cctor_nv_scvector_6_for_10_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      & operator_32_8_true_AC_TRN_AC_WRAP_6_less_6_tmp;
  assign nl_Gelu_for_1_else_else_else_if_mul_cmp_7_b = {Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_7_nl
      , reg_nv_scvector_cctor_nv_scvector_6_for_10_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_10_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1};
  wire[1:0] mux_503_nl;
  wire[2:0] mux_504_nl;
  wire[1:0] mux_505_nl;
  wire [24:0] nl_Gelu_for_1_else_else_else_if_mul_cmp_8_a;
  assign mux_503_nl = MUX_v_2_2_2(2'b10, 2'b01, operator_32_8_true_AC_TRN_AC_WRAP_6_less_7_tmp);
  assign mux_504_nl = MUX_v_3_2_2(3'b100, 3'b011, operator_32_8_true_AC_TRN_AC_WRAP_6_less_7_tmp);
  assign mux_505_nl = MUX_v_2_2_2(2'b01, 2'b10, operator_32_8_true_AC_TRN_AC_WRAP_6_less_7_tmp);
  assign nl_Gelu_for_1_else_else_else_if_mul_cmp_8_a = {mux_7_rmff , 2'b01 , mux_503_nl
      , 1'b0 , (signext_4_3(mux_504_nl)) , 3'b110 , mux_505_nl , 1'b1 , ({{1{mux_7_rmff[2]}},
      mux_7_rmff}) , 3'b001};
  wire Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_8_nl;
  wire [25:0] nl_Gelu_for_1_else_else_else_if_mul_cmp_8_b;
  assign Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_8_nl = reg_nv_scvector_cctor_nv_scvector_6_for_9_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      & operator_32_8_true_AC_TRN_AC_WRAP_6_less_7_tmp;
  assign nl_Gelu_for_1_else_else_else_if_mul_cmp_8_b = {Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_8_nl
      , reg_nv_scvector_cctor_nv_scvector_6_for_9_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_9_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1};
  wire[1:0] mux_499_nl;
  wire[2:0] mux_500_nl;
  wire[1:0] mux_501_nl;
  wire [24:0] nl_Gelu_for_1_else_else_else_if_mul_cmp_9_a;
  assign mux_499_nl = MUX_v_2_2_2(2'b10, 2'b01, operator_32_8_true_AC_TRN_AC_WRAP_6_less_8_tmp);
  assign mux_500_nl = MUX_v_3_2_2(3'b100, 3'b011, operator_32_8_true_AC_TRN_AC_WRAP_6_less_8_tmp);
  assign mux_501_nl = MUX_v_2_2_2(2'b01, 2'b10, operator_32_8_true_AC_TRN_AC_WRAP_6_less_8_tmp);
  assign nl_Gelu_for_1_else_else_else_if_mul_cmp_9_a = {mux_6_rmff , 2'b01 , mux_499_nl
      , 1'b0 , (signext_4_3(mux_500_nl)) , 3'b110 , mux_501_nl , 1'b1 , ({{1{mux_6_rmff[2]}},
      mux_6_rmff}) , 3'b001};
  wire Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_9_nl;
  wire [25:0] nl_Gelu_for_1_else_else_else_if_mul_cmp_9_b;
  assign Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_9_nl = reg_nv_scvector_cctor_nv_scvector_6_for_8_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      & operator_32_8_true_AC_TRN_AC_WRAP_6_less_8_tmp;
  assign nl_Gelu_for_1_else_else_else_if_mul_cmp_9_b = {Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_9_nl
      , reg_nv_scvector_cctor_nv_scvector_6_for_8_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_8_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1};
  wire[1:0] mux_495_nl;
  wire[2:0] mux_496_nl;
  wire[1:0] mux_497_nl;
  wire [24:0] nl_Gelu_for_1_else_else_else_if_mul_cmp_10_a;
  assign mux_495_nl = MUX_v_2_2_2(2'b10, 2'b01, operator_32_8_true_AC_TRN_AC_WRAP_6_less_9_tmp);
  assign mux_496_nl = MUX_v_3_2_2(3'b100, 3'b011, operator_32_8_true_AC_TRN_AC_WRAP_6_less_9_tmp);
  assign mux_497_nl = MUX_v_2_2_2(2'b01, 2'b10, operator_32_8_true_AC_TRN_AC_WRAP_6_less_9_tmp);
  assign nl_Gelu_for_1_else_else_else_if_mul_cmp_10_a = {mux_5_rmff , 2'b01 , mux_495_nl
      , 1'b0 , (signext_4_3(mux_496_nl)) , 3'b110 , mux_497_nl , 1'b1 , ({{1{mux_5_rmff[2]}},
      mux_5_rmff}) , 3'b001};
  wire Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_10_nl;
  wire [25:0] nl_Gelu_for_1_else_else_else_if_mul_cmp_10_b;
  assign Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_10_nl = reg_nv_scvector_cctor_nv_scvector_6_for_7_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      & operator_32_8_true_AC_TRN_AC_WRAP_6_less_9_tmp;
  assign nl_Gelu_for_1_else_else_else_if_mul_cmp_10_b = {Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_10_nl
      , reg_nv_scvector_cctor_nv_scvector_6_for_7_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_7_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1};
  wire[1:0] mux_491_nl;
  wire[2:0] mux_492_nl;
  wire[1:0] mux_493_nl;
  wire [24:0] nl_Gelu_for_1_else_else_else_if_mul_cmp_11_a;
  assign mux_491_nl = MUX_v_2_2_2(2'b10, 2'b01, operator_32_8_true_AC_TRN_AC_WRAP_6_less_10_tmp);
  assign mux_492_nl = MUX_v_3_2_2(3'b100, 3'b011, operator_32_8_true_AC_TRN_AC_WRAP_6_less_10_tmp);
  assign mux_493_nl = MUX_v_2_2_2(2'b01, 2'b10, operator_32_8_true_AC_TRN_AC_WRAP_6_less_10_tmp);
  assign nl_Gelu_for_1_else_else_else_if_mul_cmp_11_a = {mux_4_rmff , 2'b01 , mux_491_nl
      , 1'b0 , (signext_4_3(mux_492_nl)) , 3'b110 , mux_493_nl , 1'b1 , ({{1{mux_4_rmff[2]}},
      mux_4_rmff}) , 3'b001};
  wire Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_11_nl;
  wire [25:0] nl_Gelu_for_1_else_else_else_if_mul_cmp_11_b;
  assign Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_11_nl = reg_nv_scvector_cctor_nv_scvector_6_for_6_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      & operator_32_8_true_AC_TRN_AC_WRAP_6_less_10_tmp;
  assign nl_Gelu_for_1_else_else_else_if_mul_cmp_11_b = {Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_11_nl
      , reg_nv_scvector_cctor_nv_scvector_6_for_6_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_6_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1};
  wire[1:0] mux_487_nl;
  wire[2:0] mux_488_nl;
  wire[1:0] mux_489_nl;
  wire [24:0] nl_Gelu_for_1_else_else_else_if_mul_cmp_12_a;
  assign mux_487_nl = MUX_v_2_2_2(2'b10, 2'b01, operator_32_8_true_AC_TRN_AC_WRAP_6_less_11_tmp);
  assign mux_488_nl = MUX_v_3_2_2(3'b100, 3'b011, operator_32_8_true_AC_TRN_AC_WRAP_6_less_11_tmp);
  assign mux_489_nl = MUX_v_2_2_2(2'b01, 2'b10, operator_32_8_true_AC_TRN_AC_WRAP_6_less_11_tmp);
  assign nl_Gelu_for_1_else_else_else_if_mul_cmp_12_a = {mux_3_rmff , 2'b01 , mux_487_nl
      , 1'b0 , (signext_4_3(mux_488_nl)) , 3'b110 , mux_489_nl , 1'b1 , ({{1{mux_3_rmff[2]}},
      mux_3_rmff}) , 3'b001};
  wire Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_12_nl;
  wire [25:0] nl_Gelu_for_1_else_else_else_if_mul_cmp_12_b;
  assign Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_12_nl = reg_nv_scvector_cctor_nv_scvector_6_for_5_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      & operator_32_8_true_AC_TRN_AC_WRAP_6_less_11_tmp;
  assign nl_Gelu_for_1_else_else_else_if_mul_cmp_12_b = {Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_12_nl
      , reg_nv_scvector_cctor_nv_scvector_6_for_5_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_5_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1};
  wire[1:0] mux_483_nl;
  wire[2:0] mux_484_nl;
  wire[1:0] mux_485_nl;
  wire [24:0] nl_Gelu_for_1_else_else_else_if_mul_cmp_13_a;
  assign mux_483_nl = MUX_v_2_2_2(2'b10, 2'b01, operator_32_8_true_AC_TRN_AC_WRAP_6_less_12_tmp);
  assign mux_484_nl = MUX_v_3_2_2(3'b100, 3'b011, operator_32_8_true_AC_TRN_AC_WRAP_6_less_12_tmp);
  assign mux_485_nl = MUX_v_2_2_2(2'b01, 2'b10, operator_32_8_true_AC_TRN_AC_WRAP_6_less_12_tmp);
  assign nl_Gelu_for_1_else_else_else_if_mul_cmp_13_a = {mux_2_rmff , 2'b01 , mux_483_nl
      , 1'b0 , (signext_4_3(mux_484_nl)) , 3'b110 , mux_485_nl , 1'b1 , ({{1{mux_2_rmff[2]}},
      mux_2_rmff}) , 3'b001};
  wire Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_13_nl;
  wire [25:0] nl_Gelu_for_1_else_else_else_if_mul_cmp_13_b;
  assign Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_13_nl = reg_nv_scvector_cctor_nv_scvector_6_for_4_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      & operator_32_8_true_AC_TRN_AC_WRAP_6_less_12_tmp;
  assign nl_Gelu_for_1_else_else_else_if_mul_cmp_13_b = {Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_13_nl
      , reg_nv_scvector_cctor_nv_scvector_6_for_4_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_4_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1};
  wire[1:0] mux_479_nl;
  wire[2:0] mux_480_nl;
  wire[1:0] mux_481_nl;
  wire [24:0] nl_Gelu_for_1_else_else_else_if_mul_cmp_14_a;
  assign mux_479_nl = MUX_v_2_2_2(2'b10, 2'b01, operator_32_8_true_AC_TRN_AC_WRAP_6_less_13_tmp);
  assign mux_480_nl = MUX_v_3_2_2(3'b100, 3'b011, operator_32_8_true_AC_TRN_AC_WRAP_6_less_13_tmp);
  assign mux_481_nl = MUX_v_2_2_2(2'b01, 2'b10, operator_32_8_true_AC_TRN_AC_WRAP_6_less_13_tmp);
  assign nl_Gelu_for_1_else_else_else_if_mul_cmp_14_a = {mux_1_rmff , 2'b01 , mux_479_nl
      , 1'b0 , (signext_4_3(mux_480_nl)) , 3'b110 , mux_481_nl , 1'b1 , ({{1{mux_1_rmff[2]}},
      mux_1_rmff}) , 3'b001};
  wire Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_14_nl;
  wire [25:0] nl_Gelu_for_1_else_else_else_if_mul_cmp_14_b;
  assign Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_14_nl = reg_nv_scvector_cctor_nv_scvector_6_for_3_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      & operator_32_8_true_AC_TRN_AC_WRAP_6_less_13_tmp;
  assign nl_Gelu_for_1_else_else_else_if_mul_cmp_14_b = {Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_14_nl
      , reg_nv_scvector_cctor_nv_scvector_6_for_3_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_3_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1};
  wire[1:0] mux_475_nl;
  wire[2:0] mux_476_nl;
  wire[1:0] mux_477_nl;
  wire [24:0] nl_Gelu_for_1_else_else_else_if_mul_cmp_15_a;
  assign mux_475_nl = MUX_v_2_2_2(2'b10, 2'b01, operator_32_8_true_AC_TRN_AC_WRAP_6_less_14_tmp);
  assign mux_476_nl = MUX_v_3_2_2(3'b100, 3'b011, operator_32_8_true_AC_TRN_AC_WRAP_6_less_14_tmp);
  assign mux_477_nl = MUX_v_2_2_2(2'b01, 2'b10, operator_32_8_true_AC_TRN_AC_WRAP_6_less_14_tmp);
  assign nl_Gelu_for_1_else_else_else_if_mul_cmp_15_a = {mux_rmff , 2'b01 , mux_475_nl
      , 1'b0 , (signext_4_3(mux_476_nl)) , 3'b110 , mux_477_nl , 1'b1 , ({{1{mux_rmff[2]}},
      mux_rmff}) , 3'b001};
  wire Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_15_nl;
  wire [25:0] nl_Gelu_for_1_else_else_else_if_mul_cmp_15_b;
  assign Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_15_nl = reg_nv_scvector_cctor_nv_scvector_6_for_2_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      & operator_32_8_true_AC_TRN_AC_WRAP_6_less_14_tmp;
  assign nl_Gelu_for_1_else_else_else_if_mul_cmp_15_b = {Gelu_for_else_else_else_if_Gelu_for_else_else_else_if_and_15_nl
      , reg_nv_scvector_cctor_nv_scvector_6_for_2_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_2_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1};
  wire [24:0] nl_Gelu_for_1_else_else_if_mul_cmp_b;
  assign nl_Gelu_for_1_else_else_if_mul_cmp_b = {reg_ActUnit_RunInst_case_15_nv_scvector_cctor_data_0_ftd_rsp_1
      , reg_ActUnit_RunInst_case_15_nv_scvector_cctor_data_0_ftd_1};
  wire [24:0] nl_Gelu_for_1_else_else_if_mul_cmp_1_b;
  assign nl_Gelu_for_1_else_else_if_mul_cmp_1_b = {reg_nv_scvector_cctor_nv_scvector_6_for_16_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_16_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1};
  wire [24:0] nl_Gelu_for_1_else_else_if_mul_cmp_2_b;
  assign nl_Gelu_for_1_else_else_if_mul_cmp_2_b = {reg_nv_scvector_cctor_nv_scvector_6_for_15_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_15_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1};
  wire [24:0] nl_Gelu_for_1_else_else_if_mul_cmp_3_b;
  assign nl_Gelu_for_1_else_else_if_mul_cmp_3_b = {reg_nv_scvector_cctor_nv_scvector_6_for_14_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_14_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1};
  wire [24:0] nl_Gelu_for_1_else_else_if_mul_cmp_4_b;
  assign nl_Gelu_for_1_else_else_if_mul_cmp_4_b = {reg_nv_scvector_cctor_nv_scvector_6_for_13_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_13_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1};
  wire [24:0] nl_Gelu_for_1_else_else_if_mul_cmp_5_b;
  assign nl_Gelu_for_1_else_else_if_mul_cmp_5_b = {reg_nv_scvector_cctor_nv_scvector_6_for_12_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_12_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1};
  wire [24:0] nl_Gelu_for_1_else_else_if_mul_cmp_6_b;
  assign nl_Gelu_for_1_else_else_if_mul_cmp_6_b = {reg_nv_scvector_cctor_nv_scvector_6_for_11_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_11_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1};
  wire [24:0] nl_Gelu_for_1_else_else_if_mul_cmp_7_b;
  assign nl_Gelu_for_1_else_else_if_mul_cmp_7_b = {reg_nv_scvector_cctor_nv_scvector_6_for_10_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_10_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1};
  wire [24:0] nl_Gelu_for_1_else_else_if_mul_cmp_8_b;
  assign nl_Gelu_for_1_else_else_if_mul_cmp_8_b = {reg_nv_scvector_cctor_nv_scvector_6_for_9_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_9_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1};
  wire [24:0] nl_Gelu_for_1_else_else_if_mul_cmp_9_b;
  assign nl_Gelu_for_1_else_else_if_mul_cmp_9_b = {reg_nv_scvector_cctor_nv_scvector_6_for_8_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_8_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1};
  wire [24:0] nl_Gelu_for_1_else_else_if_mul_cmp_10_b;
  assign nl_Gelu_for_1_else_else_if_mul_cmp_10_b = {reg_nv_scvector_cctor_nv_scvector_6_for_7_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_7_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1};
  wire [24:0] nl_Gelu_for_1_else_else_if_mul_cmp_11_b;
  assign nl_Gelu_for_1_else_else_if_mul_cmp_11_b = {reg_nv_scvector_cctor_nv_scvector_6_for_6_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_6_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1};
  wire [24:0] nl_Gelu_for_1_else_else_if_mul_cmp_12_b;
  assign nl_Gelu_for_1_else_else_if_mul_cmp_12_b = {reg_nv_scvector_cctor_nv_scvector_6_for_5_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_5_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1};
  wire [24:0] nl_Gelu_for_1_else_else_if_mul_cmp_13_b;
  assign nl_Gelu_for_1_else_else_if_mul_cmp_13_b = {reg_nv_scvector_cctor_nv_scvector_6_for_4_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_4_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1};
  wire [24:0] nl_Gelu_for_1_else_else_if_mul_cmp_14_b;
  assign nl_Gelu_for_1_else_else_if_mul_cmp_14_b = {reg_nv_scvector_cctor_nv_scvector_6_for_3_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_3_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1};
  wire [24:0] nl_Gelu_for_1_else_else_if_mul_cmp_15_b;
  assign nl_Gelu_for_1_else_else_if_mul_cmp_15_b = {reg_nv_scvector_cctor_nv_scvector_6_for_2_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_2_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1};
  wire [20:0] nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_a;
  assign nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_a = {Silu_for_else_if_Silu_for_else_if_or_itm
      , 20'b00110011001100110011};
  wire Silu_for_else_if_mux1h_23_nl;
  wire[2:0] Silu_for_else_if_mux1h_49_nl;
  wire[21:0] Silu_for_else_if_mux1h_41_nl;
  wire [26:0] nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_b;
  assign Silu_for_else_if_mux1h_23_nl = MUX1HOT_s_1_4_2(nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3,
      nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3,
      reg_nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0,
      reg_nv_scvector_cctor_nv_scvector_6_for_16_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0,
      {Silu_for_else_if_and_1_cse , Silu_for_else_if_and_2_cse , and_dcpl_852 , and_dcpl_855});
  assign Silu_for_else_if_mux1h_49_nl = MUX1HOT_v_3_4_2(nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0,
      nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0,
      reg_nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1,
      reg_nv_scvector_cctor_nv_scvector_6_for_16_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1,
      {Silu_for_else_if_and_1_cse , Silu_for_else_if_and_2_cse , and_dcpl_852 , and_dcpl_855});
  assign Silu_for_else_if_mux1h_41_nl = MUX1HOT_v_22_4_2(nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm,
      nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm,
      reg_nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1,
      reg_nv_scvector_cctor_nv_scvector_6_for_16_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1,
      {Silu_for_else_if_and_1_cse , Silu_for_else_if_and_2_cse , and_dcpl_852 , and_dcpl_855});
  assign nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_b = {1'b1 , Silu_for_else_if_mux1h_23_nl
      , Silu_for_else_if_mux1h_49_nl , Silu_for_else_if_mux1h_41_nl};
  wire [20:0] nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_1_a;
  assign nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_1_a = {Silu_for_else_if_Silu_for_else_if_or_itm
      , 20'b00110011001100110011};
  wire Silu_for_else_if_mux1h_20_nl;
  wire[2:0] Silu_for_else_if_mux1h_50_nl;
  wire[21:0] Silu_for_else_if_mux1h_42_nl;
  wire [26:0] nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_1_b;
  assign Silu_for_else_if_mux1h_20_nl = MUX1HOT_s_1_3_2(nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3,
      reg_nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0,
      reg_nv_scvector_cctor_nv_scvector_6_for_15_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0,
      {and_dcpl_847 , and_dcpl_852 , and_dcpl_855});
  assign Silu_for_else_if_mux1h_50_nl = MUX1HOT_v_3_3_2(nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0,
      reg_nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1,
      reg_nv_scvector_cctor_nv_scvector_6_for_15_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1,
      {and_dcpl_847 , and_dcpl_852 , and_dcpl_855});
  assign Silu_for_else_if_mux1h_42_nl = MUX1HOT_v_22_3_2(nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm,
      reg_nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1,
      reg_nv_scvector_cctor_nv_scvector_6_for_15_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1,
      {and_dcpl_847 , and_dcpl_852 , and_dcpl_855});
  assign nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_1_b = {1'b1 , Silu_for_else_if_mux1h_20_nl
      , Silu_for_else_if_mux1h_50_nl , Silu_for_else_if_mux1h_42_nl};
  wire [20:0] nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_2_a;
  assign nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_2_a = {Silu_for_else_if_Silu_for_else_if_or_itm
      , 20'b00110011001100110011};
  wire Silu_for_else_if_mux1h_17_nl;
  wire[2:0] Silu_for_else_if_mux1h_51_nl;
  wire[21:0] Silu_for_else_if_mux1h_43_nl;
  wire [26:0] nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_2_b;
  assign Silu_for_else_if_mux1h_17_nl = MUX1HOT_s_1_3_2(nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3,
      reg_nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0,
      reg_nv_scvector_cctor_nv_scvector_6_for_14_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0,
      {and_dcpl_847 , and_dcpl_852 , and_dcpl_855});
  assign Silu_for_else_if_mux1h_51_nl = MUX1HOT_v_3_3_2(nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0,
      reg_nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1,
      reg_nv_scvector_cctor_nv_scvector_6_for_14_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1,
      {and_dcpl_847 , and_dcpl_852 , and_dcpl_855});
  assign Silu_for_else_if_mux1h_43_nl = MUX1HOT_v_22_3_2(nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm,
      reg_nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1,
      reg_nv_scvector_cctor_nv_scvector_6_for_14_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1,
      {and_dcpl_847 , and_dcpl_852 , and_dcpl_855});
  assign nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_2_b = {1'b1 , Silu_for_else_if_mux1h_17_nl
      , Silu_for_else_if_mux1h_51_nl , Silu_for_else_if_mux1h_43_nl};
  wire [20:0] nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_3_a;
  assign nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_3_a = {Silu_for_else_if_Silu_for_else_if_or_itm
      , 20'b00110011001100110011};
  wire Silu_for_else_if_mux1h_14_nl;
  wire[2:0] Silu_for_else_if_mux1h_52_nl;
  wire[21:0] Silu_for_else_if_mux1h_44_nl;
  wire [26:0] nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_3_b;
  assign Silu_for_else_if_mux1h_14_nl = MUX1HOT_s_1_3_2(nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3,
      reg_nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0,
      reg_nv_scvector_cctor_nv_scvector_6_for_13_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0,
      {and_dcpl_847 , and_dcpl_852 , and_dcpl_855});
  assign Silu_for_else_if_mux1h_52_nl = MUX1HOT_v_3_3_2(nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0,
      reg_nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1,
      reg_nv_scvector_cctor_nv_scvector_6_for_13_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1,
      {and_dcpl_847 , and_dcpl_852 , and_dcpl_855});
  assign Silu_for_else_if_mux1h_44_nl = MUX1HOT_v_22_3_2(nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm,
      reg_nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1,
      reg_nv_scvector_cctor_nv_scvector_6_for_13_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1,
      {and_dcpl_847 , and_dcpl_852 , and_dcpl_855});
  assign nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_3_b = {1'b1 , Silu_for_else_if_mux1h_14_nl
      , Silu_for_else_if_mux1h_52_nl , Silu_for_else_if_mux1h_44_nl};
  wire [20:0] nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_4_a;
  assign nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_4_a = {Silu_for_else_if_Silu_for_else_if_or_itm
      , 20'b00110011001100110011};
  wire Silu_for_else_if_mux1h_11_nl;
  wire[2:0] Silu_for_else_if_mux1h_53_nl;
  wire[21:0] Silu_for_else_if_mux1h_45_nl;
  wire [26:0] nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_4_b;
  assign Silu_for_else_if_mux1h_11_nl = MUX1HOT_s_1_3_2(nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3,
      reg_nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0,
      reg_nv_scvector_cctor_nv_scvector_6_for_12_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0,
      {and_dcpl_847 , and_dcpl_852 , and_dcpl_855});
  assign Silu_for_else_if_mux1h_53_nl = MUX1HOT_v_3_3_2(nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0,
      reg_nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1,
      reg_nv_scvector_cctor_nv_scvector_6_for_12_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1,
      {and_dcpl_847 , and_dcpl_852 , and_dcpl_855});
  assign Silu_for_else_if_mux1h_45_nl = MUX1HOT_v_22_3_2(nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm,
      reg_nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1,
      reg_nv_scvector_cctor_nv_scvector_6_for_12_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1,
      {and_dcpl_847 , and_dcpl_852 , and_dcpl_855});
  assign nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_4_b = {1'b1 , Silu_for_else_if_mux1h_11_nl
      , Silu_for_else_if_mux1h_53_nl , Silu_for_else_if_mux1h_45_nl};
  wire [20:0] nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_5_a;
  assign nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_5_a = {Silu_for_else_if_Silu_for_else_if_or_itm
      , 20'b00110011001100110011};
  wire Silu_for_else_if_mux1h_8_nl;
  wire[2:0] Silu_for_else_if_mux1h_54_nl;
  wire[21:0] Silu_for_else_if_mux1h_46_nl;
  wire [26:0] nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_5_b;
  assign Silu_for_else_if_mux1h_8_nl = MUX1HOT_s_1_3_2(nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3,
      reg_nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0,
      reg_nv_scvector_cctor_nv_scvector_6_for_11_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0,
      {and_dcpl_847 , and_dcpl_852 , and_dcpl_855});
  assign Silu_for_else_if_mux1h_54_nl = MUX1HOT_v_3_3_2(nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0,
      reg_nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1,
      reg_nv_scvector_cctor_nv_scvector_6_for_11_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1,
      {and_dcpl_847 , and_dcpl_852 , and_dcpl_855});
  assign Silu_for_else_if_mux1h_46_nl = MUX1HOT_v_22_3_2(nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm,
      reg_nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1,
      reg_nv_scvector_cctor_nv_scvector_6_for_11_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1,
      {and_dcpl_847 , and_dcpl_852 , and_dcpl_855});
  assign nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_5_b = {1'b1 , Silu_for_else_if_mux1h_8_nl
      , Silu_for_else_if_mux1h_54_nl , Silu_for_else_if_mux1h_46_nl};
  wire [20:0] nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_6_a;
  assign nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_6_a = {Silu_for_else_if_Silu_for_else_if_or_itm
      , 20'b00110011001100110011};
  wire Silu_for_else_if_mux1h_5_nl;
  wire[2:0] Silu_for_else_if_mux1h_55_nl;
  wire[21:0] Silu_for_else_if_mux1h_47_nl;
  wire [26:0] nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_6_b;
  assign Silu_for_else_if_mux1h_5_nl = MUX1HOT_s_1_3_2(nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3,
      reg_nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0,
      reg_nv_scvector_cctor_nv_scvector_6_for_10_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0,
      {and_dcpl_847 , and_dcpl_852 , and_dcpl_855});
  assign Silu_for_else_if_mux1h_55_nl = MUX1HOT_v_3_3_2(nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0,
      reg_nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1,
      reg_nv_scvector_cctor_nv_scvector_6_for_10_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1,
      {and_dcpl_847 , and_dcpl_852 , and_dcpl_855});
  assign Silu_for_else_if_mux1h_47_nl = MUX1HOT_v_22_3_2(nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm,
      reg_nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1,
      reg_nv_scvector_cctor_nv_scvector_6_for_10_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1,
      {and_dcpl_847 , and_dcpl_852 , and_dcpl_855});
  assign nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_6_b = {1'b1 , Silu_for_else_if_mux1h_5_nl
      , Silu_for_else_if_mux1h_55_nl , Silu_for_else_if_mux1h_47_nl};
  wire [20:0] nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_7_a;
  assign nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_7_a = {Silu_for_else_if_Silu_for_else_if_or_itm
      , 20'b00110011001100110011};
  wire Silu_for_else_if_mux1h_2_nl;
  wire[2:0] Silu_for_else_if_mux1h_56_nl;
  wire[21:0] Silu_for_else_if_mux1h_48_nl;
  wire [26:0] nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_7_b;
  assign Silu_for_else_if_mux1h_2_nl = MUX1HOT_s_1_4_2(nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3,
      nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3,
      reg_nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0,
      reg_nv_scvector_cctor_nv_scvector_6_for_9_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0,
      {Silu_for_else_if_and_1_cse , Silu_for_else_if_and_2_cse , and_dcpl_852 , and_dcpl_855});
  assign Silu_for_else_if_mux1h_56_nl = MUX1HOT_v_3_4_2(nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0,
      nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0,
      reg_nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1,
      reg_nv_scvector_cctor_nv_scvector_6_for_9_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1,
      {Silu_for_else_if_and_1_cse , Silu_for_else_if_and_2_cse , and_dcpl_852 , and_dcpl_855});
  assign Silu_for_else_if_mux1h_48_nl = MUX1HOT_v_22_4_2(nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm,
      nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm,
      reg_nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1,
      reg_nv_scvector_cctor_nv_scvector_6_for_9_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1,
      {Silu_for_else_if_and_1_cse , Silu_for_else_if_and_2_cse , and_dcpl_852 , and_dcpl_855});
  assign nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_7_b = {1'b1 , Silu_for_else_if_mux1h_2_nl
      , Silu_for_else_if_mux1h_56_nl , Silu_for_else_if_mux1h_48_nl};
  wire  nl_ActUnit_ActUnitRun_rva_out_Push_mioi_inst_ActUnitRun_wten;
  assign nl_ActUnit_ActUnitRun_rva_out_Push_mioi_inst_ActUnitRun_wten = ~ ActUnitRun_wen;
  wire[31:0] ActUnit_PushAxiRsp_if_mux_11_nl;
  wire[31:0] ActUnit_PushAxiRsp_if_mux_10_nl;
  wire[31:0] ActUnit_PushAxiRsp_if_mux_9_nl;
  wire[31:0] ActUnit_PushAxiRsp_if_mux_8_nl;
  wire[31:0] ActUnit_PushAxiRsp_if_mux_7_nl;
  wire[31:0] ActUnit_PushAxiRsp_if_mux_6_nl;
  wire[31:0] ActUnit_PushAxiRsp_if_mux_5_nl;
  wire[31:0] ActUnit_PushAxiRsp_if_mux_4_nl;
  wire[31:0] ActUnit_PushAxiRsp_if_mux_3_nl;
  wire[31:0] ActUnit_PushAxiRsp_if_mux_2_nl;
  wire[31:0] ActUnit_PushAxiRsp_if_mux_1_nl;
  wire[31:0] ActUnit_PushAxiRsp_if_mux_nl;
  wire[7:0] act_mem_banks_read_read_data_mux_19_nl;
  wire[7:0] act_mem_banks_read_read_data_mux_18_nl;
  wire[7:0] act_mem_banks_read_read_data_mux_17_nl;
  wire[7:0] act_mem_banks_read_read_data_mux_16_nl;
  wire[7:0] act_mem_banks_read_read_data_mux_15_nl;
  wire[7:0] act_mem_banks_read_read_data_mux_14_nl;
  wire[7:0] act_mem_banks_read_read_data_mux_13_nl;
  wire[2:0] act_mem_banks_read_read_data_mux_12_nl;
  wire[4:0] act_mem_banks_read_read_data_mux_36_nl;
  wire[7:0] act_mem_banks_read_read_data_mux_11_nl;
  wire[2:0] act_mem_banks_read_read_data_mux_10_nl;
  wire[4:0] act_mem_banks_read_read_data_mux_9_nl;
  wire[7:0] act_mem_banks_read_read_data_mux_8_nl;
  wire[3:0] act_mem_banks_read_read_data_mux_7_nl;
  wire act_mem_banks_read_read_data_mux_37_nl;
  wire[2:0] act_mem_banks_read_read_data_mux_39_nl;
  wire[1:0] act_mem_banks_read_read_data_mux_6_nl;
  wire[1:0] act_mem_banks_read_read_data_mux_5_nl;
  wire act_mem_banks_read_read_data_mux_38_nl;
  wire[2:0] act_mem_banks_read_read_data_mux_40_nl;
  wire[7:0] act_mem_banks_read_read_data_mux_4_nl;
  wire[6:0] act_mem_banks_read_read_data_mux_3_nl;
  wire act_mem_banks_read_read_data_mux_2_nl;
  wire[6:0] act_mem_banks_read_read_data_mux_1_nl;
  wire act_mem_banks_read_read_data_mux_nl;
  wire [511:0] nl_ActUnit_ActUnitRun_rva_out_Push_mioi_inst_rva_out_Push_mioi_m_data_rsc_dat_ActUnitRun;
  assign ActUnit_PushAxiRsp_if_mux_11_nl = MUX_v_32_2_2(rva_out_reg_data_511_480_sva_dfm_3,
      act_mem_banks_read_read_data_lpi_1_dfm_1_511_480_mx1, act_read_req_valid_lpi_1_dfm_6);
  assign ActUnit_PushAxiRsp_if_mux_10_nl = MUX_v_32_2_2(rva_out_reg_data_479_448_sva_dfm_3,
      act_mem_banks_read_read_data_lpi_1_dfm_1_479_448_mx1, act_read_req_valid_lpi_1_dfm_6);
  assign ActUnit_PushAxiRsp_if_mux_9_nl = MUX_v_32_2_2(rva_out_reg_data_447_416_sva_dfm_3,
      act_mem_banks_read_read_data_lpi_1_dfm_1_447_416_mx1, act_read_req_valid_lpi_1_dfm_6);
  assign ActUnit_PushAxiRsp_if_mux_8_nl = MUX_v_32_2_2(rva_out_reg_data_415_384_sva_dfm_3,
      act_mem_banks_read_read_data_lpi_1_dfm_1_415_384_mx1, act_read_req_valid_lpi_1_dfm_6);
  assign ActUnit_PushAxiRsp_if_mux_7_nl = MUX_v_32_2_2(rva_out_reg_data_383_352_sva_dfm_3,
      act_mem_banks_read_read_data_lpi_1_dfm_1_383_352_mx1, act_read_req_valid_lpi_1_dfm_6);
  assign ActUnit_PushAxiRsp_if_mux_6_nl = MUX_v_32_2_2(rva_out_reg_data_351_320_sva_dfm_3,
      act_mem_banks_read_read_data_lpi_1_dfm_1_351_320_mx1, act_read_req_valid_lpi_1_dfm_6);
  assign ActUnit_PushAxiRsp_if_mux_5_nl = MUX_v_32_2_2(rva_out_reg_data_319_288_sva_dfm_3,
      act_mem_banks_read_read_data_lpi_1_dfm_1_319_288_mx1, act_read_req_valid_lpi_1_dfm_6);
  assign ActUnit_PushAxiRsp_if_mux_4_nl = MUX_v_32_2_2(rva_out_reg_data_287_256_sva_dfm_3,
      act_mem_banks_read_read_data_lpi_1_dfm_1_287_256_mx1, act_read_req_valid_lpi_1_dfm_6);
  assign ActUnit_PushAxiRsp_if_mux_3_nl = MUX_v_32_2_2(rva_out_reg_data_255_224_sva_dfm_3,
      act_mem_banks_read_read_data_lpi_1_dfm_1_255_224_mx1, act_read_req_valid_lpi_1_dfm_6);
  assign ActUnit_PushAxiRsp_if_mux_2_nl = MUX_v_32_2_2(rva_out_reg_data_223_192_sva_dfm_3,
      act_mem_banks_read_read_data_lpi_1_dfm_1_223_192_mx1, act_read_req_valid_lpi_1_dfm_6);
  assign ActUnit_PushAxiRsp_if_mux_1_nl = MUX_v_32_2_2(rva_out_reg_data_191_160_sva_dfm_3,
      act_mem_banks_read_read_data_lpi_1_dfm_1_191_160_mx1, act_read_req_valid_lpi_1_dfm_6);
  assign ActUnit_PushAxiRsp_if_mux_nl = MUX_v_32_2_2(rva_out_reg_data_159_128_sva_dfm_3,
      act_mem_banks_read_read_data_lpi_1_dfm_1_159_128_mx1, act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_19_nl = MUX_v_8_2_2(rva_out_reg_data_127_120_sva_dfm_3,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_127_96_mx1[31:24]), act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_18_nl = MUX_v_8_2_2(rva_out_reg_data_119_112_sva_dfm_3,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_127_96_mx1[23:16]), act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_17_nl = MUX_v_8_2_2(rva_out_reg_data_111_104_sva_dfm_3,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_127_96_mx1[15:8]), act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_16_nl = MUX_v_8_2_2(rva_out_reg_data_103_96_sva_dfm_3,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_127_96_mx1[7:0]), act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_15_nl = MUX_v_8_2_2(rva_out_reg_data_95_88_sva_dfm_3,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_95_64_mx1[31:24]), act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_14_nl = MUX_v_8_2_2(rva_out_reg_data_87_80_sva_dfm_3,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_95_64_mx1[23:16]), act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_13_nl = MUX_v_8_2_2(rva_out_reg_data_79_72_sva_dfm_3,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_95_64_mx1[15:8]), act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_12_nl = MUX_v_3_2_2(rva_out_reg_data_71_64_sva_dfm_3_7_5,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_95_64_mx1[7:5]), act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_36_nl = MUX_v_5_2_2(rva_out_reg_data_71_64_sva_dfm_3_4_0,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_95_64_mx1[4:0]), act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_11_nl = MUX_v_8_2_2(rva_out_reg_data_63_56_sva_dfm_3,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_63_32_mx1[31:24]), act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_10_nl = MUX_v_3_2_2(rva_out_reg_data_55_53_sva_dfm_3,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_63_32_mx1[23:21]), act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_9_nl = MUX_v_5_2_2(rva_out_reg_data_52_48_sva_dfm_3,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_63_32_mx1[20:16]), act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_8_nl = MUX_v_8_2_2(rva_out_reg_data_47_40_sva_dfm_3,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_63_32_mx1[15:8]), act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_7_nl = MUX_v_4_2_2(rva_out_reg_data_39_32_sva_dfm_3_7_4,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_63_32_mx1[7:4]), act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_37_nl = MUX_s_1_2_2(rva_out_reg_data_39_32_sva_dfm_3_3,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_63_32_mx1[3]), act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_39_nl = MUX_v_3_2_2(rva_out_reg_data_39_32_sva_dfm_3_2_0,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_63_32_mx1[2:0]), act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_6_nl = MUX_v_2_2_2(rva_out_reg_data_31_30_sva_dfm_3,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_31_0_mx1[31:30]), act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_5_nl = MUX_v_2_2_2(rva_out_reg_data_29_24_sva_dfm_3_5_4,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_31_0_mx1[29:28]), act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_38_nl = MUX_s_1_2_2(rva_out_reg_data_29_24_sva_dfm_3_3,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_31_0_mx1[27]), act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_40_nl = MUX_v_3_2_2(rva_out_reg_data_29_24_sva_dfm_3_2_0,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_31_0_mx1[26:24]), act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_4_nl = MUX_v_8_2_2(rva_out_reg_data_23_16_sva_dfm_3,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_31_0_mx1[23:16]), act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_3_nl = MUX_v_7_2_2(rva_out_reg_data_15_9_sva_dfm_3,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_31_0_mx1[15:9]), act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_2_nl = MUX_s_1_2_2(rva_out_reg_data_8_sva_dfm_3,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_31_0_mx1[8]), act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_1_nl = MUX_v_7_2_2(rva_out_reg_data_7_1_sva_dfm_3,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_31_0_mx1[7:1]), act_read_req_valid_lpi_1_dfm_6);
  assign act_mem_banks_read_read_data_mux_nl = MUX_s_1_2_2(rva_out_reg_data_0_sva_dfm_3,
      (act_mem_banks_read_read_data_lpi_1_dfm_1_31_0_mx1[0]), act_read_req_valid_lpi_1_dfm_6);
  assign nl_ActUnit_ActUnitRun_rva_out_Push_mioi_inst_rva_out_Push_mioi_m_data_rsc_dat_ActUnitRun
      = {ActUnit_PushAxiRsp_if_mux_11_nl , ActUnit_PushAxiRsp_if_mux_10_nl , ActUnit_PushAxiRsp_if_mux_9_nl
      , ActUnit_PushAxiRsp_if_mux_8_nl , ActUnit_PushAxiRsp_if_mux_7_nl , ActUnit_PushAxiRsp_if_mux_6_nl
      , ActUnit_PushAxiRsp_if_mux_5_nl , ActUnit_PushAxiRsp_if_mux_4_nl , ActUnit_PushAxiRsp_if_mux_3_nl
      , ActUnit_PushAxiRsp_if_mux_2_nl , ActUnit_PushAxiRsp_if_mux_1_nl , ActUnit_PushAxiRsp_if_mux_nl
      , act_mem_banks_read_read_data_mux_19_nl , act_mem_banks_read_read_data_mux_18_nl
      , act_mem_banks_read_read_data_mux_17_nl , act_mem_banks_read_read_data_mux_16_nl
      , act_mem_banks_read_read_data_mux_15_nl , act_mem_banks_read_read_data_mux_14_nl
      , act_mem_banks_read_read_data_mux_13_nl , act_mem_banks_read_read_data_mux_12_nl
      , act_mem_banks_read_read_data_mux_36_nl , act_mem_banks_read_read_data_mux_11_nl
      , act_mem_banks_read_read_data_mux_10_nl , act_mem_banks_read_read_data_mux_9_nl
      , act_mem_banks_read_read_data_mux_8_nl , act_mem_banks_read_read_data_mux_7_nl
      , act_mem_banks_read_read_data_mux_37_nl , act_mem_banks_read_read_data_mux_39_nl
      , act_mem_banks_read_read_data_mux_6_nl , act_mem_banks_read_read_data_mux_5_nl
      , act_mem_banks_read_read_data_mux_38_nl , act_mem_banks_read_read_data_mux_40_nl
      , act_mem_banks_read_read_data_mux_4_nl , act_mem_banks_read_read_data_mux_3_nl
      , act_mem_banks_read_read_data_mux_2_nl , act_mem_banks_read_read_data_mux_1_nl
      , act_mem_banks_read_read_data_mux_nl};
  wire  nl_ActUnit_ActUnitRun_output_port_Push_mioi_inst_ActUnitRun_wten;
  assign nl_ActUnit_ActUnitRun_output_port_Push_mioi_inst_ActUnitRun_wten = ~ ActUnitRun_wen;
  wire ActUnit_PushOutput_if_for_ActUnit_PushOutput_if_for_and_3_nl;
  wire[4:0] ActUnit_PushOutput_if_for_ActUnit_PushOutput_if_for_and_1_nl;
  wire[3:0] ActUnit_PushOutput_if_for_ActUnit_PushOutput_if_for_and_nl;
  wire[21:0] ActUnit_PushOutput_if_for_ActUnit_PushOutput_if_for_and_2_nl;
  wire [511:0] nl_ActUnit_ActUnitRun_output_port_Push_mioi_inst_output_port_Push_mioi_m_data_data_rsc_dat_ActUnitRun;
  assign ActUnit_PushOutput_if_for_ActUnit_PushOutput_if_for_and_3_nl = ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_31
      & ActUnit_PushOutput_if_for_and_27_seb_1;
  assign ActUnit_PushOutput_if_for_ActUnit_PushOutput_if_for_and_1_nl = MUX_v_5_2_2(5'b00000,
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_30_26, ActUnit_PushOutput_if_for_and_27_seb_1);
  assign ActUnit_PushOutput_if_for_ActUnit_PushOutput_if_for_and_nl = MUX_v_4_2_2(4'b0000,
      ({act_config_output_counter_sva_3 , act_config_output_counter_sva_2_0}), ActUnit_PushOutput_if_for_and_27_seb_1);
  assign ActUnit_PushOutput_if_for_ActUnit_PushOutput_if_for_and_2_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      reg_Silu_for_10_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1,
      ActUnit_PushOutput_if_for_and_27_seb_1);
  assign nl_ActUnit_ActUnitRun_output_port_Push_mioi_inst_output_port_Push_mioi_m_data_data_rsc_dat_ActUnitRun
      = {ActUnit_PushOutput_if_for_ActUnit_PushOutput_if_for_and_3_nl , ActUnit_PushOutput_if_for_ActUnit_PushOutput_if_for_and_1_nl
      , ActUnit_PushOutput_if_for_ActUnit_PushOutput_if_for_and_nl , ActUnit_PushOutput_if_for_ActUnit_PushOutput_if_for_and_2_nl
      , ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_1_31 , ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_1_30_26
      , ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_1_25 , ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_1_24_22
      , Silu_for_2_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0
      , ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_1_31 , ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_1_30_26
      , ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_1_25 , ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_1_24_22
      , reg_Silu_for_16_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1
      , ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_1_31 , ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_1_30_26
      , ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_1_25 , ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_1_24_22
      , reg_Silu_for_15_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1
      , ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_1_31 , ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_1_30_26
      , ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_1_25 , ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_1_24_22
      , reg_Silu_for_14_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1
      , ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_1_31 , ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_1_30_26
      , ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_1_25 , ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_1_24_22
      , reg_Silu_for_13_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1
      , ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_1_31 , ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_1_30_26
      , ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_1_25 , ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_1_24_22
      , Silu_for_y_8_sva_3_21_0 , ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_1_31
      , ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_1_30_26 , ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_1_25
      , ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_1_24_22 , Silu_for_y_1_sva_3_21_0
      , ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_1_31 , ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_1_30_26
      , ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_1_25 , ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_1_24_22
      , Silu_for_9_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0
      , ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_1_31 , ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_1_30_26
      , ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_1_25 , ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_1_24_22
      , Silu_for_7_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0
      , ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_1_31 , ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_1_30_26
      , ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_1_25 , ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_1_24_22
      , Silu_for_6_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0
      , ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_1_31 , ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_1_30_26
      , ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_1_25 , ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_1_24_22
      , Silu_for_5_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0
      , ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_1_31 , ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_1_30_26
      , ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_1_25 , ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_1_24_22
      , Silu_for_4_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0
      , ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_1_31 , ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_1_30_26
      , ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_1_25 , ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_1_24_22
      , Silu_for_3_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0
      , ActUnit_PushOutput_if_output_port_reg_data_data_1_sva_1_31 , rva_out_reg_data_71_64_sva_dfm_6_4_0
      , rva_out_reg_data_39_32_sva_dfm_6_3 , rva_out_reg_data_39_32_sva_dfm_6_2_0
      , reg_Silu_for_12_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1
      , ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_1_31 , ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_1_30_26
      , rva_out_reg_data_29_24_sva_dfm_6_3 , rva_out_reg_data_29_24_sva_dfm_6_2_0
      , reg_Silu_for_11_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1};
  wire [8:0] nl_ActUnit_ActUnitRun_output_port_Push_mioi_inst_output_port_Push_mioi_m_logical_addr_rsc_dat_ActUnitRun;
  assign nl_ActUnit_ActUnitRun_output_port_Push_mioi_inst_output_port_Push_mioi_m_logical_addr_rsc_dat_ActUnitRun
      = ({reg_act_config_output_counter_sva_dfm_3_ftd , reg_act_config_output_counter_sva_dfm_3_ftd_1_3
      , reg_act_config_output_counter_sva_dfm_3_ftd_1_2_0}) + act_config_output_addr_base_sva;
  wire  nl_ActUnit_ActUnitRun_done_Push_mioi_inst_ActUnitRun_wten;
  assign nl_ActUnit_ActUnitRun_done_Push_mioi_inst_ActUnitRun_wten = ~ ActUnitRun_wen;
  wire  nl_ActUnit_ActUnitRun_ActUnitRun_fsm_inst_while_C_0_tr0;
  assign nl_ActUnit_ActUnitRun_ActUnitRun_fsm_inst_while_C_0_tr0 = (act_config_in_InstFetch_mux_tmp[7:5]!=3'b001)
      | or_dcpl_450;
  wire  nl_ActUnit_ActUnitRun_ActUnitRun_fsm_inst_ActUnit_RunInst_case_2_for_C_0_tr0;
  assign nl_ActUnit_ActUnitRun_ActUnitRun_fsm_inst_ActUnit_RunInst_case_2_for_C_0_tr0
      = z_out[4];
  wire  nl_ActUnit_ActUnitRun_ActUnitRun_fsm_inst_while_C_3_tr0;
  assign nl_ActUnit_ActUnitRun_ActUnitRun_fsm_inst_while_C_3_tr0 = ~(ActUnit_RunInst_switch_lp_equal_tmp_3
      & is_start_sva);
  wire  nl_ActUnit_ActUnitRun_ActUnitRun_fsm_inst_ActUnit_PushOutput_if_for_C_0_tr0;
  assign nl_ActUnit_ActUnitRun_ActUnitRun_fsm_inst_ActUnit_PushOutput_if_for_C_0_tr0
      = z_out[4];
  wire  nl_ActUnit_ActUnitRun_ActUnitRun_fsm_inst_while_C_5_tr0;
  assign nl_ActUnit_ActUnitRun_ActUnitRun_fsm_inst_while_C_5_tr0 = (~ w_load_lpi_1_dfm_1)
      | act_config_is_zero_first_sva | (~ is_start_sva);
  wire  nl_ActUnit_ActUnitRun_ActUnitRun_fsm_inst_ActUnit_RunLoad_if_else_for_C_0_tr0;
  assign nl_ActUnit_ActUnitRun_ActUnitRun_fsm_inst_ActUnit_RunLoad_if_else_for_C_0_tr0
      = z_out[4];
  ActUnit_mgc_mul_pipe #(.width_a(32'sd25),
  .signd_a(32'sd0),
  .width_b(32'sd26),
  .signd_b(32'sd0),
  .width_z(32'sd51),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Gelu_for_1_else_else_else_if_mul_cmp (
      .a(nl_Gelu_for_1_else_else_else_if_mul_cmp_a[24:0]),
      .b(nl_Gelu_for_1_else_else_else_if_mul_cmp_b[25:0]),
      .clk(clk),
      .en(Gelu_for_1_else_else_else_if_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Gelu_for_1_else_else_else_if_mul_cmp_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd25),
  .signd_a(32'sd0),
  .width_b(32'sd26),
  .signd_b(32'sd0),
  .width_z(32'sd51),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Gelu_for_1_else_else_else_if_mul_cmp_1 (
      .a(nl_Gelu_for_1_else_else_else_if_mul_cmp_1_a[24:0]),
      .b(nl_Gelu_for_1_else_else_else_if_mul_cmp_1_b[25:0]),
      .clk(clk),
      .en(Gelu_for_1_else_else_else_if_mul_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Gelu_for_1_else_else_else_if_mul_cmp_1_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd25),
  .signd_a(32'sd0),
  .width_b(32'sd26),
  .signd_b(32'sd0),
  .width_z(32'sd51),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Gelu_for_1_else_else_else_if_mul_cmp_2 (
      .a(nl_Gelu_for_1_else_else_else_if_mul_cmp_2_a[24:0]),
      .b(nl_Gelu_for_1_else_else_else_if_mul_cmp_2_b[25:0]),
      .clk(clk),
      .en(Gelu_for_1_else_else_else_if_mul_cmp_2_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Gelu_for_1_else_else_else_if_mul_cmp_2_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd25),
  .signd_a(32'sd0),
  .width_b(32'sd26),
  .signd_b(32'sd0),
  .width_z(32'sd51),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Gelu_for_1_else_else_else_if_mul_cmp_3 (
      .a(nl_Gelu_for_1_else_else_else_if_mul_cmp_3_a[24:0]),
      .b(nl_Gelu_for_1_else_else_else_if_mul_cmp_3_b[25:0]),
      .clk(clk),
      .en(Gelu_for_1_else_else_else_if_mul_cmp_3_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Gelu_for_1_else_else_else_if_mul_cmp_3_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd25),
  .signd_a(32'sd0),
  .width_b(32'sd26),
  .signd_b(32'sd0),
  .width_z(32'sd51),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Gelu_for_1_else_else_else_if_mul_cmp_4 (
      .a(nl_Gelu_for_1_else_else_else_if_mul_cmp_4_a[24:0]),
      .b(nl_Gelu_for_1_else_else_else_if_mul_cmp_4_b[25:0]),
      .clk(clk),
      .en(Gelu_for_1_else_else_else_if_mul_cmp_4_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Gelu_for_1_else_else_else_if_mul_cmp_4_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd25),
  .signd_a(32'sd0),
  .width_b(32'sd26),
  .signd_b(32'sd0),
  .width_z(32'sd51),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Gelu_for_1_else_else_else_if_mul_cmp_5 (
      .a(nl_Gelu_for_1_else_else_else_if_mul_cmp_5_a[24:0]),
      .b(nl_Gelu_for_1_else_else_else_if_mul_cmp_5_b[25:0]),
      .clk(clk),
      .en(Gelu_for_1_else_else_else_if_mul_cmp_5_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Gelu_for_1_else_else_else_if_mul_cmp_5_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd25),
  .signd_a(32'sd0),
  .width_b(32'sd26),
  .signd_b(32'sd0),
  .width_z(32'sd51),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Gelu_for_1_else_else_else_if_mul_cmp_6 (
      .a(nl_Gelu_for_1_else_else_else_if_mul_cmp_6_a[24:0]),
      .b(nl_Gelu_for_1_else_else_else_if_mul_cmp_6_b[25:0]),
      .clk(clk),
      .en(Gelu_for_1_else_else_else_if_mul_cmp_6_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Gelu_for_1_else_else_else_if_mul_cmp_6_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd25),
  .signd_a(32'sd0),
  .width_b(32'sd26),
  .signd_b(32'sd0),
  .width_z(32'sd51),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Gelu_for_1_else_else_else_if_mul_cmp_7 (
      .a(nl_Gelu_for_1_else_else_else_if_mul_cmp_7_a[24:0]),
      .b(nl_Gelu_for_1_else_else_else_if_mul_cmp_7_b[25:0]),
      .clk(clk),
      .en(Gelu_for_1_else_else_else_if_mul_cmp_7_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Gelu_for_1_else_else_else_if_mul_cmp_7_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd25),
  .signd_a(32'sd0),
  .width_b(32'sd26),
  .signd_b(32'sd0),
  .width_z(32'sd51),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Gelu_for_1_else_else_else_if_mul_cmp_8 (
      .a(nl_Gelu_for_1_else_else_else_if_mul_cmp_8_a[24:0]),
      .b(nl_Gelu_for_1_else_else_else_if_mul_cmp_8_b[25:0]),
      .clk(clk),
      .en(Gelu_for_1_else_else_else_if_mul_cmp_8_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Gelu_for_1_else_else_else_if_mul_cmp_8_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd25),
  .signd_a(32'sd0),
  .width_b(32'sd26),
  .signd_b(32'sd0),
  .width_z(32'sd51),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Gelu_for_1_else_else_else_if_mul_cmp_9 (
      .a(nl_Gelu_for_1_else_else_else_if_mul_cmp_9_a[24:0]),
      .b(nl_Gelu_for_1_else_else_else_if_mul_cmp_9_b[25:0]),
      .clk(clk),
      .en(Gelu_for_1_else_else_else_if_mul_cmp_9_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Gelu_for_1_else_else_else_if_mul_cmp_9_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd25),
  .signd_a(32'sd0),
  .width_b(32'sd26),
  .signd_b(32'sd0),
  .width_z(32'sd51),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Gelu_for_1_else_else_else_if_mul_cmp_10 (
      .a(nl_Gelu_for_1_else_else_else_if_mul_cmp_10_a[24:0]),
      .b(nl_Gelu_for_1_else_else_else_if_mul_cmp_10_b[25:0]),
      .clk(clk),
      .en(Gelu_for_1_else_else_else_if_mul_cmp_10_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Gelu_for_1_else_else_else_if_mul_cmp_10_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd25),
  .signd_a(32'sd0),
  .width_b(32'sd26),
  .signd_b(32'sd0),
  .width_z(32'sd51),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Gelu_for_1_else_else_else_if_mul_cmp_11 (
      .a(nl_Gelu_for_1_else_else_else_if_mul_cmp_11_a[24:0]),
      .b(nl_Gelu_for_1_else_else_else_if_mul_cmp_11_b[25:0]),
      .clk(clk),
      .en(Gelu_for_1_else_else_else_if_mul_cmp_11_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Gelu_for_1_else_else_else_if_mul_cmp_11_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd25),
  .signd_a(32'sd0),
  .width_b(32'sd26),
  .signd_b(32'sd0),
  .width_z(32'sd51),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Gelu_for_1_else_else_else_if_mul_cmp_12 (
      .a(nl_Gelu_for_1_else_else_else_if_mul_cmp_12_a[24:0]),
      .b(nl_Gelu_for_1_else_else_else_if_mul_cmp_12_b[25:0]),
      .clk(clk),
      .en(Gelu_for_1_else_else_else_if_mul_cmp_12_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Gelu_for_1_else_else_else_if_mul_cmp_12_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd25),
  .signd_a(32'sd0),
  .width_b(32'sd26),
  .signd_b(32'sd0),
  .width_z(32'sd51),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Gelu_for_1_else_else_else_if_mul_cmp_13 (
      .a(nl_Gelu_for_1_else_else_else_if_mul_cmp_13_a[24:0]),
      .b(nl_Gelu_for_1_else_else_else_if_mul_cmp_13_b[25:0]),
      .clk(clk),
      .en(Gelu_for_1_else_else_else_if_mul_cmp_13_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Gelu_for_1_else_else_else_if_mul_cmp_13_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd25),
  .signd_a(32'sd0),
  .width_b(32'sd26),
  .signd_b(32'sd0),
  .width_z(32'sd51),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Gelu_for_1_else_else_else_if_mul_cmp_14 (
      .a(nl_Gelu_for_1_else_else_else_if_mul_cmp_14_a[24:0]),
      .b(nl_Gelu_for_1_else_else_else_if_mul_cmp_14_b[25:0]),
      .clk(clk),
      .en(Gelu_for_1_else_else_else_if_mul_cmp_14_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Gelu_for_1_else_else_else_if_mul_cmp_14_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd25),
  .signd_a(32'sd0),
  .width_b(32'sd26),
  .signd_b(32'sd0),
  .width_z(32'sd51),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Gelu_for_1_else_else_else_if_mul_cmp_15 (
      .a(nl_Gelu_for_1_else_else_else_if_mul_cmp_15_a[24:0]),
      .b(nl_Gelu_for_1_else_else_else_if_mul_cmp_15_b[25:0]),
      .clk(clk),
      .en(Gelu_for_1_else_else_else_if_mul_cmp_15_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Gelu_for_1_else_else_else_if_mul_cmp_15_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_b(32'sd25),
  .signd_b(32'sd1),
  .width_z(32'sd47),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Gelu_for_1_else_else_if_mul_cmp (
      .a(22'b1110111010010111100011),
      .b(nl_Gelu_for_1_else_else_if_mul_cmp_b[24:0]),
      .clk(clk),
      .en(Gelu_for_1_else_else_if_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Gelu_for_1_else_else_if_mul_cmp_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_b(32'sd25),
  .signd_b(32'sd1),
  .width_z(32'sd47),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Gelu_for_1_else_else_if_mul_cmp_1 (
      .a(22'b1110111010010111100011),
      .b(nl_Gelu_for_1_else_else_if_mul_cmp_1_b[24:0]),
      .clk(clk),
      .en(Gelu_for_1_else_else_if_mul_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Gelu_for_1_else_else_if_mul_cmp_1_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_b(32'sd25),
  .signd_b(32'sd1),
  .width_z(32'sd47),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Gelu_for_1_else_else_if_mul_cmp_2 (
      .a(22'b1110111010010111100011),
      .b(nl_Gelu_for_1_else_else_if_mul_cmp_2_b[24:0]),
      .clk(clk),
      .en(Gelu_for_1_else_else_if_mul_cmp_2_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Gelu_for_1_else_else_if_mul_cmp_2_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_b(32'sd25),
  .signd_b(32'sd1),
  .width_z(32'sd47),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Gelu_for_1_else_else_if_mul_cmp_3 (
      .a(22'b1110111010010111100011),
      .b(nl_Gelu_for_1_else_else_if_mul_cmp_3_b[24:0]),
      .clk(clk),
      .en(Gelu_for_1_else_else_if_mul_cmp_3_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Gelu_for_1_else_else_if_mul_cmp_3_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_b(32'sd25),
  .signd_b(32'sd1),
  .width_z(32'sd47),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Gelu_for_1_else_else_if_mul_cmp_4 (
      .a(22'b1110111010010111100011),
      .b(nl_Gelu_for_1_else_else_if_mul_cmp_4_b[24:0]),
      .clk(clk),
      .en(Gelu_for_1_else_else_if_mul_cmp_4_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Gelu_for_1_else_else_if_mul_cmp_4_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_b(32'sd25),
  .signd_b(32'sd1),
  .width_z(32'sd47),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Gelu_for_1_else_else_if_mul_cmp_5 (
      .a(22'b1110111010010111100011),
      .b(nl_Gelu_for_1_else_else_if_mul_cmp_5_b[24:0]),
      .clk(clk),
      .en(Gelu_for_1_else_else_if_mul_cmp_5_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Gelu_for_1_else_else_if_mul_cmp_5_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_b(32'sd25),
  .signd_b(32'sd1),
  .width_z(32'sd47),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Gelu_for_1_else_else_if_mul_cmp_6 (
      .a(22'b1110111010010111100011),
      .b(nl_Gelu_for_1_else_else_if_mul_cmp_6_b[24:0]),
      .clk(clk),
      .en(Gelu_for_1_else_else_if_mul_cmp_6_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Gelu_for_1_else_else_if_mul_cmp_6_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_b(32'sd25),
  .signd_b(32'sd1),
  .width_z(32'sd47),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Gelu_for_1_else_else_if_mul_cmp_7 (
      .a(22'b1110111010010111100011),
      .b(nl_Gelu_for_1_else_else_if_mul_cmp_7_b[24:0]),
      .clk(clk),
      .en(Gelu_for_1_else_else_if_mul_cmp_7_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Gelu_for_1_else_else_if_mul_cmp_7_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_b(32'sd25),
  .signd_b(32'sd1),
  .width_z(32'sd47),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Gelu_for_1_else_else_if_mul_cmp_8 (
      .a(22'b1110111010010111100011),
      .b(nl_Gelu_for_1_else_else_if_mul_cmp_8_b[24:0]),
      .clk(clk),
      .en(Gelu_for_1_else_else_if_mul_cmp_8_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Gelu_for_1_else_else_if_mul_cmp_8_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_b(32'sd25),
  .signd_b(32'sd1),
  .width_z(32'sd47),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Gelu_for_1_else_else_if_mul_cmp_9 (
      .a(22'b1110111010010111100011),
      .b(nl_Gelu_for_1_else_else_if_mul_cmp_9_b[24:0]),
      .clk(clk),
      .en(Gelu_for_1_else_else_if_mul_cmp_9_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Gelu_for_1_else_else_if_mul_cmp_9_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_b(32'sd25),
  .signd_b(32'sd1),
  .width_z(32'sd47),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Gelu_for_1_else_else_if_mul_cmp_10 (
      .a(22'b1110111010010111100011),
      .b(nl_Gelu_for_1_else_else_if_mul_cmp_10_b[24:0]),
      .clk(clk),
      .en(Gelu_for_1_else_else_if_mul_cmp_10_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Gelu_for_1_else_else_if_mul_cmp_10_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_b(32'sd25),
  .signd_b(32'sd1),
  .width_z(32'sd47),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Gelu_for_1_else_else_if_mul_cmp_11 (
      .a(22'b1110111010010111100011),
      .b(nl_Gelu_for_1_else_else_if_mul_cmp_11_b[24:0]),
      .clk(clk),
      .en(Gelu_for_1_else_else_if_mul_cmp_11_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Gelu_for_1_else_else_if_mul_cmp_11_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_b(32'sd25),
  .signd_b(32'sd1),
  .width_z(32'sd47),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Gelu_for_1_else_else_if_mul_cmp_12 (
      .a(22'b1110111010010111100011),
      .b(nl_Gelu_for_1_else_else_if_mul_cmp_12_b[24:0]),
      .clk(clk),
      .en(Gelu_for_1_else_else_if_mul_cmp_12_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Gelu_for_1_else_else_if_mul_cmp_12_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_b(32'sd25),
  .signd_b(32'sd1),
  .width_z(32'sd47),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Gelu_for_1_else_else_if_mul_cmp_13 (
      .a(22'b1110111010010111100011),
      .b(nl_Gelu_for_1_else_else_if_mul_cmp_13_b[24:0]),
      .clk(clk),
      .en(Gelu_for_1_else_else_if_mul_cmp_13_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Gelu_for_1_else_else_if_mul_cmp_13_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_b(32'sd25),
  .signd_b(32'sd1),
  .width_z(32'sd47),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Gelu_for_1_else_else_if_mul_cmp_14 (
      .a(22'b1110111010010111100011),
      .b(nl_Gelu_for_1_else_else_if_mul_cmp_14_b[24:0]),
      .clk(clk),
      .en(Gelu_for_1_else_else_if_mul_cmp_14_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Gelu_for_1_else_else_if_mul_cmp_14_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_b(32'sd25),
  .signd_b(32'sd1),
  .width_z(32'sd47),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Gelu_for_1_else_else_if_mul_cmp_15 (
      .a(22'b1110111010010111100011),
      .b(nl_Gelu_for_1_else_else_if_mul_cmp_15_b[24:0]),
      .clk(clk),
      .en(Gelu_for_1_else_else_if_mul_cmp_15_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Gelu_for_1_else_else_if_mul_cmp_15_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd21),
  .signd_a(32'sd1),
  .width_b(32'sd27),
  .signd_b(32'sd1),
  .width_z(32'sd48),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Silu_for_1_else_if_Silu_for_else_if_mul_cmp (
      .a(nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_a[20:0]),
      .b(nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_b[26:0]),
      .clk(clk),
      .en(Silu_for_1_else_if_Silu_for_else_if_mul_cmp_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Silu_for_1_else_if_Silu_for_else_if_mul_cmp_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd21),
  .signd_a(32'sd1),
  .width_b(32'sd27),
  .signd_b(32'sd1),
  .width_z(32'sd48),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Silu_for_1_else_if_Silu_for_else_if_mul_cmp_1 (
      .a(nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_1_a[20:0]),
      .b(nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_1_b[26:0]),
      .clk(clk),
      .en(Silu_for_1_else_if_Silu_for_else_if_mul_cmp_1_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Silu_for_1_else_if_Silu_for_else_if_mul_cmp_1_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd21),
  .signd_a(32'sd1),
  .width_b(32'sd27),
  .signd_b(32'sd1),
  .width_z(32'sd48),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Silu_for_1_else_if_Silu_for_else_if_mul_cmp_2 (
      .a(nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_2_a[20:0]),
      .b(nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_2_b[26:0]),
      .clk(clk),
      .en(Silu_for_1_else_if_Silu_for_else_if_mul_cmp_2_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Silu_for_1_else_if_Silu_for_else_if_mul_cmp_2_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd21),
  .signd_a(32'sd1),
  .width_b(32'sd27),
  .signd_b(32'sd1),
  .width_z(32'sd48),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Silu_for_1_else_if_Silu_for_else_if_mul_cmp_3 (
      .a(nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_3_a[20:0]),
      .b(nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_3_b[26:0]),
      .clk(clk),
      .en(Silu_for_1_else_if_Silu_for_else_if_mul_cmp_3_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Silu_for_1_else_if_Silu_for_else_if_mul_cmp_3_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd21),
  .signd_a(32'sd1),
  .width_b(32'sd27),
  .signd_b(32'sd1),
  .width_z(32'sd48),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Silu_for_1_else_if_Silu_for_else_if_mul_cmp_4 (
      .a(nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_4_a[20:0]),
      .b(nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_4_b[26:0]),
      .clk(clk),
      .en(Silu_for_1_else_if_Silu_for_else_if_mul_cmp_4_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Silu_for_1_else_if_Silu_for_else_if_mul_cmp_4_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd21),
  .signd_a(32'sd1),
  .width_b(32'sd27),
  .signd_b(32'sd1),
  .width_z(32'sd48),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Silu_for_1_else_if_Silu_for_else_if_mul_cmp_5 (
      .a(nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_5_a[20:0]),
      .b(nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_5_b[26:0]),
      .clk(clk),
      .en(Silu_for_1_else_if_Silu_for_else_if_mul_cmp_5_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Silu_for_1_else_if_Silu_for_else_if_mul_cmp_5_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd21),
  .signd_a(32'sd1),
  .width_b(32'sd27),
  .signd_b(32'sd1),
  .width_z(32'sd48),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Silu_for_1_else_if_Silu_for_else_if_mul_cmp_6 (
      .a(nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_6_a[20:0]),
      .b(nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_6_b[26:0]),
      .clk(clk),
      .en(Silu_for_1_else_if_Silu_for_else_if_mul_cmp_6_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Silu_for_1_else_if_Silu_for_else_if_mul_cmp_6_z)
    );
  ActUnit_mgc_mul_pipe #(.width_a(32'sd21),
  .signd_a(32'sd1),
  .width_b(32'sd27),
  .signd_b(32'sd1),
  .width_z(32'sd48),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd1)) Silu_for_1_else_if_Silu_for_else_if_mul_cmp_7 (
      .a(nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_7_a[20:0]),
      .b(nl_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_7_b[26:0]),
      .clk(clk),
      .en(Silu_for_1_else_if_Silu_for_else_if_mul_cmp_7_en),
      .a_rst(rst),
      .s_rst(1'b1),
      .z(Silu_for_1_else_if_Silu_for_else_if_mul_cmp_7_z)
    );
  ActUnit_ActUnit_ActUnitRun_rva_in_PopNB_mioi ActUnit_ActUnitRun_rva_in_PopNB_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_in_vld(rva_in_vld),
      .rva_in_rdy(rva_in_rdy),
      .rva_in_dat(rva_in_dat),
      .ActUnitRun_wen(ActUnitRun_wen),
      .ActUnitRun_wten(ActUnitRun_wten),
      .rva_in_PopNB_mioi_oswt(reg_rva_in_PopNB_mioi_iswt0_cse),
      .rva_in_PopNB_mioi_data_data_rsc_z_mxwt(rva_in_PopNB_mioi_data_data_rsc_z_mxwt),
      .rva_in_PopNB_mioi_data_addr_rsc_z_mxwt(rva_in_PopNB_mioi_data_addr_rsc_z_mxwt),
      .rva_in_PopNB_mioi_data_rw_rsc_z_mxwt(rva_in_PopNB_mioi_data_rw_rsc_z_mxwt),
      .rva_in_PopNB_mioi_return_rsc_z_mxwt(rva_in_PopNB_mioi_return_rsc_z_mxwt),
      .rva_in_PopNB_mioi_oswt_pff(and_1116_rmff)
    );
  ActUnit_ActUnit_ActUnitRun_act_port_PopNB_mioi ActUnit_ActUnitRun_act_port_PopNB_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .act_port_vld(act_port_vld),
      .act_port_rdy(act_port_rdy),
      .act_port_dat(act_port_dat),
      .ActUnitRun_wen(ActUnitRun_wen),
      .ActUnitRun_wten(ActUnitRun_wten),
      .act_port_PopNB_mioi_oswt(reg_act_port_PopNB_mioi_iswt0_cse),
      .act_port_PopNB_mioi_data_data_rsc_z_mxwt(act_port_PopNB_mioi_data_data_rsc_z_mxwt),
      .act_port_PopNB_mioi_return_rsc_z_mxwt(act_port_PopNB_mioi_return_rsc_z_mxwt),
      .act_port_PopNB_mioi_oswt_pff(and_1113_rmff)
    );
  ActUnit_ActUnit_ActUnitRun_rva_out_Push_mioi ActUnit_ActUnitRun_rva_out_Push_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .rva_out_vld(rva_out_vld),
      .rva_out_rdy(rva_out_rdy),
      .rva_out_dat(rva_out_dat),
      .ActUnitRun_wten(nl_ActUnit_ActUnitRun_rva_out_Push_mioi_inst_ActUnitRun_wten),
      .rva_out_Push_mioi_oswt(reg_rva_out_Push_mioi_iswt0_cse),
      .rva_out_Push_mioi_wen_comp(rva_out_Push_mioi_wen_comp),
      .rva_out_Push_mioi_m_data_rsc_dat_ActUnitRun(nl_ActUnit_ActUnitRun_rva_out_Push_mioi_inst_rva_out_Push_mioi_m_data_rsc_dat_ActUnitRun[511:0]),
      .rva_out_Push_mioi_oswt_pff(and_1108_rmff)
    );
  ActUnit_ActUnit_ActUnitRun_start_PopNB_mioi ActUnit_ActUnitRun_start_PopNB_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .start_vld(start_vld),
      .start_rdy(start_rdy),
      .start_dat(start_dat),
      .ActUnitRun_wen(ActUnitRun_wen),
      .ActUnitRun_wten(ActUnitRun_wten),
      .start_PopNB_mioi_oswt(reg_start_PopNB_mioi_iswt0_cse),
      .start_PopNB_mioi_data_rsc_z_mxwt(start_PopNB_mioi_data_rsc_z_mxwt),
      .start_PopNB_mioi_return_rsc_z_mxwt(start_PopNB_mioi_return_rsc_z_mxwt),
      .start_PopNB_mioi_oswt_pff(and_1106_rmff)
    );
  ActUnit_ActUnit_ActUnitRun_output_port_Push_mioi ActUnit_ActUnitRun_output_port_Push_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .output_port_vld(output_port_vld),
      .output_port_rdy(output_port_rdy),
      .output_port_dat(output_port_dat),
      .ActUnitRun_wten(nl_ActUnit_ActUnitRun_output_port_Push_mioi_inst_ActUnitRun_wten),
      .output_port_Push_mioi_oswt(reg_output_port_Push_mioi_iswt0_cse),
      .output_port_Push_mioi_wen_comp(output_port_Push_mioi_wen_comp),
      .output_port_Push_mioi_m_data_data_rsc_dat_ActUnitRun(nl_ActUnit_ActUnitRun_output_port_Push_mioi_inst_output_port_Push_mioi_m_data_data_rsc_dat_ActUnitRun[511:0]),
      .output_port_Push_mioi_m_logical_addr_rsc_dat_ActUnitRun(nl_ActUnit_ActUnitRun_output_port_Push_mioi_inst_output_port_Push_mioi_m_logical_addr_rsc_dat_ActUnitRun[7:0]),
      .output_port_Push_mioi_oswt_pff(and_1102_rmff)
    );
  ActUnit_ActUnit_ActUnitRun_done_Push_mioi ActUnit_ActUnitRun_done_Push_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .done_vld(done_vld),
      .done_rdy(done_rdy),
      .done_dat(done_dat),
      .ActUnitRun_wten(nl_ActUnit_ActUnitRun_done_Push_mioi_inst_ActUnitRun_wten),
      .done_Push_mioi_oswt(reg_done_Push_mioi_iswt0_cse),
      .done_Push_mioi_wen_comp(done_Push_mioi_wen_comp),
      .done_Push_mioi_oswt_pff(and_1097_rmff)
    );
  ActUnit_ActUnit_ActUnitRun_wait_dp ActUnit_ActUnitRun_wait_dp_inst (
      .ActUnitRun_wen(ActUnitRun_wen),
      .Gelu_for_1_else_else_else_if_mul_cmp_cgo(reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_cse),
      .Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg(and_1088_rmff),
      .Gelu_for_1_else_else_else_if_mul_cmp_en(Gelu_for_1_else_else_else_if_mul_cmp_en),
      .Gelu_for_1_else_else_else_if_mul_cmp_cgo_1(reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_1_cse),
      .Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_1(and_1082_rmff),
      .Gelu_for_1_else_else_else_if_mul_cmp_1_en(Gelu_for_1_else_else_else_if_mul_cmp_1_en),
      .Gelu_for_1_else_else_else_if_mul_cmp_cgo_2(reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_2_cse),
      .Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_2(and_1076_rmff),
      .Gelu_for_1_else_else_else_if_mul_cmp_2_en(Gelu_for_1_else_else_else_if_mul_cmp_2_en),
      .Gelu_for_1_else_else_else_if_mul_cmp_cgo_3(reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_3_cse),
      .Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_3(and_1070_rmff),
      .Gelu_for_1_else_else_else_if_mul_cmp_3_en(Gelu_for_1_else_else_else_if_mul_cmp_3_en),
      .Gelu_for_1_else_else_else_if_mul_cmp_cgo_4(reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_4_cse),
      .Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_4(and_1064_rmff),
      .Gelu_for_1_else_else_else_if_mul_cmp_4_en(Gelu_for_1_else_else_else_if_mul_cmp_4_en),
      .Gelu_for_1_else_else_else_if_mul_cmp_cgo_5(reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_5_cse),
      .Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_5(and_1058_rmff),
      .Gelu_for_1_else_else_else_if_mul_cmp_5_en(Gelu_for_1_else_else_else_if_mul_cmp_5_en),
      .Gelu_for_1_else_else_else_if_mul_cmp_cgo_6(reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_6_cse),
      .Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_6(and_1052_rmff),
      .Gelu_for_1_else_else_else_if_mul_cmp_6_en(Gelu_for_1_else_else_else_if_mul_cmp_6_en),
      .Gelu_for_1_else_else_else_if_mul_cmp_cgo_7(reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_7_cse),
      .Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_7(and_1046_rmff),
      .Gelu_for_1_else_else_else_if_mul_cmp_7_en(Gelu_for_1_else_else_else_if_mul_cmp_7_en),
      .Gelu_for_1_else_else_else_if_mul_cmp_cgo_8(reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_8_cse),
      .Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_8(and_1040_rmff),
      .Gelu_for_1_else_else_else_if_mul_cmp_8_en(Gelu_for_1_else_else_else_if_mul_cmp_8_en),
      .Gelu_for_1_else_else_else_if_mul_cmp_cgo_9(reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_9_cse),
      .Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_9(and_1034_rmff),
      .Gelu_for_1_else_else_else_if_mul_cmp_9_en(Gelu_for_1_else_else_else_if_mul_cmp_9_en),
      .Gelu_for_1_else_else_else_if_mul_cmp_cgo_10(reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_10_cse),
      .Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_10(and_1028_rmff),
      .Gelu_for_1_else_else_else_if_mul_cmp_10_en(Gelu_for_1_else_else_else_if_mul_cmp_10_en),
      .Gelu_for_1_else_else_else_if_mul_cmp_cgo_11(reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_11_cse),
      .Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_11(and_1022_rmff),
      .Gelu_for_1_else_else_else_if_mul_cmp_11_en(Gelu_for_1_else_else_else_if_mul_cmp_11_en),
      .Gelu_for_1_else_else_else_if_mul_cmp_cgo_12(reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_12_cse),
      .Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_12(and_1016_rmff),
      .Gelu_for_1_else_else_else_if_mul_cmp_12_en(Gelu_for_1_else_else_else_if_mul_cmp_12_en),
      .Gelu_for_1_else_else_else_if_mul_cmp_cgo_13(reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_13_cse),
      .Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_13(and_1010_rmff),
      .Gelu_for_1_else_else_else_if_mul_cmp_13_en(Gelu_for_1_else_else_else_if_mul_cmp_13_en),
      .Gelu_for_1_else_else_else_if_mul_cmp_cgo_14(reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_14_cse),
      .Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_14(and_1004_rmff),
      .Gelu_for_1_else_else_else_if_mul_cmp_14_en(Gelu_for_1_else_else_else_if_mul_cmp_14_en),
      .Gelu_for_1_else_else_else_if_mul_cmp_cgo_15(reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_15_cse),
      .Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_unreg_15(and_998_rmff),
      .Gelu_for_1_else_else_else_if_mul_cmp_15_en(Gelu_for_1_else_else_else_if_mul_cmp_15_en),
      .Gelu_for_1_else_else_if_mul_cmp_cgo(reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_cse),
      .Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg(and_990_rmff),
      .Gelu_for_1_else_else_if_mul_cmp_en(Gelu_for_1_else_else_if_mul_cmp_en),
      .Gelu_for_1_else_else_if_mul_cmp_cgo_1(reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_1_cse),
      .Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_1(and_985_rmff),
      .Gelu_for_1_else_else_if_mul_cmp_1_en(Gelu_for_1_else_else_if_mul_cmp_1_en),
      .Gelu_for_1_else_else_if_mul_cmp_cgo_2(reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_2_cse),
      .Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_2(and_980_rmff),
      .Gelu_for_1_else_else_if_mul_cmp_2_en(Gelu_for_1_else_else_if_mul_cmp_2_en),
      .Gelu_for_1_else_else_if_mul_cmp_cgo_3(reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_3_cse),
      .Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_3(and_975_rmff),
      .Gelu_for_1_else_else_if_mul_cmp_3_en(Gelu_for_1_else_else_if_mul_cmp_3_en),
      .Gelu_for_1_else_else_if_mul_cmp_cgo_4(reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_4_cse),
      .Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_4(and_970_rmff),
      .Gelu_for_1_else_else_if_mul_cmp_4_en(Gelu_for_1_else_else_if_mul_cmp_4_en),
      .Gelu_for_1_else_else_if_mul_cmp_cgo_5(reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_5_cse),
      .Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_5(and_965_rmff),
      .Gelu_for_1_else_else_if_mul_cmp_5_en(Gelu_for_1_else_else_if_mul_cmp_5_en),
      .Gelu_for_1_else_else_if_mul_cmp_cgo_6(reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_6_cse),
      .Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_6(and_960_rmff),
      .Gelu_for_1_else_else_if_mul_cmp_6_en(Gelu_for_1_else_else_if_mul_cmp_6_en),
      .Gelu_for_1_else_else_if_mul_cmp_cgo_7(reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_7_cse),
      .Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_7(and_955_rmff),
      .Gelu_for_1_else_else_if_mul_cmp_7_en(Gelu_for_1_else_else_if_mul_cmp_7_en),
      .Gelu_for_1_else_else_if_mul_cmp_cgo_8(reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_8_cse),
      .Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_8(and_950_rmff),
      .Gelu_for_1_else_else_if_mul_cmp_8_en(Gelu_for_1_else_else_if_mul_cmp_8_en),
      .Gelu_for_1_else_else_if_mul_cmp_cgo_9(reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_9_cse),
      .Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_9(and_945_rmff),
      .Gelu_for_1_else_else_if_mul_cmp_9_en(Gelu_for_1_else_else_if_mul_cmp_9_en),
      .Gelu_for_1_else_else_if_mul_cmp_cgo_10(reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_10_cse),
      .Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_10(and_940_rmff),
      .Gelu_for_1_else_else_if_mul_cmp_10_en(Gelu_for_1_else_else_if_mul_cmp_10_en),
      .Gelu_for_1_else_else_if_mul_cmp_cgo_11(reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_11_cse),
      .Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_11(and_935_rmff),
      .Gelu_for_1_else_else_if_mul_cmp_11_en(Gelu_for_1_else_else_if_mul_cmp_11_en),
      .Gelu_for_1_else_else_if_mul_cmp_cgo_12(reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_12_cse),
      .Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_12(and_930_rmff),
      .Gelu_for_1_else_else_if_mul_cmp_12_en(Gelu_for_1_else_else_if_mul_cmp_12_en),
      .Gelu_for_1_else_else_if_mul_cmp_cgo_13(reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_13_cse),
      .Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_13(and_925_rmff),
      .Gelu_for_1_else_else_if_mul_cmp_13_en(Gelu_for_1_else_else_if_mul_cmp_13_en),
      .Gelu_for_1_else_else_if_mul_cmp_cgo_14(reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_14_cse),
      .Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_14(and_920_rmff),
      .Gelu_for_1_else_else_if_mul_cmp_14_en(Gelu_for_1_else_else_if_mul_cmp_14_en),
      .Gelu_for_1_else_else_if_mul_cmp_cgo_15(reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_15_cse),
      .Gelu_for_1_else_else_if_mul_cmp_cgo_ir_unreg_15(and_915_rmff),
      .Gelu_for_1_else_else_if_mul_cmp_15_en(Gelu_for_1_else_else_if_mul_cmp_15_en),
      .Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo(reg_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_cse),
      .Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_unreg(and_906_rmff),
      .Silu_for_1_else_if_Silu_for_else_if_mul_cmp_en(Silu_for_1_else_if_Silu_for_else_if_mul_cmp_en),
      .Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_1(reg_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_1_cse),
      .Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_unreg_1(and_905_rmff),
      .Silu_for_1_else_if_Silu_for_else_if_mul_cmp_1_en(Silu_for_1_else_if_Silu_for_else_if_mul_cmp_1_en),
      .Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_2(reg_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_2_cse),
      .Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_unreg_2(and_904_rmff),
      .Silu_for_1_else_if_Silu_for_else_if_mul_cmp_2_en(Silu_for_1_else_if_Silu_for_else_if_mul_cmp_2_en),
      .Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_3(reg_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_3_cse),
      .Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_unreg_3(and_903_rmff),
      .Silu_for_1_else_if_Silu_for_else_if_mul_cmp_3_en(Silu_for_1_else_if_Silu_for_else_if_mul_cmp_3_en),
      .Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_4(reg_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_4_cse),
      .Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_unreg_4(and_902_rmff),
      .Silu_for_1_else_if_Silu_for_else_if_mul_cmp_4_en(Silu_for_1_else_if_Silu_for_else_if_mul_cmp_4_en),
      .Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_5(reg_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_5_cse),
      .Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_unreg_5(and_901_rmff),
      .Silu_for_1_else_if_Silu_for_else_if_mul_cmp_5_en(Silu_for_1_else_if_Silu_for_else_if_mul_cmp_5_en),
      .Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_6(reg_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_6_cse),
      .Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_unreg_6(and_900_rmff),
      .Silu_for_1_else_if_Silu_for_else_if_mul_cmp_6_en(Silu_for_1_else_if_Silu_for_else_if_mul_cmp_6_en),
      .Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_7(reg_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_7_cse),
      .Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_unreg_7(and_899_rmff),
      .Silu_for_1_else_if_Silu_for_else_if_mul_cmp_7_en(Silu_for_1_else_if_Silu_for_else_if_mul_cmp_7_en)
    );
  ActUnit_ActUnit_ActUnitRun_staller ActUnit_ActUnitRun_staller_inst (
      .clk(clk),
      .rst(rst),
      .ActUnitRun_wen(ActUnitRun_wen),
      .ActUnitRun_wten(ActUnitRun_wten),
      .rva_out_Push_mioi_wen_comp(rva_out_Push_mioi_wen_comp),
      .output_port_Push_mioi_wen_comp(output_port_Push_mioi_wen_comp),
      .done_Push_mioi_wen_comp(done_Push_mioi_wen_comp)
    );
  ActUnit_ActUnit_ActUnitRun_ActUnitRun_fsm ActUnit_ActUnitRun_ActUnitRun_fsm_inst
      (
      .clk(clk),
      .rst(rst),
      .ActUnitRun_wen(ActUnitRun_wen),
      .fsm_output(fsm_output),
      .while_C_0_tr0(nl_ActUnit_ActUnitRun_ActUnitRun_fsm_inst_while_C_0_tr0),
      .ActUnit_RunInst_case_2_for_C_0_tr0(nl_ActUnit_ActUnitRun_ActUnitRun_fsm_inst_ActUnit_RunInst_case_2_for_C_0_tr0),
      .while_C_3_tr0(nl_ActUnit_ActUnitRun_ActUnitRun_fsm_inst_while_C_3_tr0),
      .ActUnit_PushOutput_if_for_C_0_tr0(nl_ActUnit_ActUnitRun_ActUnitRun_fsm_inst_ActUnit_PushOutput_if_for_C_0_tr0),
      .while_C_5_tr0(nl_ActUnit_ActUnitRun_ActUnitRun_fsm_inst_while_C_5_tr0),
      .ActUnit_RunLoad_if_else_for_C_0_tr0(nl_ActUnit_ActUnitRun_ActUnitRun_fsm_inst_ActUnit_RunLoad_if_else_for_C_0_tr0)
    );
  assign act_mem_banks_write_if_for_if_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_332);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb = act_mem_banks_write_if_for_if_mux_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 146
  // psl default clock = (posedge clk);
  // psl ActUnit_ActUnitRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb );
  assign act_mem_banks_write_if_for_if_mux_1_cse = MUX1HOT_s_1_1_2(ActUnitRun_wen,
      and_dcpl_332);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb = act_mem_banks_write_if_for_if_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb = act_mem_banks_write_if_for_if_mux_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 147
  // psl ActUnit_ActUnitRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb = act_mem_banks_write_if_for_if_mux_1_cse;
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb
      = act_mem_banks_write_if_for_if_mux_cse;
  // assert(bankread_req_valid[bank] == false && "Bank read and write valid cannot be true simultaneously for single-port RAM") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/ArbitratedScratchpadDP.h: line 196
  // psl ActUnit_ActUnitRun_ArbitratedScratchpadDP_h_ln196_assert_bankread_req_validOS_bank_CS_eq_false_and_Bankreadandwritevalidcannotbetruesimultaneouslyforsingle_m_portRAM : assert always ( rst &&  pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb  -> pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_prb );
  assign pbankread_req_valid_bank_false_Bank_read_and_write_valid_cannot_be_true_simultaneously_for_single_port_RAM_ctrl_prb
      = act_mem_banks_write_if_for_if_mux_1_cse;
  assign act_mem_banks_read_for_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_dcpl_337);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_1 = act_mem_banks_read_for_mux_cse;
  // assert(bank_sel<NumBanks && "bank index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 126
  // psl ActUnit_ActUnitRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bankindexoutofbounds : assert always ( rst &&  pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_1  -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_1 );
  assign act_mem_banks_read_for_mux_1_cse = MUX1HOT_s_1_1_2(ActUnitRun_wen, and_dcpl_337);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_1 = act_mem_banks_read_for_mux_1_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_1 = act_mem_banks_read_for_mux_cse;
  // assert(idx<NumEntriesPerBank && "local index out of bounds") - /cad/mentor/2024.2_1/Mgc_home/shared/pkgs/matchlib/cmod/include/mem_array.h: line 127
  // psl ActUnit_ActUnitRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_localindexoutofbounds : assert always ( rst &&  pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_1  -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_1 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_1 = act_mem_banks_read_for_mux_1_cse;
  assign or_866_nl = (act_config_in_InstFetch_return_sva_7_2[2]) | (~ (fsm_output[0]));
  assign mux_330_nl = MUX_s_1_2_2((fsm_output[0]), or_866_nl, fsm_output[1]);
  assign Silu_for_else_if_Silu_for_else_if_or_itm = ((act_config_in_InstFetch_mux_tmp[4])
      & (~((~ mux_330_nl) | or_dcpl_457))) | and_dcpl_855;
  assign or_872_nl = (~ Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)
      | Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign mux_337_nl = MUX_s_1_2_2(mux_tmp_318, nand_tmp_23, or_872_nl);
  assign or_871_nl = (~ Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)
      | Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign mux_338_nl = MUX_s_1_2_2(mux_tmp_317, mux_337_nl, or_871_nl);
  assign nor_143_nl = ~(Gelu_for_1_else_slc_32_svs | (~ Gelu_for_1_slc_32_1_svs));
  assign mux_335_nl = MUX_s_1_2_2(nand_tmp_23, mux_tmp_318, nor_143_nl);
  assign nor_142_nl = ~(Gelu_for_9_else_slc_32_svs | (~ Gelu_for_9_slc_32_1_svs));
  assign mux_336_nl = MUX_s_1_2_2(mux_335_nl, mux_tmp_317, nor_142_nl);
  assign mux_339_nl = MUX_s_1_2_2(mux_338_nl, mux_336_nl, act_config_in_InstFetch_return_sva_7_2[2]);
  assign mux_340_nl = MUX_s_1_2_2(nand_tmp_23, mux_339_nl, and_1648_cse);
  assign and_899_rmff = (~ mux_340_nl) & and_dcpl_856;
  assign or_877_nl = (~ Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)
      | Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign mux_347_nl = MUX_s_1_2_2(mux_tmp_328, nand_tmp_25, or_877_nl);
  assign or_876_nl = (~ Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)
      | Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign mux_348_nl = MUX_s_1_2_2(mux_tmp_327, mux_347_nl, or_876_nl);
  assign nor_147_nl = ~(Gelu_for_3_else_slc_32_svs | (~ Gelu_for_3_slc_32_1_svs));
  assign mux_345_nl = MUX_s_1_2_2(nand_tmp_25, mux_tmp_328, nor_147_nl);
  assign nor_146_nl = ~(Gelu_for_10_else_slc_32_svs | (~ Gelu_for_10_slc_32_1_svs));
  assign mux_346_nl = MUX_s_1_2_2(mux_345_nl, mux_tmp_327, nor_146_nl);
  assign mux_349_nl = MUX_s_1_2_2(mux_348_nl, mux_346_nl, act_config_in_InstFetch_return_sva_7_2[2]);
  assign mux_350_nl = MUX_s_1_2_2(nand_tmp_25, mux_349_nl, and_1648_cse);
  assign and_900_rmff = (~ mux_350_nl) & and_dcpl_856;
  assign or_882_nl = (~ Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)
      | Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign mux_357_nl = MUX_s_1_2_2(mux_tmp_338, nand_tmp_27, or_882_nl);
  assign or_881_nl = (~ Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)
      | Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign mux_358_nl = MUX_s_1_2_2(mux_tmp_337, mux_357_nl, or_881_nl);
  assign nor_151_nl = ~(Gelu_for_4_else_slc_32_svs | (~ Gelu_for_4_slc_32_1_svs));
  assign mux_355_nl = MUX_s_1_2_2(nand_tmp_27, mux_tmp_338, nor_151_nl);
  assign nor_150_nl = ~(Gelu_for_11_else_slc_32_svs | (~ Gelu_for_11_slc_32_1_svs));
  assign mux_356_nl = MUX_s_1_2_2(mux_355_nl, mux_tmp_337, nor_150_nl);
  assign mux_359_nl = MUX_s_1_2_2(mux_358_nl, mux_356_nl, act_config_in_InstFetch_return_sva_7_2[2]);
  assign mux_360_nl = MUX_s_1_2_2(nand_tmp_27, mux_359_nl, and_1648_cse);
  assign and_901_rmff = (~ mux_360_nl) & and_dcpl_856;
  assign or_887_nl = (~ Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)
      | Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign mux_367_nl = MUX_s_1_2_2(mux_tmp_348, nand_tmp_29, or_887_nl);
  assign or_886_nl = (~ Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)
      | Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign mux_368_nl = MUX_s_1_2_2(mux_tmp_347, mux_367_nl, or_886_nl);
  assign nor_155_nl = ~(Gelu_for_5_else_slc_32_svs | (~ Gelu_for_5_slc_32_1_svs));
  assign mux_365_nl = MUX_s_1_2_2(nand_tmp_29, mux_tmp_348, nor_155_nl);
  assign nor_154_nl = ~(Gelu_for_12_else_slc_32_svs | (~ Gelu_for_12_slc_32_1_svs));
  assign mux_366_nl = MUX_s_1_2_2(mux_365_nl, mux_tmp_347, nor_154_nl);
  assign mux_369_nl = MUX_s_1_2_2(mux_368_nl, mux_366_nl, act_config_in_InstFetch_return_sva_7_2[2]);
  assign mux_370_nl = MUX_s_1_2_2(nand_tmp_29, mux_369_nl, and_1648_cse);
  assign and_902_rmff = (~ mux_370_nl) & and_dcpl_856;
  assign or_892_nl = (~ Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)
      | Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign mux_377_nl = MUX_s_1_2_2(mux_tmp_358, nand_tmp_31, or_892_nl);
  assign or_891_nl = (~ Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)
      | Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign mux_378_nl = MUX_s_1_2_2(mux_tmp_357, mux_377_nl, or_891_nl);
  assign nor_159_nl = ~(Gelu_for_6_else_slc_32_svs | (~ Gelu_for_6_slc_32_1_svs));
  assign mux_375_nl = MUX_s_1_2_2(nand_tmp_31, mux_tmp_358, nor_159_nl);
  assign nor_158_nl = ~(Gelu_for_13_else_slc_32_svs | (~ Gelu_for_13_slc_32_1_svs));
  assign mux_376_nl = MUX_s_1_2_2(mux_375_nl, mux_tmp_357, nor_158_nl);
  assign mux_379_nl = MUX_s_1_2_2(mux_378_nl, mux_376_nl, act_config_in_InstFetch_return_sva_7_2[2]);
  assign mux_380_nl = MUX_s_1_2_2(nand_tmp_31, mux_379_nl, and_1648_cse);
  assign and_903_rmff = (~ mux_380_nl) & and_dcpl_856;
  assign or_897_nl = (~ Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)
      | Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign mux_387_nl = MUX_s_1_2_2(mux_tmp_368, nand_tmp_33, or_897_nl);
  assign or_896_nl = (~ Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)
      | Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign mux_388_nl = MUX_s_1_2_2(mux_tmp_367, mux_387_nl, or_896_nl);
  assign nor_163_nl = ~(Gelu_for_7_else_slc_32_svs | (~ Gelu_for_7_slc_32_1_svs));
  assign mux_385_nl = MUX_s_1_2_2(nand_tmp_33, mux_tmp_368, nor_163_nl);
  assign nor_162_nl = ~(Gelu_for_14_else_slc_32_svs | (~ Gelu_for_14_slc_32_1_svs));
  assign mux_386_nl = MUX_s_1_2_2(mux_385_nl, mux_tmp_367, nor_162_nl);
  assign mux_389_nl = MUX_s_1_2_2(mux_388_nl, mux_386_nl, act_config_in_InstFetch_return_sva_7_2[2]);
  assign mux_390_nl = MUX_s_1_2_2(nand_tmp_33, mux_389_nl, and_1648_cse);
  assign and_904_rmff = (~ mux_390_nl) & and_dcpl_856;
  assign or_902_nl = (~ Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)
      | Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign mux_397_nl = MUX_s_1_2_2(mux_tmp_378, nand_tmp_35, or_902_nl);
  assign or_901_nl = (~ Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)
      | Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign mux_398_nl = MUX_s_1_2_2(mux_tmp_377, mux_397_nl, or_901_nl);
  assign nor_167_nl = ~(Gelu_for_8_else_slc_32_svs | (~ Gelu_for_8_slc_32_1_svs));
  assign mux_395_nl = MUX_s_1_2_2(nand_tmp_35, mux_tmp_378, nor_167_nl);
  assign nor_166_nl = ~(Gelu_for_15_else_slc_32_svs | (~ Gelu_for_15_slc_32_1_svs));
  assign mux_396_nl = MUX_s_1_2_2(mux_395_nl, mux_tmp_377, nor_166_nl);
  assign mux_399_nl = MUX_s_1_2_2(mux_398_nl, mux_396_nl, act_config_in_InstFetch_return_sva_7_2[2]);
  assign mux_400_nl = MUX_s_1_2_2(nand_tmp_35, mux_399_nl, and_1648_cse);
  assign and_905_rmff = (~ mux_400_nl) & and_dcpl_856;
  assign or_907_nl = (~ Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)
      | Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign mux_407_nl = MUX_s_1_2_2(mux_tmp_388, nand_tmp_37, or_907_nl);
  assign or_906_nl = (~ Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)
      | Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign mux_408_nl = MUX_s_1_2_2(mux_tmp_387, mux_407_nl, or_906_nl);
  assign nor_171_nl = ~(Gelu_for_2_else_slc_32_svs | (~ Gelu_for_2_slc_32_1_svs));
  assign mux_405_nl = MUX_s_1_2_2(nand_tmp_37, mux_tmp_388, nor_171_nl);
  assign nor_170_nl = ~(Gelu_for_16_else_slc_32_svs | (~ Gelu_for_16_slc_32_1_svs));
  assign mux_406_nl = MUX_s_1_2_2(mux_405_nl, mux_tmp_387, nor_170_nl);
  assign mux_409_nl = MUX_s_1_2_2(mux_408_nl, mux_406_nl, act_config_in_InstFetch_return_sva_7_2[2]);
  assign mux_410_nl = MUX_s_1_2_2(nand_tmp_37, mux_409_nl, and_1648_cse);
  assign and_906_rmff = (~ mux_410_nl) & and_dcpl_856;
  assign and_915_rmff = and_dcpl_872 & and_dcpl_867 & Gelu_for_2_slc_32_1_svs & Gelu_for_2_else_slc_32_svs
      & (~ Gelu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs)
      & (~ (fsm_output[3]));
  assign and_920_rmff = and_dcpl_872 & and_dcpl_867 & Gelu_for_3_slc_32_1_svs & Gelu_for_3_else_slc_32_svs
      & (~ Gelu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs)
      & (~ (fsm_output[3]));
  assign and_925_rmff = and_dcpl_872 & and_dcpl_867 & Gelu_for_4_slc_32_1_svs & Gelu_for_4_else_slc_32_svs
      & (~ Gelu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs)
      & (~ (fsm_output[3]));
  assign and_930_rmff = and_dcpl_872 & and_dcpl_867 & Gelu_for_5_slc_32_1_svs & Gelu_for_5_else_slc_32_svs
      & (~ Gelu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs)
      & (~ (fsm_output[3]));
  assign and_935_rmff = and_dcpl_872 & and_dcpl_867 & Gelu_for_6_slc_32_1_svs & Gelu_for_6_else_slc_32_svs
      & (~ Gelu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs)
      & (~ (fsm_output[3]));
  assign and_940_rmff = and_dcpl_872 & and_dcpl_867 & Gelu_for_7_slc_32_1_svs & Gelu_for_7_else_slc_32_svs
      & (~ Gelu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs)
      & (~ (fsm_output[3]));
  assign and_945_rmff = and_dcpl_872 & and_dcpl_867 & Gelu_for_8_slc_32_1_svs & Gelu_for_8_else_slc_32_svs
      & (~ Gelu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs)
      & (~ (fsm_output[3]));
  assign and_950_rmff = and_dcpl_872 & and_dcpl_867 & Gelu_for_9_slc_32_1_svs & Gelu_for_9_else_slc_32_svs
      & (~ Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & (~ (fsm_output[3]));
  assign and_955_rmff = and_dcpl_872 & and_dcpl_867 & Gelu_for_10_slc_32_1_svs &
      Gelu_for_10_else_slc_32_svs & (~ Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & (~ (fsm_output[3]));
  assign and_960_rmff = and_dcpl_872 & and_dcpl_867 & Gelu_for_11_slc_32_1_svs &
      Gelu_for_11_else_slc_32_svs & (~ Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & (~ (fsm_output[3]));
  assign and_965_rmff = and_dcpl_872 & and_dcpl_867 & Gelu_for_12_slc_32_1_svs &
      Gelu_for_12_else_slc_32_svs & (~ Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & (~ (fsm_output[3]));
  assign and_970_rmff = and_dcpl_872 & and_dcpl_867 & Gelu_for_13_slc_32_1_svs &
      Gelu_for_13_else_slc_32_svs & (~ Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & (~ (fsm_output[3]));
  assign and_975_rmff = and_dcpl_872 & and_dcpl_867 & Gelu_for_14_slc_32_1_svs &
      Gelu_for_14_else_slc_32_svs & (~ Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & (~ (fsm_output[3]));
  assign and_980_rmff = and_dcpl_872 & and_dcpl_867 & Gelu_for_15_slc_32_1_svs &
      Gelu_for_15_else_slc_32_svs & (~ Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & (~ (fsm_output[3]));
  assign and_985_rmff = and_dcpl_872 & and_dcpl_867 & Gelu_for_16_slc_32_1_svs &
      Gelu_for_16_else_slc_32_svs & (~ Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & (~ (fsm_output[3]));
  assign and_990_rmff = and_dcpl_872 & and_dcpl_867 & Gelu_for_1_slc_32_1_svs & Gelu_for_1_else_slc_32_svs
      & (~ Gelu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs)
      & (~ (fsm_output[3]));
  assign mux_rmff = MUX_v_3_2_2(3'b011, 3'b100, operator_32_8_true_AC_TRN_AC_WRAP_6_less_14_tmp);
  assign and_1658_nl = (~(operator_32_8_true_AC_TRN_AC_WRAP_6_less_14_tmp & operator_32_8_true_AC_TRN_AC_WRAP_7_less_14_tmp))
      & and_2371_cse;
  assign nor_431_nl = ~((Gelu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      | (fsm_output[1:0]!=2'b00));
  assign mux_412_nl = MUX_s_1_2_2(and_1658_nl, nor_431_nl, fsm_output[2]);
  assign and_998_rmff = mux_412_nl & (act_config_in_InstFetch_return_sva_7_2[4])
      & and_dcpl_953 & Gelu_for_2_slc_32_1_svs & Gelu_for_2_else_slc_32_svs & Gelu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
      & (~ (fsm_output[3]));
  assign mux_1_rmff = MUX_v_3_2_2(3'b011, 3'b100, operator_32_8_true_AC_TRN_AC_WRAP_6_less_13_tmp);
  assign and_1661_nl = (~(operator_32_8_true_AC_TRN_AC_WRAP_6_less_13_tmp & operator_32_8_true_AC_TRN_AC_WRAP_7_less_13_tmp))
      & and_2371_cse;
  assign nor_432_nl = ~((Gelu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      | (fsm_output[1:0]!=2'b00));
  assign mux_413_nl = MUX_s_1_2_2(and_1661_nl, nor_432_nl, fsm_output[2]);
  assign and_1004_rmff = mux_413_nl & (act_config_in_InstFetch_return_sva_7_2[4])
      & and_dcpl_953 & Gelu_for_3_slc_32_1_svs & Gelu_for_3_else_slc_32_svs & Gelu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
      & (~ (fsm_output[3]));
  assign mux_2_rmff = MUX_v_3_2_2(3'b011, 3'b100, operator_32_8_true_AC_TRN_AC_WRAP_6_less_12_tmp);
  assign and_1664_nl = (~(operator_32_8_true_AC_TRN_AC_WRAP_6_less_12_tmp & operator_32_8_true_AC_TRN_AC_WRAP_7_less_12_tmp))
      & and_2371_cse;
  assign nor_433_nl = ~((Gelu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      | (fsm_output[1:0]!=2'b00));
  assign mux_414_nl = MUX_s_1_2_2(and_1664_nl, nor_433_nl, fsm_output[2]);
  assign and_1010_rmff = mux_414_nl & (act_config_in_InstFetch_return_sva_7_2[4])
      & and_dcpl_953 & Gelu_for_4_slc_32_1_svs & Gelu_for_4_else_slc_32_svs & Gelu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
      & (~ (fsm_output[3]));
  assign mux_3_rmff = MUX_v_3_2_2(3'b011, 3'b100, operator_32_8_true_AC_TRN_AC_WRAP_6_less_11_tmp);
  assign and_1667_nl = (~(operator_32_8_true_AC_TRN_AC_WRAP_6_less_11_tmp & operator_32_8_true_AC_TRN_AC_WRAP_7_less_11_tmp))
      & and_2371_cse;
  assign nor_434_nl = ~((Gelu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      | (fsm_output[1:0]!=2'b00));
  assign mux_415_nl = MUX_s_1_2_2(and_1667_nl, nor_434_nl, fsm_output[2]);
  assign and_1016_rmff = mux_415_nl & (act_config_in_InstFetch_return_sva_7_2[4])
      & and_dcpl_953 & Gelu_for_5_slc_32_1_svs & Gelu_for_5_else_slc_32_svs & Gelu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
      & (~ (fsm_output[3]));
  assign mux_4_rmff = MUX_v_3_2_2(3'b011, 3'b100, operator_32_8_true_AC_TRN_AC_WRAP_6_less_10_tmp);
  assign and_1670_nl = (~(operator_32_8_true_AC_TRN_AC_WRAP_6_less_10_tmp & operator_32_8_true_AC_TRN_AC_WRAP_7_less_10_tmp))
      & and_2371_cse;
  assign nor_435_nl = ~((Gelu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      | (fsm_output[1:0]!=2'b00));
  assign mux_416_nl = MUX_s_1_2_2(and_1670_nl, nor_435_nl, fsm_output[2]);
  assign and_1022_rmff = mux_416_nl & (act_config_in_InstFetch_return_sva_7_2[4])
      & and_dcpl_953 & Gelu_for_6_slc_32_1_svs & Gelu_for_6_else_slc_32_svs & Gelu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
      & (~ (fsm_output[3]));
  assign mux_5_rmff = MUX_v_3_2_2(3'b011, 3'b100, operator_32_8_true_AC_TRN_AC_WRAP_6_less_9_tmp);
  assign and_1673_nl = (~(operator_32_8_true_AC_TRN_AC_WRAP_6_less_9_tmp & operator_32_8_true_AC_TRN_AC_WRAP_7_less_9_tmp))
      & and_2371_cse;
  assign nor_436_nl = ~((Gelu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      | (fsm_output[1:0]!=2'b00));
  assign mux_417_nl = MUX_s_1_2_2(and_1673_nl, nor_436_nl, fsm_output[2]);
  assign and_1028_rmff = mux_417_nl & (act_config_in_InstFetch_return_sva_7_2[4])
      & and_dcpl_953 & Gelu_for_7_slc_32_1_svs & Gelu_for_7_else_slc_32_svs & Gelu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
      & (~ (fsm_output[3]));
  assign mux_6_rmff = MUX_v_3_2_2(3'b011, 3'b100, operator_32_8_true_AC_TRN_AC_WRAP_6_less_8_tmp);
  assign and_1676_nl = (~(operator_32_8_true_AC_TRN_AC_WRAP_6_less_8_tmp & operator_32_8_true_AC_TRN_AC_WRAP_7_less_8_tmp))
      & and_2371_cse;
  assign nor_437_nl = ~((Gelu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      | (fsm_output[1:0]!=2'b00));
  assign mux_418_nl = MUX_s_1_2_2(and_1676_nl, nor_437_nl, fsm_output[2]);
  assign and_1034_rmff = mux_418_nl & (act_config_in_InstFetch_return_sva_7_2[4])
      & and_dcpl_953 & Gelu_for_8_slc_32_1_svs & Gelu_for_8_else_slc_32_svs & Gelu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
      & (~ (fsm_output[3]));
  assign mux_7_rmff = MUX_v_3_2_2(3'b011, 3'b100, operator_32_8_true_AC_TRN_AC_WRAP_6_less_7_tmp);
  assign and_1679_nl = (~(operator_32_8_true_AC_TRN_AC_WRAP_6_less_7_tmp & operator_32_8_true_AC_TRN_AC_WRAP_7_less_7_tmp))
      & and_2371_cse;
  assign nor_438_nl = ~((Gelu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      | (fsm_output[1:0]!=2'b00));
  assign mux_419_nl = MUX_s_1_2_2(and_1679_nl, nor_438_nl, fsm_output[2]);
  assign and_1040_rmff = mux_419_nl & (act_config_in_InstFetch_return_sva_7_2[4])
      & and_dcpl_953 & Gelu_for_9_slc_32_1_svs & Gelu_for_9_else_slc_32_svs & Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & (~ (fsm_output[3]));
  assign mux_8_rmff = MUX_v_3_2_2(3'b011, 3'b100, operator_32_8_true_AC_TRN_AC_WRAP_6_less_6_tmp);
  assign and_1682_nl = (~(operator_32_8_true_AC_TRN_AC_WRAP_6_less_6_tmp & operator_32_8_true_AC_TRN_AC_WRAP_7_less_6_tmp))
      & and_2371_cse;
  assign nor_439_nl = ~((Gelu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      | (fsm_output[1:0]!=2'b00));
  assign mux_420_nl = MUX_s_1_2_2(and_1682_nl, nor_439_nl, fsm_output[2]);
  assign and_1046_rmff = mux_420_nl & (act_config_in_InstFetch_return_sva_7_2[4])
      & and_dcpl_953 & Gelu_for_10_slc_32_1_svs & Gelu_for_10_else_slc_32_svs & Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & (~ (fsm_output[3]));
  assign mux_9_rmff = MUX_v_3_2_2(3'b011, 3'b100, operator_32_8_true_AC_TRN_AC_WRAP_6_less_5_tmp);
  assign and_1685_nl = (~(operator_32_8_true_AC_TRN_AC_WRAP_6_less_5_tmp & operator_32_8_true_AC_TRN_AC_WRAP_7_less_5_tmp))
      & and_2371_cse;
  assign nor_440_nl = ~((Gelu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      | (fsm_output[1:0]!=2'b00));
  assign mux_421_nl = MUX_s_1_2_2(and_1685_nl, nor_440_nl, fsm_output[2]);
  assign and_1052_rmff = mux_421_nl & (act_config_in_InstFetch_return_sva_7_2[4])
      & and_dcpl_953 & Gelu_for_11_slc_32_1_svs & Gelu_for_11_else_slc_32_svs & Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & (~ (fsm_output[3]));
  assign mux_10_rmff = MUX_v_3_2_2(3'b011, 3'b100, operator_32_8_true_AC_TRN_AC_WRAP_6_less_4_tmp);
  assign and_1688_nl = (~(operator_32_8_true_AC_TRN_AC_WRAP_6_less_4_tmp & operator_32_8_true_AC_TRN_AC_WRAP_7_less_4_tmp))
      & and_2371_cse;
  assign nor_441_nl = ~((Gelu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      | (fsm_output[1:0]!=2'b00));
  assign mux_422_nl = MUX_s_1_2_2(and_1688_nl, nor_441_nl, fsm_output[2]);
  assign and_1058_rmff = mux_422_nl & (act_config_in_InstFetch_return_sva_7_2[4])
      & and_dcpl_953 & Gelu_for_12_slc_32_1_svs & Gelu_for_12_else_slc_32_svs & Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & (~ (fsm_output[3]));
  assign mux_11_rmff = MUX_v_3_2_2(3'b011, 3'b100, operator_32_8_true_AC_TRN_AC_WRAP_6_less_3_tmp);
  assign and_1691_nl = (~(operator_32_8_true_AC_TRN_AC_WRAP_6_less_3_tmp & operator_32_8_true_AC_TRN_AC_WRAP_7_less_3_tmp))
      & and_2371_cse;
  assign nor_442_nl = ~((Gelu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      | (fsm_output[1:0]!=2'b00));
  assign mux_423_nl = MUX_s_1_2_2(and_1691_nl, nor_442_nl, fsm_output[2]);
  assign and_1064_rmff = mux_423_nl & (act_config_in_InstFetch_return_sva_7_2[4])
      & and_dcpl_953 & Gelu_for_13_slc_32_1_svs & Gelu_for_13_else_slc_32_svs & Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & (~ (fsm_output[3]));
  assign mux_12_rmff = MUX_v_3_2_2(3'b011, 3'b100, operator_32_8_true_AC_TRN_AC_WRAP_6_less_2_tmp);
  assign and_1694_nl = (~(operator_32_8_true_AC_TRN_AC_WRAP_6_less_2_tmp & operator_32_8_true_AC_TRN_AC_WRAP_7_less_2_tmp))
      & and_2371_cse;
  assign nor_443_nl = ~((Gelu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      | (fsm_output[1:0]!=2'b00));
  assign mux_424_nl = MUX_s_1_2_2(and_1694_nl, nor_443_nl, fsm_output[2]);
  assign and_1070_rmff = mux_424_nl & (act_config_in_InstFetch_return_sva_7_2[4])
      & and_dcpl_953 & Gelu_for_14_slc_32_1_svs & Gelu_for_14_else_slc_32_svs & Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & (~ (fsm_output[3]));
  assign mux_13_rmff = MUX_v_3_2_2(3'b011, 3'b100, operator_32_8_true_AC_TRN_AC_WRAP_6_less_1_tmp);
  assign and_1697_nl = (~(operator_32_8_true_AC_TRN_AC_WRAP_6_less_1_tmp & operator_32_8_true_AC_TRN_AC_WRAP_7_less_1_tmp))
      & and_2371_cse;
  assign nor_444_nl = ~((Gelu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      | (fsm_output[1:0]!=2'b00));
  assign mux_425_nl = MUX_s_1_2_2(and_1697_nl, nor_444_nl, fsm_output[2]);
  assign and_1076_rmff = mux_425_nl & (act_config_in_InstFetch_return_sva_7_2[4])
      & and_dcpl_953 & Gelu_for_15_slc_32_1_svs & Gelu_for_15_else_slc_32_svs & Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & (~ (fsm_output[3]));
  assign mux_14_rmff = MUX_v_3_2_2(3'b011, 3'b100, operator_32_8_true_AC_TRN_AC_WRAP_6_less_tmp);
  assign and_1701_nl = (fsm_output[1]) & (~(operator_32_8_true_AC_TRN_AC_WRAP_6_less_tmp
      & operator_32_8_true_AC_TRN_AC_WRAP_7_less_tmp)) & (fsm_output[0]);
  assign nor_445_nl = ~((fsm_output[1]) | (Gelu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      | (fsm_output[0]));
  assign mux_426_nl = MUX_s_1_2_2(and_1701_nl, nor_445_nl, fsm_output[2]);
  assign and_1082_rmff = mux_426_nl & (act_config_in_InstFetch_return_sva_7_2[4])
      & and_dcpl_953 & Gelu_for_16_slc_32_1_svs & Gelu_for_16_else_slc_32_svs & Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & (~ (fsm_output[3]));
  assign mux_15_rmff = MUX_v_3_2_2(3'b011, 3'b100, operator_32_8_true_AC_TRN_AC_WRAP_6_less_15_tmp);
  assign and_1704_nl = (~(operator_32_8_true_AC_TRN_AC_WRAP_6_less_15_tmp & operator_32_8_true_AC_TRN_AC_WRAP_7_less_15_tmp))
      & and_2371_cse;
  assign nor_446_nl = ~((Gelu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      | (fsm_output[1:0]!=2'b00));
  assign mux_427_nl = MUX_s_1_2_2(and_1704_nl, nor_446_nl, fsm_output[2]);
  assign and_1088_rmff = mux_427_nl & (act_config_in_InstFetch_return_sva_7_2[4])
      & and_dcpl_953 & Gelu_for_1_slc_32_1_svs & Gelu_for_1_else_slc_32_svs & Gelu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
      & (~ (fsm_output[3]));
  assign and_1097_rmff = nor_447_cse & act_config_InstIncr_if_equal_1_tmp & and_dcpl_1051
      & and_dcpl_1048 & (fsm_output[3]) & act_config_InstIncr_if_act_config_InstIncr_if_if_nor_tmp
      & is_incr_lpi_1_dfm_1;
  assign and_1102_rmff = and_dcpl_469 & (fsm_output[0]) & and_dcpl_1056 & (~ (fsm_output[3]));
  assign and_1106_rmff = and_dcpl_1063 & and_dcpl_1061;
  assign and_1108_rmff = and_dcpl_1063 & and_dcpl_1061 & w_axi_rsp_lpi_1_dfm_1;
  assign and_1113_rmff = (act_config_in_InstFetch_mux_tmp[7:4]==4'b0011) & is_start_sva
      & and_dcpl_847;
  assign and_1116_rmff = and_dcpl_1072 & (~ (fsm_output[1])) & nor_1441_cse;
  assign nor_223_nl = ~((~ (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[8])
      | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[10]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[9])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]));
  assign or_359_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[8])
      | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[10]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[9])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]);
  assign mux_102_nl = MUX_s_1_2_2(nor_223_nl, or_359_nl, act_config_is_valid_sva);
  assign nor_42_nl = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1:0]!=2'b01));
  assign mux_103_nl = MUX_s_1_2_2(act_config_is_valid_sva, mux_102_nl, nor_42_nl);
  assign ActUnit_DecodeAxi_if_and_37_cse = ActUnitRun_wen & and_dcpl_331 & (mux_103_nl
      | is_start_sva);
  assign and_1521_nl = ActUnit_CheckStart_start_reg_sva & act_config_is_valid_sva;
  assign mux_319_nl = MUX_s_1_2_2(is_start_sva, or_dcpl_28, and_1521_nl);
  assign or_695_nl = (z_out[4]) | act_config_is_zero_first_sva | (~ and_dcpl_333);
  assign or_656_nl = act_config_is_zero_first_sva | (~ and_dcpl_333);
  assign mux_314_nl = MUX_s_1_2_2(or_tmp_397, (~ or_dcpl_28), w_load_lpi_1_dfm_1);
  assign mux_315_nl = MUX_s_1_2_2(mux_314_nl, or_tmp_397, act_config_is_zero_first_sva);
  assign mux_316_nl = MUX_s_1_2_2(or_656_nl, mux_315_nl, act_config_is_valid_sva);
  assign or_692_nl = (~ act_config_is_valid_sva) | is_start_sva | (~ ActUnit_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva);
  assign mux_317_nl = MUX_s_1_2_2(mux_316_nl, or_692_nl, z_out[4]);
  assign mux_318_nl = MUX_s_1_2_2(or_695_nl, mux_317_nl, ActUnit_CheckStart_start_reg_sva);
  assign mux_320_nl = MUX_s_1_2_2((~ mux_319_nl), mux_318_nl, is_incr_lpi_1_dfm_1);
  assign act_config_inst_regs_and_36_cse = ActUnitRun_wen & and_dcpl_1090 & mux_320_nl;
  assign act_config_num_inst_and_cse = ActUnitRun_wen & (~(or_dcpl_485 | or_dcpl_475
      | or_dcpl_457 | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1:0]!=2'b01)));
  assign rva_out_reg_data_and_ssc = ActUnitRun_wen & ((~ mux_tmp_413) | and_dcpl_1094
      | and_dcpl_1096);
  assign or_1427_cse = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0!=4'b0000);
  assign or_1527_tmp = and_dcpl_1426 | mux_tmp_413;
  assign nor_1405_cse = ~((fsm_output[2:0]!=3'b010));
  assign or_3395_cse = (fsm_output[2:1]!=2'b00);
  assign and_1720_cse = and_dcpl_1236 & (~ or_dcpl_1012);
  assign nor_1406_cse = ~((ActUnit_PushOutput_if_for_i_4_0_sva_3_0!=4'b0001));
  assign act_mem_banks_bank_a_and_cse = ActUnitRun_wen & (~(or_dcpl_498 | or_dcpl_496
      | or_dcpl_494));
  assign act_mem_banks_bank_a_and_1_cse = ActUnitRun_wen & (~(or_dcpl_498 | or_dcpl_496
      | or_dcpl_501));
  assign act_mem_banks_bank_a_and_2_cse = ActUnitRun_wen & (~(or_dcpl_498 | or_dcpl_496
      | or_dcpl_505));
  assign act_mem_banks_bank_a_and_3_cse = ActUnitRun_wen & (~(or_dcpl_498 | or_dcpl_496
      | or_dcpl_509));
  assign act_mem_banks_bank_a_and_4_cse = ActUnitRun_wen & (~(or_dcpl_498 | or_dcpl_496
      | or_dcpl_513));
  assign act_mem_banks_bank_a_and_5_cse = ActUnitRun_wen & (~(or_dcpl_498 | or_dcpl_496
      | or_dcpl_516));
  assign act_mem_banks_bank_a_and_6_cse = ActUnitRun_wen & (~(or_dcpl_498 | or_dcpl_496
      | or_dcpl_519));
  assign act_mem_banks_bank_a_and_7_cse = ActUnitRun_wen & (~(or_dcpl_498 | or_dcpl_496
      | or_dcpl_522));
  assign act_mem_banks_bank_a_and_8_cse = ActUnitRun_wen & (~(or_dcpl_498 | or_dcpl_496
      | or_dcpl_526));
  assign act_mem_banks_bank_a_and_9_cse = ActUnitRun_wen & (~(or_dcpl_498 | or_dcpl_496
      | or_dcpl_529));
  assign act_mem_banks_bank_a_and_10_cse = ActUnitRun_wen & (~(or_dcpl_498 | or_dcpl_496
      | or_dcpl_532));
  assign act_mem_banks_bank_a_and_11_cse = ActUnitRun_wen & (~(or_dcpl_498 | or_dcpl_496
      | or_dcpl_535));
  assign act_mem_banks_bank_a_and_12_cse = ActUnitRun_wen & (~(or_dcpl_498 | or_dcpl_496
      | or_dcpl_539));
  assign act_mem_banks_bank_a_and_13_cse = ActUnitRun_wen & (~(or_dcpl_498 | or_dcpl_496
      | or_dcpl_542));
  assign act_mem_banks_bank_a_and_14_cse = ActUnitRun_wen & (~(or_dcpl_498 | or_dcpl_496
      | or_dcpl_545));
  assign act_mem_banks_bank_a_and_15_cse = ActUnitRun_wen & (~(or_dcpl_498 | or_dcpl_496
      | or_dcpl_548));
  assign act_mem_banks_bank_a_and_16_cse = ActUnitRun_wen & (~(or_dcpl_498 | or_dcpl_552
      | or_dcpl_494));
  assign act_mem_banks_bank_a_and_17_cse = ActUnitRun_wen & (~(or_dcpl_498 | or_dcpl_552
      | or_dcpl_501));
  assign act_mem_banks_bank_a_and_18_cse = ActUnitRun_wen & (~(or_dcpl_498 | or_dcpl_552
      | or_dcpl_505));
  assign act_mem_banks_bank_a_and_19_cse = ActUnitRun_wen & (~(or_dcpl_498 | or_dcpl_552
      | or_dcpl_509));
  assign act_mem_banks_bank_a_and_20_cse = ActUnitRun_wen & (~(or_dcpl_498 | or_dcpl_552
      | or_dcpl_513));
  assign act_mem_banks_bank_a_and_21_cse = ActUnitRun_wen & (~(or_dcpl_498 | or_dcpl_552
      | or_dcpl_516));
  assign act_mem_banks_bank_a_and_22_cse = ActUnitRun_wen & (~(or_dcpl_498 | or_dcpl_552
      | or_dcpl_519));
  assign act_mem_banks_bank_a_and_23_cse = ActUnitRun_wen & (~(or_dcpl_498 | or_dcpl_552
      | or_dcpl_522));
  assign act_mem_banks_bank_a_and_24_cse = ActUnitRun_wen & (~(or_dcpl_498 | or_dcpl_552
      | or_dcpl_526));
  assign act_mem_banks_bank_a_and_25_cse = ActUnitRun_wen & (~(or_dcpl_498 | or_dcpl_552
      | or_dcpl_529));
  assign act_mem_banks_bank_a_and_26_cse = ActUnitRun_wen & (~(or_dcpl_498 | or_dcpl_552
      | or_dcpl_532));
  assign act_mem_banks_bank_a_and_27_cse = ActUnitRun_wen & (~(or_dcpl_498 | or_dcpl_552
      | or_dcpl_535));
  assign act_mem_banks_bank_a_and_28_cse = ActUnitRun_wen & (~(or_dcpl_498 | or_dcpl_552
      | or_dcpl_539));
  assign act_mem_banks_bank_a_and_29_cse = ActUnitRun_wen & (~(or_dcpl_498 | or_dcpl_552
      | or_dcpl_542));
  assign act_mem_banks_bank_a_and_30_cse = ActUnitRun_wen & (~(or_dcpl_498 | or_dcpl_552
      | or_dcpl_545));
  assign act_mem_banks_bank_a_and_31_cse = ActUnitRun_wen & (~(or_dcpl_498 | or_dcpl_552
      | or_dcpl_548));
  assign act_config_inst_regs_and_4_cse = ActUnitRun_wen & (~(or_dcpl_586 | (fsm_output[3])
      | not_tmp_503));
  assign act_config_inst_regs_and_20_cse = ActUnitRun_wen & (~(or_dcpl_485 | or_dcpl_475
      | or_dcpl_457 | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1:0]!=2'b10)));
  assign nl_operator_8_false_acc_sdt = ({reg_act_config_output_counter_sva_dfm_3_ftd
      , reg_act_config_output_counter_sva_dfm_3_ftd_1_3 , reg_act_config_output_counter_sva_dfm_3_ftd_1_2_0})
      + 8'b00000001;
  assign operator_8_false_acc_sdt = nl_operator_8_false_acc_sdt[7:0];
  assign act_config_output_counter_and_ssc = ActUnitRun_wen & (act_config_output_counter_sva_mx0c0
      | act_config_output_counter_sva_mx0c1 | act_config_output_counter_sva_mx0c2);
  assign nl_Silu_for_11_else_else_else_else_if_acc_sdt = ({reg_nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1})
      + 4'b1111;
  assign Silu_for_11_else_else_else_else_if_acc_sdt = nl_Silu_for_11_else_else_else_else_if_acc_sdt[3:0];
  assign act_config_output_counter_and_3_ssc = (~ and_dcpl_1235) & act_config_output_counter_sva_mx0c0;
  assign act_config_output_counter_and_2_ssc = act_config_output_counter_and_ssc
      & (~ and_dcpl_1112);
  assign act_regs_data_and_ssc = ActUnitRun_wen & and_dcpl_1104;
  assign act_regs_data_and_2530_enex5 = act_regs_data_and_ssc & (reg_act_config_is_zero_first_sva_dfm_4_enexo
      | reg_act_regs_data_2_2_sva_8_30_26_enexo | reg_w_load_lpi_1_dfm_1_enexo |
      reg_is_start_enexo | reg_act_regs_data_3_15_sva_8_30_26_enexo | reg_act_regs_data_3_15_sva_dfm_2_30_26_enexo);
  assign act_regs_data_and_2531_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_2_2_sva_8_25_22_enexo
      | reg_is_start_enexo_1 | reg_act_regs_data_3_15_sva_8_25_22_enexo | reg_w_load_lpi_1_dfm_1_enexo_1
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_1 | reg_act_regs_data_3_15_sva_dfm_2_25_22_enexo);
  assign act_regs_data_and_2532_enex5 = act_regs_data_and_ssc & (reg_w_load_lpi_1_dfm_1_enexo_2
      | reg_is_start_enexo_2 | reg_act_regs_data_3_15_sva_8_21_0_enexo | reg_act_regs_data_3_15_sva_dfm_2_21_0_enexo
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_2 | reg_act_regs_data_2_2_sva_8_21_0_enexo);
  assign act_regs_data_and_2533_enex5 = act_regs_data_and_ssc & (reg_act_config_is_zero_first_sva_dfm_4_enexo_3
      | reg_act_regs_data_3_14_sva_8_30_26_enexo | reg_act_regs_data_3_14_sva_dfm_2_30_26_enexo
      | reg_w_load_lpi_1_dfm_1_enexo_3 | reg_act_regs_data_2_15_sva_8_30_26_enexo
      | reg_is_start_enexo_3);
  assign act_regs_data_and_2534_enex5 = act_regs_data_and_ssc & (reg_w_load_lpi_1_dfm_1_enexo_4
      | reg_act_regs_data_3_14_sva_8_25_22_enexo | reg_act_config_is_zero_first_sva_dfm_4_enexo_4
      | reg_act_regs_data_3_14_sva_dfm_2_25_22_enexo | reg_act_regs_data_2_15_sva_8_25_22_enexo
      | reg_is_start_enexo_4);
  assign act_regs_data_and_2535_enex5 = act_regs_data_and_ssc & (reg_act_config_is_zero_first_sva_dfm_4_enexo_5
      | reg_act_regs_data_2_15_sva_8_21_0_enexo | reg_w_load_lpi_1_dfm_1_enexo_5
      | reg_is_start_enexo_5 | reg_act_regs_data_3_14_sva_dfm_2_21_0_enexo | reg_act_regs_data_3_14_sva_8_21_0_enexo);
  assign act_regs_data_and_2536_enex5 = act_regs_data_and_ssc & (reg_w_load_lpi_1_dfm_1_enexo_6
      | reg_is_start_enexo_6 | reg_act_regs_data_2_14_sva_8_30_26_enexo | reg_act_config_is_zero_first_sva_dfm_4_enexo_6
      | reg_act_regs_data_3_13_sva_dfm_2_30_26_enexo | reg_act_regs_data_3_13_sva_8_30_26_enexo);
  assign act_regs_data_and_2537_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_3_13_sva_8_25_22_enexo
      | reg_act_regs_data_2_14_sva_8_25_22_enexo | reg_w_load_lpi_1_dfm_1_enexo_7
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_7 | reg_is_start_enexo_7 | reg_act_regs_data_3_13_sva_dfm_2_25_22_enexo);
  assign act_regs_data_and_2538_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_2_14_sva_8_21_0_enexo
      | reg_act_regs_data_3_13_sva_dfm_2_21_0_enexo | reg_act_regs_data_3_13_sva_8_21_0_enexo
      | reg_w_load_lpi_1_dfm_1_enexo_8 | reg_is_start_enexo_8 | reg_act_config_is_zero_first_sva_dfm_4_enexo_8);
  assign act_regs_data_and_2539_enex5 = act_regs_data_and_ssc & (reg_act_config_is_zero_first_sva_dfm_4_enexo_9
      | reg_act_regs_data_2_13_sva_8_30_26_enexo | reg_is_start_enexo_9 | reg_act_regs_data_3_12_sva_8_30_26_enexo
      | reg_act_regs_data_3_12_sva_dfm_2_30_26_enexo | reg_w_load_lpi_1_dfm_1_enexo_9);
  assign act_regs_data_and_2540_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_3_12_sva_dfm_2_25_22_enexo
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_10 | reg_act_regs_data_3_12_sva_8_25_22_enexo
      | reg_is_start_enexo_10 | reg_w_load_lpi_1_dfm_1_enexo_10 | reg_act_regs_data_2_13_sva_8_25_22_enexo);
  assign act_regs_data_and_2541_enex5 = act_regs_data_and_ssc & (reg_w_load_lpi_1_dfm_1_enexo_11
      | reg_act_regs_data_3_12_sva_dfm_2_21_0_enexo | reg_act_regs_data_2_13_sva_8_21_0_enexo
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_11 | reg_act_regs_data_3_12_sva_8_21_0_enexo
      | reg_is_start_enexo_11);
  assign act_regs_data_and_2542_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_3_11_sva_dfm_2_30_26_enexo
      | reg_w_load_lpi_1_dfm_1_enexo_12 | reg_act_regs_data_2_12_sva_8_30_26_enexo
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_12 | reg_is_start_enexo_12 |
      reg_act_regs_data_3_11_sva_8_30_26_enexo);
  assign act_regs_data_and_2543_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_3_11_sva_dfm_2_25_22_enexo
      | reg_w_load_lpi_1_dfm_1_enexo_13 | reg_act_regs_data_2_12_sva_8_25_22_enexo
      | reg_act_regs_data_3_11_sva_8_25_22_enexo | reg_is_start_enexo_13 | reg_act_config_is_zero_first_sva_dfm_4_enexo_13);
  assign act_regs_data_and_2544_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_3_11_sva_dfm_2_21_0_enexo
      | reg_act_regs_data_2_12_sva_8_21_0_enexo | reg_is_start_enexo_14 | reg_w_load_lpi_1_dfm_1_enexo_14
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_14 | reg_act_regs_data_3_11_sva_8_21_0_enexo);
  assign act_regs_data_and_2545_enex5 = act_regs_data_and_ssc & (reg_w_load_lpi_1_dfm_1_enexo_15
      | reg_act_regs_data_2_11_sva_8_30_26_enexo | reg_act_config_is_zero_first_sva_dfm_4_enexo_15
      | reg_act_regs_data_3_10_sva_8_30_26_enexo | reg_is_start_enexo_15 | reg_act_regs_data_3_10_sva_dfm_2_30_26_enexo);
  assign act_regs_data_and_2546_enex5 = act_regs_data_and_ssc & (reg_w_load_lpi_1_dfm_1_enexo_16
      | reg_is_start_enexo_16 | reg_act_config_is_zero_first_sva_dfm_4_enexo_16 |
      reg_act_regs_data_3_10_sva_dfm_2_25_22_enexo | reg_act_regs_data_2_11_sva_8_25_22_enexo
      | reg_act_regs_data_3_10_sva_8_25_22_enexo);
  assign act_regs_data_and_2547_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_2_11_sva_8_21_0_enexo
      | reg_w_load_lpi_1_dfm_1_enexo_17 | reg_act_regs_data_3_10_sva_dfm_2_21_0_enexo
      | reg_is_start_enexo_17 | reg_act_regs_data_3_10_sva_8_21_0_enexo | reg_act_config_is_zero_first_sva_dfm_4_enexo_17);
  assign act_regs_data_and_2548_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_3_9_sva_8_30_26_enexo
      | reg_act_regs_data_3_9_sva_dfm_2_30_26_enexo | reg_act_regs_data_3_0_sva_8_30_26_enexo
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_18 | reg_is_start_enexo_18 |
      reg_w_load_lpi_1_dfm_1_enexo_18);
  assign act_regs_data_and_2549_enex5 = act_regs_data_and_ssc & (reg_w_load_lpi_1_dfm_1_enexo_19
      | reg_act_regs_data_3_9_sva_8_25_22_enexo | reg_act_regs_data_3_9_sva_dfm_2_25_22_enexo
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_19 | reg_is_start_enexo_19 |
      reg_act_regs_data_3_0_sva_8_25_22_enexo);
  assign act_regs_data_and_2550_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_3_9_sva_dfm_2_21_0_enexo
      | reg_act_regs_data_3_9_sva_8_21_0_enexo | reg_is_start_enexo_20 | reg_w_load_lpi_1_dfm_1_enexo_20
      | reg_act_regs_data_3_0_sva_8_21_0_enexo | reg_act_config_is_zero_first_sva_dfm_4_enexo_20);
  assign act_regs_data_and_2551_enex5 = act_regs_data_and_ssc & (reg_is_start_enexo_21
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_21 | reg_act_regs_data_3_8_sva_dfm_2_30_26_enexo
      | reg_act_regs_data_2_9_sva_8_30_26_enexo | reg_w_load_lpi_1_dfm_1_enexo_21
      | reg_act_regs_data_3_8_sva_8_30_26_enexo);
  assign act_regs_data_and_2552_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_2_9_sva_8_25_22_enexo
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_22 | reg_act_regs_data_3_8_sva_8_25_22_enexo
      | reg_is_start_enexo_22 | reg_act_regs_data_3_8_sva_dfm_2_25_22_enexo | reg_w_load_lpi_1_dfm_1_enexo_22);
  assign act_regs_data_and_2553_enex5 = act_regs_data_and_ssc & (reg_w_load_lpi_1_dfm_1_enexo_23
      | reg_act_regs_data_3_8_sva_8_21_0_enexo | reg_is_start_enexo_23 | reg_act_config_is_zero_first_sva_dfm_4_enexo_23
      | reg_act_regs_data_2_9_sva_8_21_0_enexo | reg_act_regs_data_3_8_sva_dfm_2_21_0_enexo);
  assign act_regs_data_and_2554_enex5 = act_regs_data_and_ssc & (reg_w_load_lpi_1_dfm_1_enexo_24
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_24 | reg_act_regs_data_2_8_sva_8_30_26_enexo
      | reg_act_regs_data_3_7_sva_dfm_2_30_26_enexo | reg_is_start_enexo_24 | reg_act_regs_data_3_7_sva_8_30_26_enexo);
  assign act_regs_data_and_2555_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_3_7_sva_8_25_22_enexo
      | reg_w_load_lpi_1_dfm_1_enexo_25 | reg_act_regs_data_3_7_sva_dfm_2_25_22_enexo
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_25 | reg_is_start_enexo_25 |
      reg_act_regs_data_2_8_sva_8_25_22_enexo);
  assign act_regs_data_and_2556_enex5 = act_regs_data_and_ssc & (reg_is_start_enexo_26
      | reg_w_load_lpi_1_dfm_1_enexo_26 | reg_act_config_is_zero_first_sva_dfm_4_enexo_26
      | reg_act_regs_data_3_7_sva_dfm_2_21_0_enexo | reg_act_regs_data_2_8_sva_8_21_0_enexo
      | reg_act_regs_data_3_7_sva_8_21_0_enexo);
  assign act_regs_data_and_2557_enex5 = act_regs_data_and_ssc & (reg_is_start_enexo_27
      | reg_act_regs_data_2_7_sva_8_30_26_enexo | reg_act_config_is_zero_first_sva_dfm_4_enexo_27
      | reg_w_load_lpi_1_dfm_1_enexo_27 | reg_act_regs_data_3_6_sva_dfm_2_30_26_enexo
      | reg_act_regs_data_3_6_sva_8_30_26_enexo);
  assign act_regs_data_and_2558_enex5 = act_regs_data_and_ssc & (reg_act_config_is_zero_first_sva_dfm_4_enexo_28
      | reg_is_start_enexo_28 | reg_act_regs_data_2_7_sva_8_25_22_enexo | reg_act_regs_data_3_6_sva_dfm_2_25_22_enexo
      | reg_act_regs_data_3_6_sva_8_25_22_enexo | reg_w_load_lpi_1_dfm_1_enexo_28);
  assign act_regs_data_and_2559_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_3_6_sva_dfm_2_21_0_enexo
      | reg_w_load_lpi_1_dfm_1_enexo_29 | reg_act_config_is_zero_first_sva_dfm_4_enexo_29
      | reg_act_regs_data_3_6_sva_8_21_0_enexo | reg_act_regs_data_2_7_sva_8_21_0_enexo
      | reg_is_start_enexo_29);
  assign act_regs_data_and_2560_enex5 = act_regs_data_and_ssc & (reg_w_load_lpi_1_dfm_1_enexo_30
      | reg_is_start_enexo_30 | reg_act_regs_data_3_5_sva_8_30_26_enexo | reg_act_config_is_zero_first_sva_dfm_4_enexo_30
      | reg_act_regs_data_2_6_sva_8_30_26_enexo | reg_act_regs_data_3_5_sva_dfm_2_30_26_enexo);
  assign act_regs_data_and_2561_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_3_5_sva_8_25_22_enexo
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_31 | reg_act_regs_data_2_6_sva_8_25_22_enexo
      | reg_is_start_enexo_31 | reg_w_load_lpi_1_dfm_1_enexo_31 | reg_act_regs_data_3_5_sva_dfm_2_25_22_enexo);
  assign act_regs_data_and_2562_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_3_5_sva_dfm_2_21_0_enexo
      | reg_act_regs_data_2_6_sva_8_21_0_enexo | reg_act_config_is_zero_first_sva_dfm_4_enexo_32
      | reg_act_regs_data_3_5_sva_8_21_0_enexo | reg_is_start_enexo_32 | reg_w_load_lpi_1_dfm_1_enexo_32);
  assign act_regs_data_and_2563_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_2_5_sva_8_30_26_enexo
      | reg_act_regs_data_3_4_sva_dfm_2_30_26_enexo | reg_w_load_lpi_1_dfm_1_enexo_33
      | reg_is_start_enexo_33 | reg_act_regs_data_3_4_sva_8_30_26_enexo | reg_act_config_is_zero_first_sva_dfm_4_enexo_33);
  assign act_regs_data_and_2564_enex5 = act_regs_data_and_ssc & (reg_act_config_is_zero_first_sva_dfm_4_enexo_34
      | reg_w_load_lpi_1_dfm_1_enexo_34 | reg_is_start_enexo_34 | reg_act_regs_data_3_4_sva_8_25_22_enexo
      | reg_act_regs_data_2_5_sva_8_25_22_enexo | reg_act_regs_data_3_4_sva_dfm_2_25_22_enexo);
  assign act_regs_data_and_2565_enex5 = act_regs_data_and_ssc & (reg_is_start_enexo_35
      | reg_act_regs_data_2_5_sva_8_21_0_enexo | reg_w_load_lpi_1_dfm_1_enexo_35
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_35 | reg_act_regs_data_3_4_sva_dfm_2_21_0_enexo
      | reg_act_regs_data_3_4_sva_8_21_0_enexo);
  assign act_regs_data_and_2566_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_3_3_sva_dfm_2_30_26_enexo
      | reg_act_regs_data_2_4_sva_8_30_26_enexo | reg_w_load_lpi_1_dfm_1_enexo_36
      | reg_act_regs_data_3_3_sva_8_30_26_enexo | reg_is_start_enexo_36 | reg_act_config_is_zero_first_sva_dfm_4_enexo_36);
  assign act_regs_data_and_2567_enex5 = act_regs_data_and_ssc & (reg_is_start_enexo_37
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_37 | reg_act_regs_data_2_4_sva_8_25_22_enexo
      | reg_act_regs_data_3_3_sva_8_25_22_enexo | reg_act_regs_data_3_3_sva_dfm_2_25_22_enexo
      | reg_w_load_lpi_1_dfm_1_enexo_37);
  assign act_regs_data_and_2568_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_3_3_sva_8_21_0_enexo
      | reg_w_load_lpi_1_dfm_1_enexo_38 | reg_is_start_enexo_38 | reg_act_config_is_zero_first_sva_dfm_4_enexo_38
      | reg_act_regs_data_2_4_sva_8_21_0_enexo | reg_act_regs_data_3_3_sva_dfm_2_21_0_enexo);
  assign act_regs_data_and_2569_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_2_3_sva_8_30_26_enexo
      | reg_act_regs_data_3_2_sva_8_30_26_enexo | reg_act_config_is_zero_first_sva_dfm_4_enexo_39
      | reg_act_regs_data_3_2_sva_dfm_2_30_26_enexo | reg_w_load_lpi_1_dfm_1_enexo_39
      | reg_is_start_enexo_39);
  assign act_regs_data_and_2570_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_2_3_sva_8_25_22_enexo
      | reg_act_regs_data_3_2_sva_8_25_22_enexo | reg_is_start_enexo_40 | reg_w_load_lpi_1_dfm_1_enexo_40
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_40 | reg_act_regs_data_3_2_sva_dfm_2_25_22_enexo);
  assign act_regs_data_and_2571_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_3_2_sva_8_21_0_enexo
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_41 | reg_is_start_enexo_41 |
      reg_act_regs_data_2_3_sva_8_21_0_enexo | reg_w_load_lpi_1_dfm_1_enexo_41 |
      reg_act_regs_data_3_2_sva_dfm_2_21_0_enexo);
  assign act_regs_data_and_2572_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_3_1_sva_dfm_2_30_26_enexo
      | reg_is_start_enexo_42 | reg_act_regs_data_3_1_sva_8_30_26_enexo | reg_act_regs_data_2_10_sva_8_30_26_enexo
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_42 | reg_w_load_lpi_1_dfm_1_enexo_42);
  assign act_regs_data_and_2573_enex5 = act_regs_data_and_ssc & (reg_act_config_is_zero_first_sva_dfm_4_enexo_43
      | reg_w_load_lpi_1_dfm_1_enexo_43 | reg_act_regs_data_2_10_sva_8_25_22_enexo
      | reg_act_regs_data_3_1_sva_dfm_2_25_22_enexo | reg_is_start_enexo_43 | reg_act_regs_data_3_1_sva_8_25_22_enexo);
  assign act_regs_data_and_2574_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_3_1_sva_8_21_0_enexo
      | reg_is_start_enexo_44 | reg_act_config_is_zero_first_sva_dfm_4_enexo_44 |
      reg_act_regs_data_2_10_sva_8_21_0_enexo | reg_act_regs_data_3_1_sva_dfm_2_21_0_enexo
      | reg_w_load_lpi_1_dfm_1_enexo_44);
  assign act_regs_data_and_2575_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_3_0_sva_dfm_2_30_26_enexo
      | reg_act_regs_data_2_1_sva_8_30_26_enexo | reg_w_load_lpi_1_dfm_1_enexo_45
      | reg_act_regs_data_3_0_sva_8_30_26_enexo_1 | reg_act_config_is_zero_first_sva_dfm_4_enexo_45
      | reg_is_start_enexo_45);
  assign act_regs_data_and_2576_enex5 = act_regs_data_and_ssc & (reg_act_config_is_zero_first_sva_dfm_4_enexo_46
      | reg_act_regs_data_3_0_sva_8_25_22_enexo_1 | reg_is_start_enexo_46 | reg_w_load_lpi_1_dfm_1_enexo_46
      | reg_act_regs_data_3_0_sva_dfm_2_25_22_enexo | reg_act_regs_data_2_1_sva_8_25_22_enexo);
  assign act_regs_data_and_2577_enex5 = act_regs_data_and_ssc & (reg_w_load_lpi_1_dfm_1_enexo_47
      | reg_is_start_enexo_47 | reg_act_regs_data_3_0_sva_dfm_2_21_0_enexo | reg_act_regs_data_2_1_sva_8_21_0_enexo
      | reg_act_regs_data_3_0_sva_8_21_0_enexo_1 | reg_act_config_is_zero_first_sva_dfm_4_enexo_47);
  assign act_regs_data_and_2578_enex5 = act_regs_data_and_ssc & (reg_act_config_is_zero_first_sva_dfm_4_enexo_48
      | reg_act_regs_data_2_15_sva_dfm_2_30_26_enexo | reg_act_regs_data_1_2_sva_8_30_26_enexo
      | reg_act_regs_data_2_15_sva_8_30_26_enexo_1 | reg_is_start_enexo_48 | reg_w_load_lpi_1_dfm_1_enexo_48);
  assign act_regs_data_and_2579_enex5 = act_regs_data_and_ssc & (reg_is_start_enexo_49
      | reg_act_regs_data_2_15_sva_dfm_2_25_22_enexo | reg_w_load_lpi_1_dfm_1_enexo_49
      | reg_act_regs_data_1_2_sva_8_25_22_enexo | reg_act_regs_data_2_15_sva_8_25_22_enexo_1
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_49);
  assign act_regs_data_and_2580_enex5 = act_regs_data_and_ssc & (reg_w_load_lpi_1_dfm_1_enexo_50
      | reg_is_start_enexo_50 | reg_act_regs_data_1_2_sva_8_21_0_enexo | reg_act_regs_data_2_15_sva_dfm_2_21_0_enexo
      | reg_act_regs_data_2_15_sva_8_21_0_enexo_1 | reg_act_config_is_zero_first_sva_dfm_4_enexo_50);
  assign act_regs_data_and_2581_enex5 = act_regs_data_and_ssc & (reg_w_load_lpi_1_dfm_1_enexo_51
      | reg_is_start_enexo_51 | reg_act_regs_data_1_15_sva_8_30_26_enexo | reg_act_config_is_zero_first_sva_dfm_4_enexo_51
      | reg_act_regs_data_2_14_sva_dfm_2_30_26_enexo | reg_act_regs_data_2_14_sva_8_30_26_enexo_1);
  assign act_regs_data_and_2582_enex5 = act_regs_data_and_ssc & (reg_act_config_is_zero_first_sva_dfm_4_enexo_52
      | reg_w_load_lpi_1_dfm_1_enexo_52 | reg_act_regs_data_1_15_sva_8_25_22_enexo
      | reg_act_regs_data_2_14_sva_8_25_22_enexo_1 | reg_act_regs_data_2_14_sva_dfm_2_25_22_enexo
      | reg_is_start_enexo_52);
  assign act_regs_data_and_2583_enex5 = act_regs_data_and_ssc & (reg_act_config_is_zero_first_sva_dfm_4_enexo_53
      | reg_act_regs_data_2_14_sva_8_21_0_enexo_1 | reg_act_regs_data_1_15_sva_8_21_0_enexo
      | reg_w_load_lpi_1_dfm_1_enexo_53 | reg_is_start_enexo_53 | reg_act_regs_data_2_14_sva_dfm_2_21_0_enexo);
  assign act_regs_data_and_2584_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_2_13_sva_dfm_2_30_26_enexo
      | reg_act_regs_data_1_14_sva_8_30_26_enexo | reg_act_regs_data_2_13_sva_8_30_26_enexo_1
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_54 | reg_w_load_lpi_1_dfm_1_enexo_54
      | reg_is_start_enexo_54);
  assign act_regs_data_and_2585_enex5 = act_regs_data_and_ssc & (reg_act_config_is_zero_first_sva_dfm_4_enexo_55
      | reg_act_regs_data_2_13_sva_8_25_22_enexo_1 | reg_act_regs_data_1_14_sva_8_25_22_enexo
      | reg_is_start_enexo_55 | reg_act_regs_data_2_13_sva_dfm_2_25_22_enexo | reg_w_load_lpi_1_dfm_1_enexo_55);
  assign act_regs_data_and_2586_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_2_13_sva_dfm_2_21_0_enexo
      | reg_act_regs_data_2_13_sva_8_21_0_enexo_1 | reg_is_start_enexo_56 | reg_act_config_is_zero_first_sva_dfm_4_enexo_56
      | reg_act_regs_data_1_14_sva_8_21_0_enexo | reg_w_load_lpi_1_dfm_1_enexo_56);
  assign act_regs_data_and_2587_enex5 = act_regs_data_and_ssc & (reg_w_load_lpi_1_dfm_1_enexo_57
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_57 | reg_act_regs_data_2_12_sva_8_30_26_enexo_1
      | reg_act_regs_data_1_13_sva_8_30_26_enexo | reg_act_regs_data_2_12_sva_dfm_2_30_26_enexo
      | reg_is_start_enexo_57);
  assign act_regs_data_and_2588_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_1_13_sva_8_25_22_enexo
      | reg_act_regs_data_2_12_sva_dfm_2_25_22_enexo | reg_act_regs_data_2_12_sva_8_25_22_enexo_1
      | reg_is_start_enexo_58 | reg_act_config_is_zero_first_sva_dfm_4_enexo_58 |
      reg_w_load_lpi_1_dfm_1_enexo_58);
  assign act_regs_data_and_2589_enex5 = act_regs_data_and_ssc & (reg_is_start_enexo_59
      | reg_act_regs_data_2_12_sva_8_21_0_enexo_1 | reg_act_regs_data_1_13_sva_8_21_0_enexo
      | reg_act_regs_data_2_12_sva_dfm_2_21_0_enexo | reg_act_config_is_zero_first_sva_dfm_4_enexo_59
      | reg_w_load_lpi_1_dfm_1_enexo_59);
  assign act_regs_data_and_2590_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_2_11_sva_8_30_26_enexo_1
      | reg_w_load_lpi_1_dfm_1_enexo_60 | reg_act_regs_data_1_12_sva_8_30_26_enexo
      | reg_is_start_enexo_60 | reg_act_regs_data_2_11_sva_dfm_2_30_26_enexo | reg_act_config_is_zero_first_sva_dfm_4_enexo_60);
  assign act_regs_data_and_2591_enex5 = act_regs_data_and_ssc & (reg_act_config_is_zero_first_sva_dfm_4_enexo_61
      | reg_act_regs_data_1_12_sva_8_25_22_enexo | reg_w_load_lpi_1_dfm_1_enexo_61
      | reg_act_regs_data_2_11_sva_8_25_22_enexo_1 | reg_is_start_enexo_61 | reg_act_regs_data_2_11_sva_dfm_2_25_22_enexo);
  assign act_regs_data_and_2592_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_2_11_sva_dfm_2_21_0_enexo
      | reg_act_regs_data_2_11_sva_8_21_0_enexo_1 | reg_act_regs_data_1_12_sva_8_21_0_enexo
      | reg_w_load_lpi_1_dfm_1_enexo_62 | reg_act_config_is_zero_first_sva_dfm_4_enexo_62
      | reg_is_start_enexo_62);
  assign act_regs_data_and_2593_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_2_10_sva_8_30_26_enexo_1
      | reg_act_regs_data_2_10_sva_dfm_2_30_26_enexo | reg_act_regs_data_1_11_sva_8_30_26_enexo
      | reg_w_load_lpi_1_dfm_1_enexo_63 | reg_act_config_is_zero_first_sva_dfm_4_enexo_63
      | reg_is_start_enexo_63);
  assign act_regs_data_and_2594_enex5 = act_regs_data_and_ssc & (reg_w_load_lpi_1_dfm_1_enexo_64
      | reg_act_regs_data_2_10_sva_8_25_22_enexo_1 | reg_act_config_is_zero_first_sva_dfm_4_enexo_64
      | reg_act_regs_data_1_11_sva_8_25_22_enexo | reg_is_start_enexo_64 | reg_act_regs_data_2_10_sva_dfm_2_25_22_enexo);
  assign act_regs_data_and_2595_enex5 = act_regs_data_and_ssc & (reg_act_config_is_zero_first_sva_dfm_4_enexo_65
      | reg_act_regs_data_1_11_sva_8_21_0_enexo | reg_is_start_enexo_65 | reg_w_load_lpi_1_dfm_1_enexo_65
      | reg_act_regs_data_2_10_sva_8_21_0_enexo_1 | reg_act_regs_data_2_10_sva_dfm_2_21_0_enexo);
  assign act_regs_data_and_2596_enex5 = act_regs_data_and_ssc & (reg_is_start_enexo_66
      | reg_act_regs_data_2_9_sva_dfm_2_30_26_enexo | reg_act_regs_data_2_9_sva_8_30_26_enexo_1
      | reg_w_load_lpi_1_dfm_1_enexo_66 | reg_act_regs_data_2_0_sva_8_30_26_enexo
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_66);
  assign act_regs_data_and_2597_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_2_0_sva_8_25_22_enexo
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_67 | reg_act_regs_data_2_9_sva_dfm_2_25_22_enexo
      | reg_act_regs_data_2_9_sva_8_25_22_enexo_1 | reg_w_load_lpi_1_dfm_1_enexo_67
      | reg_is_start_enexo_67);
  assign act_regs_data_and_2598_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_2_0_sva_8_21_0_enexo
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_68 | reg_act_regs_data_2_9_sva_8_21_0_enexo_1
      | reg_act_regs_data_2_9_sva_dfm_2_21_0_enexo | reg_is_start_enexo_68 | reg_w_load_lpi_1_dfm_1_enexo_68);
  assign act_regs_data_and_2599_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_2_8_sva_dfm_2_30_26_enexo
      | reg_is_start_enexo_69 | reg_w_load_lpi_1_dfm_1_enexo_69 | reg_act_config_is_zero_first_sva_dfm_4_enexo_69
      | reg_act_regs_data_2_8_sva_8_30_26_enexo_1 | reg_act_regs_data_1_9_sva_8_30_26_enexo);
  assign act_regs_data_and_2600_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_2_8_sva_dfm_2_25_22_enexo
      | reg_w_load_lpi_1_dfm_1_enexo_70 | reg_act_config_is_zero_first_sva_dfm_4_enexo_70
      | reg_act_regs_data_2_8_sva_8_25_22_enexo_1 | reg_is_start_enexo_70 | reg_act_regs_data_1_9_sva_8_25_22_enexo);
  assign act_regs_data_and_2601_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_1_9_sva_8_21_0_enexo
      | reg_act_regs_data_2_8_sva_8_21_0_enexo_1 | reg_act_config_is_zero_first_sva_dfm_4_enexo_71
      | reg_w_load_lpi_1_dfm_1_enexo_71 | reg_is_start_enexo_71 | reg_act_regs_data_2_8_sva_dfm_2_21_0_enexo);
  assign act_regs_data_and_2602_enex5 = act_regs_data_and_ssc & (reg_w_load_lpi_1_dfm_1_enexo_72
      | reg_is_start_enexo_72 | reg_act_regs_data_1_8_sva_8_30_26_enexo | reg_act_regs_data_2_7_sva_dfm_2_30_26_enexo
      | reg_act_regs_data_2_7_sva_8_30_26_enexo_1 | reg_act_config_is_zero_first_sva_dfm_4_enexo_72);
  assign act_regs_data_and_2603_enex5 = act_regs_data_and_ssc & (reg_is_start_enexo_73
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_73 | reg_act_regs_data_2_7_sva_8_25_22_enexo_1
      | reg_act_regs_data_2_7_sva_dfm_2_25_22_enexo | reg_act_regs_data_1_8_sva_8_25_22_enexo
      | reg_w_load_lpi_1_dfm_1_enexo_73);
  assign act_regs_data_and_2604_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_2_7_sva_dfm_2_21_0_enexo
      | reg_is_start_enexo_74 | reg_w_load_lpi_1_dfm_1_enexo_74 | reg_act_config_is_zero_first_sva_dfm_4_enexo_74
      | reg_act_regs_data_2_7_sva_8_21_0_enexo_1 | reg_act_regs_data_1_8_sva_8_21_0_enexo);
  assign act_regs_data_and_2605_enex5 = act_regs_data_and_ssc & (reg_w_load_lpi_1_dfm_1_enexo_75
      | reg_act_regs_data_1_7_sva_8_30_26_enexo | reg_is_start_enexo_75 | reg_act_regs_data_2_6_sva_8_30_26_enexo_1
      | reg_act_regs_data_2_6_sva_dfm_2_30_26_enexo | reg_act_config_is_zero_first_sva_dfm_4_enexo_75);
  assign act_regs_data_and_2606_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_2_6_sva_8_25_22_enexo_1
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_76 | reg_act_regs_data_1_7_sva_8_25_22_enexo
      | reg_act_regs_data_2_6_sva_dfm_2_25_22_enexo | reg_w_load_lpi_1_dfm_1_enexo_76
      | reg_is_start_enexo_76);
  assign act_regs_data_and_2607_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_1_7_sva_8_21_0_enexo
      | reg_w_load_lpi_1_dfm_1_enexo_77 | reg_act_config_is_zero_first_sva_dfm_4_enexo_77
      | reg_act_regs_data_2_6_sva_dfm_2_21_0_enexo | reg_is_start_enexo_77 | reg_act_regs_data_2_6_sva_8_21_0_enexo_1);
  assign act_regs_data_and_2608_enex5 = act_regs_data_and_ssc & (reg_w_load_lpi_1_dfm_1_enexo_78
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_78 | reg_is_start_enexo_78 |
      reg_act_regs_data_1_6_sva_8_30_26_enexo | reg_act_regs_data_2_5_sva_dfm_2_30_26_enexo
      | reg_act_regs_data_2_5_sva_8_30_26_enexo_1);
  assign act_regs_data_and_2609_enex5 = act_regs_data_and_ssc & (reg_w_load_lpi_1_dfm_1_enexo_79
      | reg_is_start_enexo_79 | reg_act_config_is_zero_first_sva_dfm_4_enexo_79 |
      reg_act_regs_data_1_6_sva_8_25_22_enexo | reg_act_regs_data_2_5_sva_8_25_22_enexo_1
      | reg_act_regs_data_2_5_sva_dfm_2_25_22_enexo);
  assign act_regs_data_and_2610_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_1_6_sva_8_21_0_enexo
      | reg_act_regs_data_2_5_sva_8_21_0_enexo_1 | reg_w_load_lpi_1_dfm_1_enexo_80
      | reg_is_start_enexo_80 | reg_act_config_is_zero_first_sva_dfm_4_enexo_80 |
      reg_act_regs_data_2_5_sva_dfm_2_21_0_enexo);
  assign act_regs_data_and_2611_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_1_5_sva_8_30_26_enexo
      | reg_is_start_enexo_81 | reg_w_load_lpi_1_dfm_1_enexo_81 | reg_act_regs_data_2_4_sva_8_30_26_enexo_1
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_81 | reg_act_regs_data_2_4_sva_dfm_2_30_26_enexo);
  assign act_regs_data_and_2612_enex5 = act_regs_data_and_ssc & (reg_act_config_is_zero_first_sva_dfm_4_enexo_82
      | reg_act_regs_data_2_4_sva_8_25_22_enexo_1 | reg_act_regs_data_2_4_sva_dfm_2_25_22_enexo
      | reg_act_regs_data_1_5_sva_8_25_22_enexo | reg_w_load_lpi_1_dfm_1_enexo_82
      | reg_is_start_enexo_82);
  assign act_regs_data_and_2613_enex5 = act_regs_data_and_ssc & (reg_is_start_enexo_83
      | reg_act_regs_data_1_5_sva_8_21_0_enexo | reg_w_load_lpi_1_dfm_1_enexo_83
      | reg_act_regs_data_2_4_sva_dfm_2_21_0_enexo | reg_act_config_is_zero_first_sva_dfm_4_enexo_83
      | reg_act_regs_data_2_4_sva_8_21_0_enexo_1);
  assign act_regs_data_and_2614_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_2_3_sva_8_30_26_enexo_1
      | reg_w_load_lpi_1_dfm_1_enexo_84 | reg_is_start_enexo_84 | reg_act_config_is_zero_first_sva_dfm_4_enexo_84
      | reg_act_regs_data_1_4_sva_8_30_26_enexo | reg_act_regs_data_2_3_sva_dfm_2_30_26_enexo);
  assign act_regs_data_and_2615_enex5 = act_regs_data_and_ssc & (reg_w_load_lpi_1_dfm_1_enexo_85
      | reg_act_regs_data_2_3_sva_dfm_2_25_22_enexo | reg_act_config_is_zero_first_sva_dfm_4_enexo_85
      | reg_is_start_enexo_85 | reg_act_regs_data_1_4_sva_8_25_22_enexo | reg_act_regs_data_2_3_sva_8_25_22_enexo_1);
  assign act_regs_data_and_2616_enex5 = act_regs_data_and_ssc & (reg_is_start_enexo_86
      | reg_act_regs_data_2_3_sva_dfm_2_21_0_enexo | reg_w_load_lpi_1_dfm_1_enexo_86
      | reg_act_regs_data_1_4_sva_8_21_0_enexo | reg_act_config_is_zero_first_sva_dfm_4_enexo_86
      | reg_act_regs_data_2_3_sva_8_21_0_enexo_1);
  assign act_regs_data_and_2617_enex5 = act_regs_data_and_ssc & (reg_act_config_is_zero_first_sva_dfm_4_enexo_87
      | reg_act_regs_data_2_2_sva_8_30_26_enexo_1 | reg_is_start_enexo_87 | reg_w_load_lpi_1_dfm_1_enexo_87
      | reg_act_regs_data_1_3_sva_8_30_26_enexo | reg_act_regs_data_2_2_sva_dfm_2_30_26_enexo);
  assign act_regs_data_and_2618_enex5 = act_regs_data_and_ssc & (reg_is_start_enexo_88
      | reg_w_load_lpi_1_dfm_1_enexo_88 | reg_act_regs_data_2_2_sva_dfm_2_25_22_enexo
      | reg_act_regs_data_2_2_sva_8_25_22_enexo_1 | reg_act_config_is_zero_first_sva_dfm_4_enexo_88
      | reg_act_regs_data_1_3_sva_8_25_22_enexo);
  assign act_regs_data_and_2619_enex5 = act_regs_data_and_ssc & (reg_w_load_lpi_1_dfm_1_enexo_89
      | reg_act_regs_data_2_2_sva_dfm_2_21_0_enexo | reg_act_regs_data_2_2_sva_8_21_0_enexo_1
      | reg_act_regs_data_1_3_sva_8_21_0_enexo | reg_act_config_is_zero_first_sva_dfm_4_enexo_89
      | reg_is_start_enexo_89);
  assign act_regs_data_and_2620_enex5 = act_regs_data_and_ssc & (reg_act_config_is_zero_first_sva_dfm_4_enexo_90
      | reg_act_regs_data_2_1_sva_8_30_26_enexo_1 | reg_is_start_enexo_90 | reg_w_load_lpi_1_dfm_1_enexo_90
      | reg_act_regs_data_1_10_sva_8_30_26_enexo | reg_act_regs_data_2_1_sva_dfm_2_30_26_enexo);
  assign act_regs_data_and_2621_enex5 = act_regs_data_and_ssc & (reg_act_config_is_zero_first_sva_dfm_4_enexo_91
      | reg_act_regs_data_1_10_sva_8_25_22_enexo | reg_is_start_enexo_91 | reg_w_load_lpi_1_dfm_1_enexo_91
      | reg_act_regs_data_2_1_sva_8_25_22_enexo_1 | reg_act_regs_data_2_1_sva_dfm_2_25_22_enexo);
  assign act_regs_data_and_2622_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_2_1_sva_dfm_2_21_0_enexo
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_92 | reg_act_regs_data_1_10_sva_8_21_0_enexo
      | reg_is_start_enexo_92 | reg_act_regs_data_2_1_sva_8_21_0_enexo_1 | reg_w_load_lpi_1_dfm_1_enexo_92);
  assign act_regs_data_and_2623_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_1_1_sva_8_30_26_enexo
      | reg_act_regs_data_2_0_sva_8_30_26_enexo_1 | reg_is_start_enexo_93 | reg_act_config_is_zero_first_sva_dfm_4_enexo_93
      | reg_w_load_lpi_1_dfm_1_enexo_93 | reg_act_regs_data_2_0_sva_dfm_2_30_26_enexo);
  assign act_regs_data_and_2624_enex5 = act_regs_data_and_ssc & (reg_is_start_enexo_94
      | reg_act_regs_data_2_0_sva_dfm_2_25_22_enexo | reg_act_regs_data_2_0_sva_8_25_22_enexo_1
      | reg_w_load_lpi_1_dfm_1_enexo_94 | reg_act_config_is_zero_first_sva_dfm_4_enexo_94
      | reg_act_regs_data_1_1_sva_8_25_22_enexo);
  assign act_regs_data_and_2625_enex5 = act_regs_data_and_ssc & (reg_act_config_is_zero_first_sva_dfm_4_enexo_95
      | reg_act_regs_data_2_0_sva_dfm_2_21_0_enexo | reg_is_start_enexo_95 | reg_w_load_lpi_1_dfm_1_enexo_95
      | reg_act_regs_data_1_1_sva_8_21_0_enexo | reg_act_regs_data_2_0_sva_8_21_0_enexo_1);
  assign act_regs_data_and_2626_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_1_15_sva_dfm_2_30_26_enexo
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_96 | reg_act_regs_data_0_2_sva_8_30_26_enexo
      | reg_w_load_lpi_1_dfm_1_enexo_96 | reg_act_regs_data_1_15_sva_8_30_26_enexo_1
      | reg_is_start_enexo_96);
  assign act_regs_data_and_2627_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_1_15_sva_dfm_2_25_22_enexo
      | reg_act_regs_data_0_2_sva_8_25_22_enexo | reg_w_load_lpi_1_dfm_1_enexo_97
      | reg_act_regs_data_1_15_sva_8_25_22_enexo_1 | reg_is_start_enexo_97 | reg_act_config_is_zero_first_sva_dfm_4_enexo_97);
  assign act_regs_data_and_2628_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_1_15_sva_dfm_2_21_0_enexo
      | reg_w_load_lpi_1_dfm_1_enexo_98 | reg_is_start_enexo_98 | reg_act_regs_data_1_15_sva_8_21_0_enexo_1
      | reg_act_regs_data_0_2_sva_8_21_0_enexo | reg_act_config_is_zero_first_sva_dfm_4_enexo_98);
  assign act_regs_data_and_2629_enex5 = act_regs_data_and_ssc & (reg_is_start_enexo_99
      | reg_act_regs_data_0_15_sva_8_30_26_enexo | reg_act_regs_data_1_14_sva_8_30_26_enexo_1
      | reg_act_regs_data_1_14_sva_dfm_2_30_26_enexo | reg_w_load_lpi_1_dfm_1_enexo_99
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_99);
  assign act_regs_data_and_2630_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_1_14_sva_dfm_2_25_22_enexo
      | reg_act_regs_data_0_15_sva_8_25_22_enexo | reg_is_start_enexo_100 | reg_w_load_lpi_1_dfm_1_enexo_100
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_100 | reg_act_regs_data_1_14_sva_8_25_22_enexo_1);
  assign act_regs_data_and_2631_enex5 = act_regs_data_and_ssc & (reg_act_config_is_zero_first_sva_dfm_4_enexo_101
      | reg_w_load_lpi_1_dfm_1_enexo_101 | reg_is_start_enexo_101 | reg_act_regs_data_0_15_sva_8_21_0_enexo
      | reg_act_regs_data_1_14_sva_dfm_2_21_0_enexo | reg_act_regs_data_1_14_sva_8_21_0_enexo_1);
  assign act_regs_data_and_2632_enex5 = act_regs_data_and_ssc & (reg_w_load_lpi_1_dfm_1_enexo_102
      | reg_act_regs_data_1_13_sva_8_30_26_enexo_1 | reg_act_regs_data_1_13_sva_dfm_2_30_26_enexo
      | reg_is_start_enexo_102 | reg_act_regs_data_0_14_sva_8_30_26_enexo | reg_act_config_is_zero_first_sva_dfm_4_enexo_102);
  assign act_regs_data_and_2633_enex5 = act_regs_data_and_ssc & (reg_act_config_is_zero_first_sva_dfm_4_enexo_103
      | reg_is_start_enexo_103 | reg_w_load_lpi_1_dfm_1_enexo_103 | reg_act_regs_data_1_13_sva_dfm_2_25_22_enexo
      | reg_act_regs_data_0_14_sva_8_25_22_enexo | reg_act_regs_data_1_13_sva_8_25_22_enexo_1);
  assign act_regs_data_and_2634_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_1_13_sva_dfm_2_21_0_enexo
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_104 | reg_is_start_enexo_104
      | reg_act_regs_data_0_14_sva_8_21_0_enexo | reg_act_regs_data_1_13_sva_8_21_0_enexo_1
      | reg_w_load_lpi_1_dfm_1_enexo_104);
  assign act_regs_data_and_2635_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_1_12_sva_8_30_26_enexo_1
      | reg_w_load_lpi_1_dfm_1_enexo_105 | reg_act_config_is_zero_first_sva_dfm_4_enexo_105
      | reg_act_regs_data_0_13_sva_8_30_26_enexo | reg_is_start_enexo_105 | reg_act_regs_data_1_12_sva_dfm_2_30_26_enexo);
  assign act_regs_data_and_2636_enex5 = act_regs_data_and_ssc & (reg_is_start_enexo_106
      | reg_act_regs_data_1_12_sva_dfm_2_25_22_enexo | reg_act_regs_data_0_13_sva_8_25_22_enexo
      | reg_w_load_lpi_1_dfm_1_enexo_106 | reg_act_config_is_zero_first_sva_dfm_4_enexo_106
      | reg_act_regs_data_1_12_sva_8_25_22_enexo_1);
  assign act_regs_data_and_2637_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_1_12_sva_dfm_2_21_0_enexo
      | reg_act_regs_data_1_12_sva_8_21_0_enexo_1 | reg_is_start_enexo_107 | reg_w_load_lpi_1_dfm_1_enexo_107
      | reg_act_regs_data_0_13_sva_8_21_0_enexo | reg_act_config_is_zero_first_sva_dfm_4_enexo_107);
  assign act_regs_data_and_2638_enex5 = act_regs_data_and_ssc & (reg_w_load_lpi_1_dfm_1_enexo_108
      | reg_is_start_enexo_108 | reg_act_regs_data_1_11_sva_dfm_2_30_26_enexo | reg_act_config_is_zero_first_sva_dfm_4_enexo_108
      | reg_act_regs_data_1_11_sva_8_30_26_enexo_1 | reg_act_regs_data_0_12_sva_8_30_26_enexo);
  assign act_regs_data_and_2639_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_1_11_sva_dfm_2_25_22_enexo
      | reg_is_start_enexo_109 | reg_act_regs_data_1_11_sva_8_25_22_enexo_1 | reg_w_load_lpi_1_dfm_1_enexo_109
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_109 | reg_act_regs_data_0_12_sva_8_25_22_enexo);
  assign act_regs_data_and_2640_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_1_11_sva_8_21_0_enexo_1
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_110 | reg_is_start_enexo_110
      | reg_w_load_lpi_1_dfm_1_enexo_110 | reg_act_regs_data_1_11_sva_dfm_2_21_0_enexo
      | reg_act_regs_data_0_12_sva_8_21_0_enexo);
  assign act_regs_data_and_2641_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_1_10_sva_dfm_2_30_26_enexo
      | reg_act_regs_data_0_11_sva_8_30_26_enexo | reg_act_regs_data_1_10_sva_8_30_26_enexo_1
      | reg_w_load_lpi_1_dfm_1_enexo_111 | reg_act_config_is_zero_first_sva_dfm_4_enexo_111
      | reg_is_start_enexo_111);
  assign act_regs_data_and_2642_enex5 = act_regs_data_and_ssc & (reg_is_start_enexo_112
      | reg_act_regs_data_1_10_sva_8_25_22_enexo_1 | reg_w_load_lpi_1_dfm_1_enexo_112
      | reg_act_regs_data_1_10_sva_dfm_2_25_22_enexo | reg_act_config_is_zero_first_sva_dfm_4_enexo_112
      | reg_act_regs_data_0_11_sva_8_25_22_enexo);
  assign act_regs_data_and_2643_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_1_10_sva_dfm_2_21_0_enexo
      | reg_act_regs_data_1_10_sva_8_21_0_enexo_1 | reg_act_regs_data_0_11_sva_8_21_0_enexo
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_113 | reg_is_start_enexo_113
      | reg_w_load_lpi_1_dfm_1_enexo_113);
  assign act_regs_data_and_2644_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_1_9_sva_8_30_26_enexo_1
      | reg_act_regs_data_1_0_sva_8_30_26_enexo | reg_act_config_is_zero_first_sva_dfm_4_enexo_114
      | reg_act_regs_data_1_9_sva_dfm_2_30_26_enexo | reg_w_load_lpi_1_dfm_1_enexo_114
      | reg_is_start_enexo_114);
  assign act_regs_data_and_2645_enex5 = act_regs_data_and_ssc & (reg_is_start_enexo_115
      | reg_w_load_lpi_1_dfm_1_enexo_115 | reg_act_config_is_zero_first_sva_dfm_4_enexo_115
      | reg_act_regs_data_1_9_sva_dfm_2_25_22_enexo | reg_act_regs_data_1_0_sva_8_25_22_enexo
      | reg_act_regs_data_1_9_sva_8_25_22_enexo_1);
  assign act_regs_data_and_2646_enex5 = act_regs_data_and_ssc & (reg_w_load_lpi_1_dfm_1_enexo_116
      | reg_act_regs_data_1_0_sva_8_21_0_enexo | reg_act_regs_data_1_9_sva_8_21_0_enexo_1
      | reg_is_start_enexo_116 | reg_act_config_is_zero_first_sva_dfm_4_enexo_116
      | reg_act_regs_data_1_9_sva_dfm_2_21_0_enexo);
  assign act_regs_data_and_2647_enex5 = act_regs_data_and_ssc & (reg_is_start_enexo_117
      | reg_act_regs_data_1_8_sva_8_30_26_enexo_1 | reg_act_config_is_zero_first_sva_dfm_4_enexo_117
      | reg_act_regs_data_0_9_sva_8_30_26_enexo | reg_w_load_lpi_1_dfm_1_enexo_117
      | reg_act_regs_data_1_8_sva_dfm_2_30_26_enexo);
  assign act_regs_data_and_2648_enex5 = act_regs_data_and_ssc & (reg_act_config_is_zero_first_sva_dfm_4_enexo_118
      | reg_act_regs_data_1_8_sva_dfm_2_25_22_enexo | reg_act_regs_data_1_8_sva_8_25_22_enexo_1
      | reg_act_regs_data_0_9_sva_8_25_22_enexo | reg_is_start_enexo_118 | reg_w_load_lpi_1_dfm_1_enexo_118);
  assign act_regs_data_and_2649_enex5 = act_regs_data_and_ssc & (reg_w_load_lpi_1_dfm_1_enexo_119
      | reg_act_regs_data_1_8_sva_8_21_0_enexo_1 | reg_act_regs_data_1_8_sva_dfm_2_21_0_enexo
      | reg_act_regs_data_0_9_sva_8_21_0_enexo | reg_is_start_enexo_119 | reg_act_config_is_zero_first_sva_dfm_4_enexo_119);
  assign act_regs_data_and_2650_enex5 = act_regs_data_and_ssc & (reg_w_load_lpi_1_dfm_1_enexo_120
      | reg_act_regs_data_1_7_sva_dfm_2_30_26_enexo | reg_is_start_enexo_120 | reg_act_config_is_zero_first_sva_dfm_4_enexo_120
      | reg_act_regs_data_0_8_sva_8_30_26_enexo | reg_act_regs_data_1_7_sva_8_30_26_enexo_1);
  assign act_regs_data_and_2651_enex5 = act_regs_data_and_ssc & (reg_w_load_lpi_1_dfm_1_enexo_121
      | reg_act_regs_data_0_8_sva_8_25_22_enexo | reg_act_regs_data_1_7_sva_8_25_22_enexo_1
      | reg_act_regs_data_1_7_sva_dfm_2_25_22_enexo | reg_act_config_is_zero_first_sva_dfm_4_enexo_121
      | reg_is_start_enexo_121);
  assign act_regs_data_and_2652_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_1_7_sva_8_21_0_enexo_1
      | reg_act_regs_data_0_8_sva_8_21_0_enexo | reg_act_regs_data_1_7_sva_dfm_2_21_0_enexo
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_122 | reg_is_start_enexo_122
      | reg_w_load_lpi_1_dfm_1_enexo_122);
  assign act_regs_data_and_2653_enex5 = act_regs_data_and_ssc & (reg_is_start_enexo_123
      | reg_act_regs_data_1_6_sva_dfm_2_30_26_enexo | reg_w_load_lpi_1_dfm_1_enexo_123
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_123 | reg_act_regs_data_0_7_sva_8_30_26_enexo
      | reg_act_regs_data_1_6_sva_8_30_26_enexo_1);
  assign act_regs_data_and_2654_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_0_7_sva_8_25_22_enexo
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_124 | reg_is_start_enexo_124
      | reg_act_regs_data_1_6_sva_dfm_2_25_22_enexo | reg_act_regs_data_1_6_sva_8_25_22_enexo_1
      | reg_w_load_lpi_1_dfm_1_enexo_124);
  assign act_regs_data_and_2655_enex5 = act_regs_data_and_ssc & (reg_act_config_is_zero_first_sva_dfm_4_enexo_125
      | reg_act_regs_data_0_7_sva_8_21_0_enexo | reg_act_regs_data_1_6_sva_dfm_2_21_0_enexo
      | reg_act_regs_data_1_6_sva_8_21_0_enexo_1 | reg_w_load_lpi_1_dfm_1_enexo_125
      | reg_is_start_enexo_125);
  assign act_regs_data_and_2656_enex5 = act_regs_data_and_ssc & (reg_is_start_enexo_126
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_126 | reg_w_load_lpi_1_dfm_1_enexo_126
      | reg_act_regs_data_1_5_sva_8_30_26_enexo_1 | reg_act_regs_data_0_6_sva_8_30_26_enexo
      | reg_act_regs_data_1_5_sva_dfm_2_30_26_enexo);
  assign act_regs_data_and_2657_enex5 = act_regs_data_and_ssc & (reg_act_config_is_zero_first_sva_dfm_4_enexo_127
      | reg_act_regs_data_1_5_sva_dfm_2_25_22_enexo | reg_act_regs_data_1_5_sva_8_25_22_enexo_1
      | reg_w_load_lpi_1_dfm_1_enexo_127 | reg_act_regs_data_0_6_sva_8_25_22_enexo
      | reg_is_start_enexo_127);
  assign act_regs_data_and_2658_enex5 = act_regs_data_and_ssc & (reg_act_config_is_zero_first_sva_dfm_4_enexo_128
      | reg_w_load_lpi_1_dfm_1_enexo_128 | reg_act_regs_data_1_5_sva_8_21_0_enexo_1
      | reg_is_start_enexo_128 | reg_act_regs_data_0_6_sva_8_21_0_enexo | reg_act_regs_data_1_5_sva_dfm_2_21_0_enexo);
  assign act_regs_data_and_2659_enex5 = act_regs_data_and_ssc & (reg_act_config_is_zero_first_sva_dfm_4_enexo_129
      | reg_act_regs_data_1_4_sva_8_30_26_enexo_1 | reg_act_regs_data_0_5_sva_8_30_26_enexo
      | reg_is_start_enexo_129 | reg_act_regs_data_1_4_sva_dfm_2_30_26_enexo | reg_w_load_lpi_1_dfm_1_enexo_129);
  assign act_regs_data_and_2660_enex5 = act_regs_data_and_ssc & (reg_is_start_enexo_130
      | reg_act_regs_data_1_4_sva_dfm_2_25_22_enexo | reg_act_regs_data_0_5_sva_8_25_22_enexo
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_130 | reg_act_regs_data_1_4_sva_8_25_22_enexo_1
      | reg_w_load_lpi_1_dfm_1_enexo_130);
  assign act_regs_data_and_2661_enex5 = act_regs_data_and_ssc & (reg_act_config_is_zero_first_sva_dfm_4_enexo_131
      | reg_act_regs_data_1_4_sva_dfm_2_21_0_enexo | reg_act_regs_data_1_4_sva_8_21_0_enexo_1
      | reg_w_load_lpi_1_dfm_1_enexo_131 | reg_is_start_enexo_131 | reg_act_regs_data_0_5_sva_8_21_0_enexo);
  assign act_regs_data_and_2662_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_1_3_sva_dfm_2_30_26_enexo
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_132 | reg_act_regs_data_1_3_sva_8_30_26_enexo_1
      | reg_is_start_enexo_132 | reg_act_regs_data_0_4_sva_8_30_26_enexo | reg_w_load_lpi_1_dfm_1_enexo_132);
  assign act_regs_data_and_2663_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_1_3_sva_dfm_2_25_22_enexo
      | reg_act_regs_data_0_4_sva_8_25_22_enexo | reg_act_regs_data_1_3_sva_8_25_22_enexo_1
      | reg_w_load_lpi_1_dfm_1_enexo_133 | reg_act_config_is_zero_first_sva_dfm_4_enexo_133
      | reg_is_start_enexo_133);
  assign act_regs_data_and_2664_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_1_3_sva_dfm_2_21_0_enexo
      | reg_act_regs_data_0_4_sva_8_21_0_enexo | reg_act_regs_data_1_3_sva_8_21_0_enexo_1
      | reg_w_load_lpi_1_dfm_1_enexo_134 | reg_is_start_enexo_134 | reg_act_config_is_zero_first_sva_dfm_4_enexo_134);
  assign act_regs_data_and_2665_enex5 = act_regs_data_and_ssc & (reg_w_load_lpi_1_dfm_1_enexo_135
      | reg_is_start_enexo_135 | reg_act_config_is_zero_first_sva_dfm_4_enexo_135
      | reg_act_regs_data_1_2_sva_dfm_2_30_26_enexo | reg_act_regs_data_1_2_sva_8_30_26_enexo_1
      | reg_act_regs_data_0_3_sva_8_30_26_enexo);
  assign act_regs_data_and_2666_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_1_2_sva_dfm_2_25_22_enexo
      | reg_act_regs_data_1_2_sva_8_25_22_enexo_1 | reg_is_start_enexo_136 | reg_act_config_is_zero_first_sva_dfm_4_enexo_136
      | reg_act_regs_data_0_3_sva_8_25_22_enexo | reg_w_load_lpi_1_dfm_1_enexo_136);
  assign act_regs_data_and_2667_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_1_2_sva_8_21_0_enexo_1
      | reg_w_load_lpi_1_dfm_1_enexo_137 | reg_act_regs_data_0_3_sva_8_21_0_enexo
      | reg_act_regs_data_1_2_sva_dfm_2_21_0_enexo | reg_is_start_enexo_137 | reg_act_config_is_zero_first_sva_dfm_4_enexo_137);
  assign act_regs_data_and_2668_enex5 = act_regs_data_and_ssc & (reg_w_load_lpi_1_dfm_1_enexo_138
      | reg_act_regs_data_1_1_sva_dfm_2_30_26_enexo | reg_act_regs_data_0_10_sva_8_30_26_enexo
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_138 | reg_act_regs_data_1_1_sva_8_30_26_enexo_1
      | reg_is_start_enexo_138);
  assign act_regs_data_and_2669_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_1_1_sva_8_25_22_enexo_1
      | reg_act_regs_data_1_1_sva_dfm_2_25_22_enexo | reg_act_config_is_zero_first_sva_dfm_4_enexo_139
      | reg_w_load_lpi_1_dfm_1_enexo_139 | reg_is_start_enexo_139 | reg_act_regs_data_0_10_sva_8_25_22_enexo);
  assign act_regs_data_and_2670_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_1_1_sva_8_21_0_enexo_1
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_140 | reg_is_start_enexo_140
      | reg_act_regs_data_1_1_sva_dfm_2_21_0_enexo | reg_w_load_lpi_1_dfm_1_enexo_140
      | reg_act_regs_data_0_10_sva_8_21_0_enexo);
  assign act_regs_data_and_2671_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_1_0_sva_8_30_26_enexo_1
      | reg_act_regs_data_1_0_sva_dfm_2_30_26_enexo | reg_is_start_enexo_141 | reg_act_regs_data_0_1_sva_8_30_26_enexo
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_141 | reg_w_load_lpi_1_dfm_1_enexo_141);
  assign act_regs_data_and_2672_enex5 = act_regs_data_and_ssc & (reg_act_config_is_zero_first_sva_dfm_4_enexo_142
      | reg_w_load_lpi_1_dfm_1_enexo_142 | reg_act_regs_data_0_1_sva_8_25_22_enexo
      | reg_is_start_enexo_142 | reg_act_regs_data_1_0_sva_dfm_2_25_22_enexo | reg_act_regs_data_1_0_sva_8_25_22_enexo_1);
  assign act_regs_data_and_2673_enex5 = act_regs_data_and_ssc & (reg_is_start_enexo_143
      | reg_w_load_lpi_1_dfm_1_enexo_143 | reg_act_regs_data_1_0_sva_8_21_0_enexo_1
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_143 | reg_act_regs_data_0_1_sva_8_21_0_enexo
      | reg_act_regs_data_1_0_sva_dfm_2_21_0_enexo);
  assign act_regs_data_and_2674_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_0_15_sva_dfm_2_30_26_enexo
      | reg_act_regs_data_0_15_sva_8_30_26_enexo_1 | reg_ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_1_30_26_enexo
      | reg_is_start_enexo_144 | reg_w_load_lpi_1_dfm_1_enexo_144 | reg_act_config_is_zero_first_sva_dfm_4_enexo_144);
  assign act_regs_data_and_2675_enex5 = act_regs_data_and_ssc & (reg_is_start_enexo_145
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_145 | reg_w_load_lpi_1_dfm_1_enexo_145
      | reg_act_regs_data_0_15_sva_8_25_22_enexo_1 | reg_ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_1_25_22_enexo
      | reg_act_regs_data_0_15_sva_dfm_2_25_22_enexo);
  assign act_regs_data_and_2676_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_0_15_sva_8_21_0_enexo_1
      | reg_is_start_enexo_146 | reg_act_config_is_zero_first_sva_dfm_4_enexo_146
      | reg_w_load_lpi_1_dfm_1_enexo_146 | reg_act_regs_data_0_15_sva_dfm_2_21_0_enexo
      | reg_Silu_for_3_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo);
  assign act_regs_data_and_2677_enex5 = act_regs_data_and_ssc & (reg_act_config_is_zero_first_sva_dfm_4_enexo_147
      | reg_is_start_enexo_147 | reg_w_load_lpi_1_dfm_1_enexo_147 | reg_act_regs_data_0_14_sva_8_30_26_enexo_1
      | reg_ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_1_30_26_enexo
      | reg_act_regs_data_0_14_sva_dfm_2_30_26_enexo);
  assign act_regs_data_and_2678_enex5 = act_regs_data_and_ssc & (reg_w_load_lpi_1_dfm_1_enexo_148
      | reg_act_regs_data_0_14_sva_8_25_22_enexo_1 | reg_is_start_enexo_148 | reg_act_config_is_zero_first_sva_dfm_4_enexo_148
      | reg_ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_1_25_22_enexo
      | reg_act_regs_data_0_14_sva_dfm_2_25_22_enexo);
  assign act_regs_data_and_2679_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_0_14_sva_dfm_2_21_0_enexo
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_149 | reg_is_start_enexo_149
      | reg_w_load_lpi_1_dfm_1_enexo_149 | reg_Silu_for_2_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo
      | reg_act_regs_data_0_14_sva_8_21_0_enexo_1);
  assign act_regs_data_and_2680_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_0_0_sva_8_30_26_enexo
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_150 | reg_is_start_enexo_150
      | reg_act_regs_data_0_9_sva_8_30_26_enexo_1 | reg_w_load_lpi_1_dfm_1_enexo_150
      | reg_act_regs_data_0_9_sva_dfm_2_30_26_enexo);
  assign act_regs_data_and_2681_enex5 = act_regs_data_and_ssc & (reg_w_load_lpi_1_dfm_1_enexo_151
      | reg_is_start_enexo_151 | reg_act_config_is_zero_first_sva_dfm_4_enexo_151
      | reg_act_regs_data_0_9_sva_8_25_22_enexo_1 | reg_act_regs_data_0_0_sva_8_25_22_enexo
      | reg_act_regs_data_0_9_sva_dfm_2_25_22_enexo);
  assign act_regs_data_and_2682_enex5 = act_regs_data_and_ssc & (reg_act_config_is_zero_first_sva_dfm_4_enexo_152
      | reg_is_start_enexo_152 | reg_act_regs_data_0_9_sva_8_21_0_enexo_1 | reg_act_regs_data_0_9_sva_dfm_2_21_0_enexo
      | reg_act_regs_data_0_0_sva_8_21_0_enexo | reg_w_load_lpi_1_dfm_1_enexo_152);
  assign act_regs_data_and_2683_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_0_8_sva_dfm_2_30_26_enexo
      | reg_w_load_lpi_1_dfm_1_enexo_153 | reg_is_start_enexo_153 | reg_act_config_is_zero_first_sva_dfm_4_enexo_153
      | reg_ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_1_30_26_enexo |
      reg_act_regs_data_0_8_sva_8_30_26_enexo_1);
  assign act_regs_data_and_2684_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_0_8_sva_8_25_22_enexo_1
      | reg_act_regs_data_0_8_sva_dfm_2_25_22_enexo | reg_w_load_lpi_1_dfm_1_enexo_154
      | reg_ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_1_25_22_enexo |
      reg_act_config_is_zero_first_sva_dfm_4_enexo_154 | reg_is_start_enexo_154);
  assign act_regs_data_and_2685_enex5 = act_regs_data_and_ssc & (reg_Silu_for_y_8_sva_3_24_0_1_enexo
      | reg_act_regs_data_0_8_sva_dfm_2_21_0_enexo | reg_act_regs_data_0_8_sva_8_21_0_enexo_1
      | reg_w_load_lpi_1_dfm_1_enexo_155 | reg_is_start_enexo_155 | reg_act_config_is_zero_first_sva_dfm_4_enexo_155);
  assign act_regs_data_and_2686_enex5 = act_regs_data_and_ssc & (reg_act_config_is_zero_first_sva_dfm_4_enexo_156
      | reg_act_regs_data_0_7_sva_8_30_26_enexo_1 | reg_act_regs_data_0_7_sva_dfm_2_30_26_enexo
      | reg_is_start_enexo_156 | reg_w_load_lpi_1_dfm_1_enexo_156 | reg_ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_1_30_26_enexo);
  assign act_regs_data_and_2687_enex5 = act_regs_data_and_ssc & (reg_is_start_enexo_157
      | reg_w_load_lpi_1_dfm_1_enexo_157 | reg_act_regs_data_0_7_sva_8_25_22_enexo_1
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_157 | reg_act_regs_data_0_7_sva_dfm_2_25_22_enexo
      | reg_ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_1_25_22_enexo);
  assign act_regs_data_and_2688_enex5 = act_regs_data_and_ssc & (reg_w_load_lpi_1_dfm_1_enexo_158
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_158 | reg_Silu_for_y_1_sva_3_24_0_1_enexo
      | reg_act_regs_data_0_7_sva_8_21_0_enexo_1 | reg_is_start_enexo_158 | reg_act_regs_data_0_7_sva_dfm_2_21_0_enexo);
  assign act_regs_data_and_2689_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_0_6_sva_8_30_26_enexo_1
      | reg_is_start_enexo_159 | reg_ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_1_30_26_enexo
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_159 | reg_w_load_lpi_1_dfm_1_enexo_159
      | reg_act_regs_data_0_6_sva_dfm_2_30_26_enexo);
  assign act_regs_data_and_2690_enex5 = act_regs_data_and_ssc & (reg_act_config_is_zero_first_sva_dfm_4_enexo_160
      | reg_w_load_lpi_1_dfm_1_enexo_160 | reg_act_regs_data_0_6_sva_dfm_2_25_22_enexo
      | reg_is_start_enexo_160 | reg_ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_1_25_22_enexo
      | reg_act_regs_data_0_6_sva_8_25_22_enexo_1);
  assign act_regs_data_and_2691_enex5 = act_regs_data_and_ssc & (reg_w_load_lpi_1_dfm_1_enexo_161
      | reg_Silu_for_9_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo
      | reg_act_regs_data_0_6_sva_8_21_0_enexo_1 | reg_is_start_enexo_161 | reg_act_config_is_zero_first_sva_dfm_4_enexo_161
      | reg_act_regs_data_0_6_sva_dfm_2_21_0_enexo);
  assign act_regs_data_and_2692_enex5 = act_regs_data_and_ssc & (reg_w_load_lpi_1_dfm_1_enexo_162
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_162 | reg_act_regs_data_0_5_sva_8_30_26_enexo_1
      | reg_act_regs_data_0_5_sva_dfm_2_30_26_enexo | reg_ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_1_30_26_enexo
      | reg_is_start_enexo_162);
  assign act_regs_data_and_2693_enex5 = act_regs_data_and_ssc & (reg_act_config_is_zero_first_sva_dfm_4_enexo_163
      | reg_act_regs_data_0_5_sva_8_25_22_enexo_1 | reg_is_start_enexo_163 | reg_w_load_lpi_1_dfm_1_enexo_163
      | reg_act_regs_data_0_5_sva_dfm_2_25_22_enexo | reg_ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_1_25_22_enexo);
  assign act_regs_data_and_2694_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_0_5_sva_dfm_2_21_0_enexo
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_164 | reg_act_regs_data_0_5_sva_8_21_0_enexo_1
      | reg_w_load_lpi_1_dfm_1_enexo_164 | reg_Silu_for_7_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo
      | reg_is_start_enexo_164);
  assign act_regs_data_and_2695_enex5 = act_regs_data_and_ssc & (reg_act_config_is_zero_first_sva_dfm_4_enexo_165
      | reg_act_regs_data_0_4_sva_8_30_26_enexo_1 | reg_ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_1_30_26_enexo
      | reg_w_load_lpi_1_dfm_1_enexo_165 | reg_act_regs_data_0_4_sva_dfm_2_30_26_enexo
      | reg_is_start_enexo_165);
  assign act_regs_data_and_2696_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_0_4_sva_8_25_22_enexo_1
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_166 | reg_ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_1_25_22_enexo
      | reg_w_load_lpi_1_dfm_1_enexo_166 | reg_act_regs_data_0_4_sva_dfm_2_25_22_enexo
      | reg_is_start_enexo_166);
  assign act_regs_data_and_2697_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_0_4_sva_8_21_0_enexo_1
      | reg_w_load_lpi_1_dfm_1_enexo_167 | reg_act_config_is_zero_first_sva_dfm_4_enexo_167
      | reg_act_regs_data_0_4_sva_dfm_2_21_0_enexo | reg_Silu_for_6_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo
      | reg_is_start_enexo_167);
  assign act_regs_data_and_2698_enex5 = act_regs_data_and_ssc & (reg_act_config_is_zero_first_sva_dfm_4_enexo_168
      | reg_w_load_lpi_1_dfm_1_enexo_168 | reg_act_regs_data_0_3_sva_dfm_2_30_26_enexo
      | reg_act_regs_data_0_3_sva_8_30_26_enexo_1 | reg_is_start_enexo_168 | reg_ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_1_30_26_enexo);
  assign act_regs_data_and_2699_enex5 = act_regs_data_and_ssc & (reg_is_start_enexo_169
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_169 | reg_act_regs_data_0_3_sva_dfm_2_25_22_enexo
      | reg_w_load_lpi_1_dfm_1_enexo_169 | reg_act_regs_data_0_3_sva_8_25_22_enexo_1
      | reg_ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_1_25_22_enexo);
  assign act_regs_data_and_2700_enex5 = act_regs_data_and_ssc & (reg_w_load_lpi_1_dfm_1_enexo_170
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_170 | reg_act_regs_data_0_3_sva_8_21_0_enexo_1
      | reg_is_start_enexo_170 | reg_act_regs_data_0_3_sva_dfm_2_21_0_enexo | reg_Silu_for_5_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo);
  assign act_regs_data_and_2701_enex5 = act_regs_data_and_ssc & (reg_is_start_enexo_171
      | reg_ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_1_30_26_enexo |
      reg_act_regs_data_0_2_sva_dfm_2_30_26_enexo | reg_act_regs_data_0_2_sva_8_30_26_enexo_1
      | reg_w_load_lpi_1_dfm_1_enexo_171 | reg_act_config_is_zero_first_sva_dfm_4_enexo_171);
  assign act_regs_data_and_2702_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_0_2_sva_dfm_2_25_22_enexo
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_172 | reg_act_regs_data_0_2_sva_8_25_22_enexo_1
      | reg_w_load_lpi_1_dfm_1_enexo_172 | reg_is_start_enexo_172 | reg_ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_1_25_22_enexo);
  assign act_regs_data_and_2703_enex5 = act_regs_data_and_ssc & (reg_is_start_enexo_173
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_173 | reg_act_regs_data_0_2_sva_8_21_0_enexo_1
      | reg_w_load_lpi_1_dfm_1_enexo_173 | reg_Silu_for_4_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo
      | reg_act_regs_data_0_2_sva_dfm_2_21_0_enexo);
  assign act_mem_banks_read_read_data_and_cse = ActUnitRun_wen & and_dcpl_1109 &
      and_dcpl_1106 & (~ act_write_req_valid_lpi_1_dfm_5);
  assign act_mem_banks_read_read_data_and_16_enex5 = act_mem_banks_read_read_data_and_cse
      & reg_act_mem_banks_read_for_mux_15_enexo;
  assign act_mem_banks_read_read_data_and_17_enex5 = act_mem_banks_read_read_data_and_cse
      & reg_act_mem_banks_read_for_mux_14_enexo;
  assign act_mem_banks_read_read_data_and_18_enex5 = act_mem_banks_read_read_data_and_cse
      & reg_act_mem_banks_read_for_mux_13_enexo;
  assign act_mem_banks_read_read_data_and_19_enex5 = act_mem_banks_read_read_data_and_cse
      & reg_act_mem_banks_read_for_mux_12_enexo;
  assign act_mem_banks_read_read_data_and_20_enex5 = act_mem_banks_read_read_data_and_cse
      & reg_act_mem_banks_read_for_mux_11_enexo;
  assign act_mem_banks_read_read_data_and_21_enex5 = act_mem_banks_read_read_data_and_cse
      & reg_act_mem_banks_read_for_mux_10_enexo;
  assign act_mem_banks_read_read_data_and_22_enex5 = act_mem_banks_read_read_data_and_cse
      & reg_act_mem_banks_read_for_mux_9_enexo;
  assign act_mem_banks_read_read_data_and_23_enex5 = act_mem_banks_read_read_data_and_cse
      & reg_act_mem_banks_read_for_mux_8_enexo;
  assign act_mem_banks_read_read_data_and_24_enex5 = act_mem_banks_read_read_data_and_cse
      & reg_act_mem_banks_read_for_mux_7_enexo;
  assign act_mem_banks_read_read_data_and_25_enex5 = act_mem_banks_read_read_data_and_cse
      & reg_act_mem_banks_read_for_mux_6_enexo;
  assign act_mem_banks_read_read_data_and_26_enex5 = act_mem_banks_read_read_data_and_cse
      & reg_act_mem_banks_read_for_mux_5_enexo;
  assign act_mem_banks_read_read_data_and_27_enex5 = act_mem_banks_read_read_data_and_cse
      & reg_act_mem_banks_read_for_mux_4_enexo;
  assign act_mem_banks_read_read_data_and_28_enex5 = act_mem_banks_read_read_data_and_cse
      & reg_act_mem_banks_read_for_mux_3_enexo;
  assign act_mem_banks_read_read_data_and_29_enex5 = act_mem_banks_read_read_data_and_cse
      & reg_act_mem_banks_read_for_mux_2_enexo;
  assign act_mem_banks_read_read_data_and_30_enex5 = act_mem_banks_read_read_data_and_cse
      & reg_act_mem_banks_read_for_mux_1_enexo;
  assign act_mem_banks_read_read_data_and_31_enex5 = act_mem_banks_read_read_data_and_cse
      & reg_act_mem_banks_read_for_mux_enexo;
  assign act_port_read_out_data_and_cse = ActUnitRun_wen & and_dcpl_1109 & and_dcpl_1106;
  assign act_port_read_out_data_and_16_enex5 = act_port_read_out_data_and_cse & (reg_act_write_req_valid_lpi_1_dfm_5_enexo
      | reg_act_mem_banks_read_read_data_lpi_1_dfm_1_31_0_enexo | reg_act_mem_banks_read_for_mux_15_enexo_1);
  assign act_port_read_out_data_and_17_enex5 = act_port_read_out_data_and_cse & (reg_act_mem_banks_read_for_mux_14_enexo_1
      | reg_act_mem_banks_read_read_data_lpi_1_dfm_1_63_32_enexo | reg_act_write_req_valid_lpi_1_dfm_5_enexo_1);
  assign act_port_read_out_data_and_18_enex5 = act_port_read_out_data_and_cse & (reg_act_mem_banks_read_for_mux_13_enexo_1
      | reg_act_write_req_valid_lpi_1_dfm_5_enexo_2 | reg_act_mem_banks_read_read_data_lpi_1_dfm_1_95_64_enexo);
  assign act_port_read_out_data_and_19_enex5 = act_port_read_out_data_and_cse & (reg_act_write_req_valid_lpi_1_dfm_5_enexo_3
      | reg_act_mem_banks_read_for_mux_12_enexo_1 | reg_act_mem_banks_read_read_data_lpi_1_dfm_1_127_96_enexo);
  assign act_port_read_out_data_and_20_enex5 = act_port_read_out_data_and_cse & (reg_act_mem_banks_read_for_mux_11_enexo_1
      | reg_act_mem_banks_read_read_data_lpi_1_dfm_1_159_128_enexo | reg_act_write_req_valid_lpi_1_dfm_5_enexo_4);
  assign act_port_read_out_data_and_21_enex5 = act_port_read_out_data_and_cse & (reg_act_write_req_valid_lpi_1_dfm_5_enexo_5
      | reg_act_mem_banks_read_for_mux_10_enexo_1 | reg_act_mem_banks_read_read_data_lpi_1_dfm_1_191_160_enexo);
  assign act_port_read_out_data_and_22_enex5 = act_port_read_out_data_and_cse & (reg_act_write_req_valid_lpi_1_dfm_5_enexo_6
      | reg_act_mem_banks_read_for_mux_9_enexo_1 | reg_act_mem_banks_read_read_data_lpi_1_dfm_1_223_192_enexo);
  assign act_port_read_out_data_and_23_enex5 = act_port_read_out_data_and_cse & (reg_act_write_req_valid_lpi_1_dfm_5_enexo_7
      | reg_act_mem_banks_read_read_data_lpi_1_dfm_1_255_224_enexo | reg_act_mem_banks_read_for_mux_8_enexo_1);
  assign act_port_read_out_data_and_24_enex5 = act_port_read_out_data_and_cse & (reg_act_write_req_valid_lpi_1_dfm_5_enexo_8
      | reg_act_mem_banks_read_for_mux_7_enexo_1 | reg_act_mem_banks_read_read_data_lpi_1_dfm_1_287_256_enexo);
  assign act_port_read_out_data_and_25_enex5 = act_port_read_out_data_and_cse & (reg_act_write_req_valid_lpi_1_dfm_5_enexo_9
      | reg_act_mem_banks_read_read_data_lpi_1_dfm_1_319_288_enexo | reg_act_mem_banks_read_for_mux_6_enexo_1);
  assign act_port_read_out_data_and_26_enex5 = act_port_read_out_data_and_cse & (reg_act_mem_banks_read_for_mux_5_enexo_1
      | reg_act_write_req_valid_lpi_1_dfm_5_enexo_10 | reg_act_mem_banks_read_read_data_lpi_1_dfm_1_351_320_enexo);
  assign act_port_read_out_data_and_27_enex5 = act_port_read_out_data_and_cse & (reg_act_mem_banks_read_read_data_lpi_1_dfm_1_383_352_enexo
      | reg_act_mem_banks_read_for_mux_4_enexo_1 | reg_act_write_req_valid_lpi_1_dfm_5_enexo_11);
  assign act_port_read_out_data_and_28_enex5 = act_port_read_out_data_and_cse & (reg_act_write_req_valid_lpi_1_dfm_5_enexo_12
      | reg_act_mem_banks_read_read_data_lpi_1_dfm_1_415_384_enexo | reg_act_mem_banks_read_for_mux_3_enexo_1);
  assign act_port_read_out_data_and_29_enex5 = act_port_read_out_data_and_cse & (reg_act_mem_banks_read_read_data_lpi_1_dfm_1_447_416_enexo
      | reg_act_mem_banks_read_for_mux_2_enexo_1 | reg_act_write_req_valid_lpi_1_dfm_5_enexo_13);
  assign act_port_read_out_data_and_30_enex5 = act_port_read_out_data_and_cse & (reg_act_mem_banks_read_read_data_lpi_1_dfm_1_479_448_enexo
      | reg_act_mem_banks_read_for_mux_1_enexo_1 | reg_act_write_req_valid_lpi_1_dfm_5_enexo_14);
  assign act_port_read_out_data_and_31_enex5 = act_port_read_out_data_and_cse & (reg_act_mem_banks_read_for_mux_enexo_1
      | reg_act_write_req_valid_lpi_1_dfm_5_enexo_15 | reg_act_mem_banks_read_read_data_lpi_1_dfm_1_511_480_enexo);
  assign nor_1441_cse = ~((fsm_output[3:2]!=2'b00));
  assign Tanh_for_and_85_m1c = w_axi_rsp_lpi_1_dfm_1 & and_dcpl_1085;
  assign Tanh_for_or_cse = and_dcpl_1083 | ((~ w_axi_rsp_lpi_1_dfm_1) & and_dcpl_1085)
      | ((~ act_read_req_valid_lpi_1_dfm_6) & Tanh_for_and_85_m1c);
  assign Tanh_for_and_87_cse = act_read_req_valid_lpi_1_dfm_6 & Tanh_for_and_85_m1c;
  assign mux_438_cse = MUX_s_1_2_2(and_2371_cse, or_1872_cse, fsm_output[2]);
  assign mux_439_nl = MUX_s_1_2_2(mux_438_cse, or_dcpl_586, fsm_output[3]);
  assign ActUnit_PushOutput_if_for_and_28_cse = ActUnitRun_wen & mux_439_nl;
  assign or_1579_cse = (fsm_output[3:2]!=2'b10);
  assign nor_1442_nl = ~((fsm_output[2:0]!=3'b011) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11:8]!=4'b1000));
  assign and_2332_nl = act_read_req_valid_lpi_1_dfm_6 & w_axi_rsp_lpi_1_dfm_1 & (fsm_output[1:0]==2'b10);
  assign nor_1443_nl = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11:8]!=4'b1000));
  assign mux_629_nl = MUX_s_1_2_2(and_2332_nl, nor_1443_nl, fsm_output[2]);
  assign mux_630_nl = MUX_s_1_2_2(nor_1442_nl, mux_629_nl, fsm_output[3]);
  assign nor_1444_nl = ~((fsm_output[3:2]!=2'b10) | (~ act_read_req_valid_lpi_1_dfm_6)
      | (~ w_axi_rsp_lpi_1_dfm_1) | (fsm_output[1:0]!=2'b10));
  assign or_1582_nl = is_start_sva | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt) | rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  assign mux_631_nl = MUX_s_1_2_2(mux_630_nl, nor_1444_nl, or_1582_nl);
  assign and_1809_cse = mux_631_nl & ActUnitRun_wen;
  assign mux_441_nl = MUX_s_1_2_2(and_dcpl_1077, (fsm_output[2]), fsm_output[3]);
  assign or_1306_nl = (fsm_output[2]) | and_dcpl_848;
  assign mux_440_nl = MUX_s_1_2_2(and_dcpl_1077, or_1306_nl, fsm_output[3]);
  assign and_1647_nl = act_read_req_valid_lpi_1_dfm_6 & w_axi_rsp_lpi_1_dfm_1;
  assign mux_442_nl = MUX_s_1_2_2(mux_441_nl, mux_440_nl, and_1647_nl);
  assign rva_out_reg_data_and_15_cse = ActUnitRun_wen & ((~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11:9]!=3'b100)
      | or_dcpl_465 | is_start_sva | (~ mux_442_nl))) | and_dcpl_1094);
  assign mux_443_nl = MUX_s_1_2_2((fsm_output[1]), (~ or_1872_cse), fsm_output[2]);
  assign ActUnit_RunInst_switch_lp_and_802_cse = ActUnitRun_wen & (~(mux_443_nl &
      (~ (fsm_output[3]))));
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc = ActUnit_RunInst_switch_lp_and_802_cse
      & is_start_sva & (~ (act_config_in_InstFetch_mux_tmp[7])) & (act_config_in_InstFetch_mux_tmp[5])
      & and_dcpl_78;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_37_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo | reg_act_config_inst_regs_4_sva_dfm_5_enexo
      | reg_act_regs_data_3_15_1_enexo | reg_act_config_inst_counter_enexo | reg_act_regs_data_2_15_1_enexo
      | reg_act_regs_data_0_15_1_enexo | reg_act_regs_data_1_15_1_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_38_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_1 | reg_act_regs_data_0_15_2_enexo
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_1 | reg_act_regs_data_1_15_2_enexo
      | reg_act_regs_data_2_15_2_enexo | reg_act_regs_data_3_15_2_enexo | reg_act_config_inst_counter_enexo_1);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_39_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_2 | reg_act_regs_data_1_15_3_enexo
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_2 | reg_act_regs_data_0_15_3_enexo
      | reg_act_config_inst_counter_enexo_2 | reg_act_regs_data_3_15_3_enexo | reg_act_regs_data_2_15_3_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_40_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_3 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_3
      | reg_act_regs_data_2_14_1_enexo | reg_act_regs_data_1_14_1_enexo | reg_act_regs_data_0_14_1_enexo
      | reg_act_config_inst_counter_enexo_3 | reg_act_regs_data_3_14_1_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_41_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_4 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_4
      | reg_act_regs_data_2_14_2_enexo | reg_act_regs_data_1_14_2_enexo | reg_act_config_inst_counter_enexo_4
      | reg_act_regs_data_3_14_2_enexo | reg_act_regs_data_0_14_2_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_42_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_5 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_5
      | reg_act_regs_data_1_14_3_enexo | reg_act_config_inst_counter_enexo_5 | reg_act_regs_data_2_14_3_enexo
      | reg_act_regs_data_0_14_3_enexo | reg_act_regs_data_3_14_3_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_43_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_6 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_6
      | reg_act_regs_data_1_13_1_enexo | reg_act_regs_data_2_13_1_enexo | reg_act_regs_data_3_13_1_enexo
      | reg_act_regs_data_0_13_1_enexo | reg_act_config_inst_counter_enexo_6);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_44_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_7 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_7
      | reg_act_config_inst_counter_enexo_7 | reg_act_regs_data_1_13_2_enexo | reg_act_regs_data_0_13_2_enexo
      | reg_act_regs_data_2_13_2_enexo | reg_act_regs_data_3_13_2_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_45_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_8 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_8
      | reg_act_regs_data_3_13_3_enexo | reg_act_config_inst_counter_enexo_8 | reg_act_regs_data_0_13_3_enexo
      | reg_act_regs_data_2_13_3_enexo | reg_act_regs_data_1_13_3_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_46_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_9 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_9
      | reg_act_regs_data_0_12_1_enexo | reg_act_regs_data_3_12_1_enexo | reg_act_regs_data_1_12_1_enexo
      | reg_act_config_inst_counter_enexo_9 | reg_act_regs_data_2_12_1_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_47_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_10 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_10
      | reg_act_regs_data_3_12_2_enexo | reg_act_regs_data_2_12_2_enexo | reg_act_regs_data_0_12_2_enexo
      | reg_act_regs_data_1_12_2_enexo | reg_act_config_inst_counter_enexo_10);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_48_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_regs_data_3_12_3_enexo | reg_act_config_inst_regs_4_sva_dfm_5_enexo_11
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_11 | reg_act_config_inst_counter_enexo_11
      | reg_act_regs_data_1_12_3_enexo | reg_act_regs_data_0_12_3_enexo | reg_act_regs_data_2_12_3_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_49_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_counter_enexo_12 | reg_act_regs_data_1_11_1_enexo |
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_12 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_12
      | reg_act_regs_data_2_11_1_enexo | reg_act_regs_data_3_11_1_enexo | reg_act_regs_data_0_11_1_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_50_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_13 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_13
      | reg_act_config_inst_counter_enexo_13 | reg_act_regs_data_2_11_2_enexo | reg_act_regs_data_3_11_2_enexo
      | reg_act_regs_data_1_11_2_enexo | reg_act_regs_data_0_11_2_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_51_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_14 | reg_act_config_inst_counter_enexo_14
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_14 | reg_act_regs_data_2_11_3_enexo
      | reg_act_regs_data_1_11_3_enexo | reg_act_regs_data_3_11_3_enexo | reg_act_regs_data_0_11_3_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_52_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_15 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_15
      | reg_act_config_inst_counter_enexo_15 | reg_act_regs_data_1_10_1_enexo | reg_act_regs_data_0_10_1_enexo
      | reg_act_regs_data_2_10_1_enexo | reg_act_regs_data_3_10_1_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_53_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_16 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_16
      | reg_act_regs_data_2_10_2_enexo | reg_act_regs_data_0_10_2_enexo | reg_act_config_inst_counter_enexo_16
      | reg_act_regs_data_1_10_2_enexo | reg_act_regs_data_3_10_2_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_54_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_17 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_17
      | reg_act_regs_data_1_10_3_enexo | reg_act_regs_data_3_10_3_enexo | reg_act_regs_data_0_10_3_enexo
      | reg_act_regs_data_2_10_3_enexo | reg_act_config_inst_counter_enexo_17);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_55_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_18 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_18
      | reg_act_regs_data_3_9_1_enexo | reg_act_regs_data_1_9_1_enexo | reg_act_config_inst_counter_enexo_18
      | reg_act_regs_data_2_9_1_enexo | reg_act_regs_data_0_9_1_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_56_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_regs_data_3_9_2_enexo | reg_act_config_inst_regs_20_sva_dfm_6_enexo_19
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_19 | reg_act_regs_data_0_9_2_enexo
      | reg_act_regs_data_2_9_2_enexo | reg_act_config_inst_counter_enexo_19 | reg_act_regs_data_1_9_2_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_57_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_regs_data_0_9_3_enexo | reg_act_config_inst_regs_4_sva_dfm_5_enexo_20
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_20 | reg_act_regs_data_2_9_3_enexo
      | reg_act_regs_data_3_9_3_enexo | reg_act_config_inst_counter_enexo_20 | reg_act_regs_data_1_9_3_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_58_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_21 | reg_act_config_inst_counter_enexo_21
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_21 | reg_act_regs_data_3_8_1_enexo
      | reg_act_regs_data_0_8_1_enexo | reg_act_regs_data_2_8_1_enexo | reg_act_regs_data_1_8_1_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_59_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_22 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_22
      | reg_act_regs_data_2_8_2_enexo | reg_act_regs_data_1_8_2_enexo | reg_act_regs_data_0_8_2_enexo
      | reg_act_regs_data_3_8_2_enexo | reg_act_config_inst_counter_enexo_22);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_60_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_23 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_23
      | reg_act_regs_data_3_8_3_enexo | reg_act_regs_data_0_8_3_enexo | reg_act_regs_data_2_8_3_enexo
      | reg_act_config_inst_counter_enexo_23 | reg_act_regs_data_1_8_3_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_61_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_24 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_24
      | reg_act_regs_data_0_7_1_enexo | reg_act_config_inst_counter_enexo_24 | reg_act_regs_data_2_7_1_enexo
      | reg_act_regs_data_1_7_1_enexo | reg_act_regs_data_3_7_1_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_62_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_25 | reg_act_config_inst_counter_enexo_25
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_25 | reg_act_regs_data_3_7_2_enexo
      | reg_act_regs_data_1_7_2_enexo | reg_act_regs_data_0_7_2_enexo | reg_act_regs_data_2_7_2_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_63_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_26 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_26
      | reg_act_regs_data_1_7_3_enexo | reg_act_regs_data_3_7_3_enexo | reg_act_config_inst_counter_enexo_26
      | reg_act_regs_data_0_7_3_enexo | reg_act_regs_data_2_7_3_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_64_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_27 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_27
      | reg_act_regs_data_0_6_1_enexo | reg_act_config_inst_counter_enexo_27 | reg_act_regs_data_1_6_1_enexo
      | reg_act_regs_data_3_6_1_enexo | reg_act_regs_data_2_6_1_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_65_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_28 | reg_act_regs_data_1_6_2_enexo
      | reg_act_regs_data_3_6_2_enexo | reg_act_config_inst_regs_4_sva_dfm_5_enexo_28
      | reg_act_config_inst_counter_enexo_28 | reg_act_regs_data_2_6_2_enexo | reg_act_regs_data_0_6_2_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_66_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_29 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_29
      | reg_act_regs_data_2_6_3_enexo | reg_act_regs_data_1_6_3_enexo | reg_act_config_inst_counter_enexo_29
      | reg_act_regs_data_3_6_3_enexo | reg_act_regs_data_0_6_3_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_67_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_30 | reg_act_regs_data_3_5_1_enexo
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_30 | reg_act_config_inst_counter_enexo_30
      | reg_act_regs_data_2_5_1_enexo | reg_act_regs_data_0_5_1_enexo | reg_act_regs_data_1_5_1_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_68_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_regs_data_3_5_2_enexo | reg_act_config_inst_regs_20_sva_dfm_6_enexo_31
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_31 | reg_act_regs_data_1_5_2_enexo
      | reg_act_config_inst_counter_enexo_31 | reg_act_regs_data_2_5_2_enexo | reg_act_regs_data_0_5_2_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_69_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_32 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_32
      | reg_act_config_inst_counter_enexo_32 | reg_act_regs_data_3_5_3_enexo | reg_act_regs_data_1_5_3_enexo
      | reg_act_regs_data_0_5_3_enexo | reg_act_regs_data_2_5_3_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_70_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_regs_data_1_4_1_enexo | reg_act_config_inst_regs_20_sva_dfm_6_enexo_33
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_33 | reg_act_regs_data_3_4_1_enexo
      | reg_act_regs_data_0_4_1_enexo | reg_act_config_inst_counter_enexo_33 | reg_act_regs_data_2_4_1_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_71_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_34 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_34
      | reg_act_config_inst_counter_enexo_34 | reg_act_regs_data_1_4_2_enexo | reg_act_regs_data_0_4_2_enexo
      | reg_act_regs_data_3_4_2_enexo | reg_act_regs_data_2_4_2_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_72_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_35 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_35
      | reg_act_regs_data_2_4_3_enexo | reg_act_regs_data_1_4_3_enexo | reg_act_regs_data_0_4_3_enexo
      | reg_act_config_inst_counter_enexo_35 | reg_act_regs_data_3_4_3_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_73_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_36 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_36
      | reg_act_config_inst_counter_enexo_36 | reg_act_regs_data_2_3_1_enexo | reg_act_regs_data_3_3_1_enexo
      | reg_act_regs_data_1_3_1_enexo | reg_act_regs_data_0_3_1_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_74_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_37 | reg_act_regs_data_0_3_2_enexo
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_37 | reg_act_config_inst_counter_enexo_37
      | reg_act_regs_data_3_3_2_enexo | reg_act_regs_data_2_3_2_enexo | reg_act_regs_data_1_3_2_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_75_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_38 | reg_act_config_inst_counter_enexo_38
      | reg_act_regs_data_0_3_3_enexo | reg_act_config_inst_regs_4_sva_dfm_5_enexo_38
      | reg_act_regs_data_2_3_3_enexo | reg_act_regs_data_3_3_3_enexo | reg_act_regs_data_1_3_3_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_76_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_counter_enexo_39 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_39
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_39 | reg_act_regs_data_3_2_1_enexo
      | reg_act_regs_data_2_2_1_enexo | reg_act_regs_data_0_2_1_enexo | reg_act_regs_data_1_2_1_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_77_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_40 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_40
      | reg_act_config_inst_counter_enexo_40 | reg_act_regs_data_2_2_2_enexo | reg_act_regs_data_0_2_2_enexo
      | reg_act_regs_data_3_2_2_enexo | reg_act_regs_data_1_2_2_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_78_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_41 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_41
      | reg_act_regs_data_2_2_3_enexo | reg_act_config_inst_counter_enexo_41 | reg_act_regs_data_1_2_3_enexo
      | reg_act_regs_data_3_2_3_enexo | reg_act_regs_data_0_2_3_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_79_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_42 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_42
      | reg_act_regs_data_0_1_1_enexo | reg_act_regs_data_2_1_1_enexo | reg_act_regs_data_1_1_1_enexo
      | reg_act_regs_data_3_1_1_enexo | reg_act_config_inst_counter_enexo_42);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_80_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_43 | reg_act_regs_data_3_1_2_enexo
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_43 | reg_act_regs_data_1_1_2_enexo
      | reg_act_regs_data_2_1_2_enexo | reg_act_regs_data_0_1_2_enexo | reg_act_config_inst_counter_enexo_43);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_81_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_regs_data_2_1_3_enexo | reg_act_config_inst_regs_20_sva_dfm_6_enexo_44
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_44 | reg_act_config_inst_counter_enexo_44
      | reg_act_regs_data_1_1_3_enexo | reg_act_regs_data_3_1_3_enexo | reg_act_regs_data_0_1_3_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_82_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_regs_data_3_0_1_enexo | reg_act_config_inst_regs_20_sva_dfm_6_enexo_45
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_45 | reg_act_config_inst_counter_enexo_45
      | reg_act_regs_data_2_0_1_enexo | reg_act_regs_data_0_0_1_enexo | reg_act_regs_data_1_0_1_enexo);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_83_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_46 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_46
      | reg_act_regs_data_1_0_2_enexo | reg_act_regs_data_0_0_2_enexo | reg_act_regs_data_2_0_2_enexo
      | reg_act_regs_data_3_0_2_enexo | reg_act_config_inst_counter_enexo_46);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_84_enex5 = nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_47 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_47
      | reg_act_regs_data_0_0_3_enexo | reg_act_config_inst_counter_enexo_47 | reg_act_regs_data_3_0_3_enexo
      | reg_act_regs_data_2_0_3_enexo | reg_act_regs_data_1_0_3_enexo);
  assign Tanh_for_and_79_ssc = ($signed({1'b0, 25'b1000000000000000000000000}) <
      $signed(({nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm})))
      & (~ Tanh_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1);
  assign Tanh_for_y_and_ssc = ActUnit_RunInst_switch_lp_and_802_cse & and_dcpl_84
      & (~ (act_config_in_InstFetch_mux_tmp[6])) & (act_config_in_InstFetch_mux_tmp[4]);
  assign Tanh_for_y_and_31_enex5 = Tanh_for_y_and_ssc & (reg_act_regs_data_1_15_enexo
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_48 | reg_act_regs_data_1_15_3_enexo_1
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_48 | reg_act_regs_data_0_15_1_enexo_1
      | reg_act_config_inst_counter_enexo_48 | reg_act_regs_data_2_15_1_enexo_1 |
      reg_act_regs_data_1_15_2_enexo_1 | reg_act_regs_data_3_15_3_enexo_1 | reg_act_regs_data_3_15_2_enexo_1
      | reg_act_regs_data_3_15_1_enexo_1 | reg_act_regs_data_2_15_2_enexo_1 | reg_act_regs_data_0_15_2_enexo_1
      | reg_act_regs_data_1_15_1_enexo_1 | reg_act_regs_data_0_15_3_enexo_1 | reg_act_regs_data_2_15_3_enexo_1);
  assign Tanh_for_y_and_32_enex5 = Tanh_for_y_and_ssc & (reg_act_regs_data_1_15_enexo_1
      | reg_act_regs_data_3_15_1_enexo_2 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_49
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_49 | reg_act_regs_data_2_15_1_enexo_2
      | reg_act_regs_data_1_15_2_enexo_2 | reg_act_regs_data_0_15_3_enexo_2 | reg_act_regs_data_1_15_1_enexo_2
      | reg_act_regs_data_3_15_2_enexo_2 | reg_act_regs_data_2_15_3_enexo_2 | reg_act_regs_data_0_15_2_enexo_2
      | reg_act_regs_data_3_15_3_enexo_2 | reg_act_regs_data_1_15_3_enexo_2 | reg_act_config_inst_counter_enexo_49
      | reg_act_regs_data_0_15_1_enexo_2 | reg_act_regs_data_2_15_2_enexo_2);
  assign Tanh_for_and_77_ssc = ($signed({1'b0, 25'b1000000000000000000000000}) <
      $signed(({nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm})))
      & (~ Tanh_for_15_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1);
  assign Tanh_for_y_and_33_enex5 = Tanh_for_y_and_ssc & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_50
      | reg_act_regs_data_0_14_enexo | reg_act_regs_data_2_14_1_enexo_1 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_50
      | reg_act_regs_data_2_14_3_enexo_1 | reg_act_regs_data_1_14_1_enexo_1 | reg_act_regs_data_1_14_3_enexo_1
      | reg_act_regs_data_0_14_2_enexo_1 | reg_act_regs_data_2_14_2_enexo_1 | reg_act_regs_data_0_14_1_enexo_1
      | reg_act_regs_data_3_14_1_enexo_1 | reg_act_regs_data_3_14_3_enexo_1 | reg_act_config_inst_counter_enexo_50
      | reg_act_regs_data_3_14_2_enexo_1 | reg_act_regs_data_0_14_3_enexo_1 | reg_act_regs_data_1_14_2_enexo_1);
  assign Tanh_for_y_and_34_enex5 = Tanh_for_y_and_ssc & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_51
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_51 | reg_act_regs_data_3_14_1_enexo_2
      | reg_act_regs_data_0_14_3_enexo_2 | reg_act_regs_data_2_14_1_enexo_2 | reg_act_regs_data_1_14_3_enexo_2
      | reg_act_regs_data_0_14_enexo_1 | reg_act_regs_data_3_14_3_enexo_2 | reg_act_config_inst_counter_enexo_51
      | reg_act_regs_data_0_14_2_enexo_2 | reg_act_regs_data_1_14_1_enexo_2 | reg_act_regs_data_1_14_2_enexo_2
      | reg_act_regs_data_0_14_1_enexo_2 | reg_act_regs_data_2_14_3_enexo_2 | reg_act_regs_data_3_14_2_enexo_2
      | reg_act_regs_data_2_14_2_enexo_2);
  assign Tanh_for_and_75_ssc = ($signed({1'b0, 25'b1000000000000000000000000}) <
      $signed(({nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm})))
      & (~ Tanh_for_14_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1);
  assign Tanh_for_y_and_35_enex5 = Tanh_for_y_and_ssc & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_52
      | reg_act_regs_data_2_13_2_enexo_1 | reg_act_regs_data_3_13_2_enexo_1 | reg_act_regs_data_0_13_1_enexo_1
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_52 | reg_act_regs_data_3_13_3_enexo_1
      | reg_act_regs_data_1_13_3_enexo_1 | reg_act_config_inst_counter_enexo_52 |
      reg_act_regs_data_0_13_3_enexo_1 | reg_act_regs_data_3_13_enexo | reg_act_regs_data_0_13_2_enexo_1
      | reg_act_regs_data_2_13_3_enexo_1 | reg_act_regs_data_3_13_1_enexo_1 | reg_act_regs_data_1_13_2_enexo_1
      | reg_act_regs_data_2_13_1_enexo_1 | reg_act_regs_data_1_13_1_enexo_1);
  assign Tanh_for_y_and_36_enex5 = Tanh_for_y_and_ssc & (reg_act_config_inst_counter_enexo_53
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_53 | reg_act_regs_data_0_13_1_enexo_2
      | reg_act_regs_data_3_13_enexo_1 | reg_act_regs_data_3_13_1_enexo_2 | reg_act_regs_data_2_13_2_enexo_2
      | reg_act_regs_data_1_13_2_enexo_2 | reg_act_regs_data_3_13_3_enexo_2 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_53
      | reg_act_regs_data_1_13_1_enexo_2 | reg_act_regs_data_0_13_2_enexo_2 | reg_act_regs_data_1_13_3_enexo_2
      | reg_act_regs_data_2_13_3_enexo_2 | reg_act_regs_data_3_13_2_enexo_2 | reg_act_regs_data_2_13_1_enexo_2
      | reg_act_regs_data_0_13_3_enexo_2);
  assign Tanh_for_and_73_ssc = ($signed({1'b0, 25'b1000000000000000000000000}) <
      $signed(({nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm})))
      & (~ Tanh_for_13_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1);
  assign Tanh_for_y_and_37_enex5 = Tanh_for_y_and_ssc & (reg_act_regs_data_2_12_1_enexo_1
      | reg_act_regs_data_3_12_3_enexo_1 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_54
      | reg_act_regs_data_1_12_1_enexo_1 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_54
      | reg_act_regs_data_0_12_enexo | reg_act_regs_data_0_12_2_enexo_1 | reg_act_regs_data_1_12_3_enexo_1
      | reg_act_regs_data_2_12_2_enexo_1 | reg_act_regs_data_3_12_1_enexo_1 | reg_act_config_inst_counter_enexo_54
      | reg_act_regs_data_1_12_2_enexo_1 | reg_act_regs_data_2_12_3_enexo_1 | reg_act_regs_data_0_12_3_enexo_1
      | reg_act_regs_data_3_12_2_enexo_1 | reg_act_regs_data_0_12_1_enexo_1);
  assign Tanh_for_y_and_38_enex5 = Tanh_for_y_and_ssc & (reg_act_regs_data_0_12_enexo_1
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_55 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_55
      | reg_act_regs_data_0_12_1_enexo_2 | reg_act_regs_data_1_12_2_enexo_2 | reg_act_regs_data_1_12_1_enexo_2
      | reg_act_regs_data_0_12_2_enexo_2 | reg_act_regs_data_3_12_2_enexo_2 | reg_act_regs_data_2_12_1_enexo_2
      | reg_act_regs_data_2_12_2_enexo_2 | reg_act_regs_data_3_12_1_enexo_2 | reg_act_regs_data_2_12_3_enexo_2
      | reg_act_config_inst_counter_enexo_55 | reg_act_regs_data_0_12_3_enexo_2 |
      reg_act_regs_data_1_12_3_enexo_2 | reg_act_regs_data_3_12_3_enexo_2);
  assign Tanh_for_and_71_ssc = ($signed({1'b0, 25'b1000000000000000000000000}) <
      $signed(({nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm})))
      & (~ Tanh_for_12_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1);
  assign Tanh_for_y_and_39_enex5 = Tanh_for_y_and_ssc & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_56
      | reg_act_config_inst_counter_enexo_56 | reg_act_regs_data_2_11_enexo | reg_act_regs_data_1_11_3_enexo_1
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_56 | reg_act_regs_data_3_11_3_enexo_1
      | reg_act_regs_data_2_11_2_enexo_1 | reg_act_regs_data_1_11_1_enexo_1 | reg_act_regs_data_0_11_1_enexo_1
      | reg_act_regs_data_2_11_1_enexo_1 | reg_act_regs_data_3_11_1_enexo_1 | reg_act_regs_data_2_11_3_enexo_1
      | reg_act_regs_data_3_11_2_enexo_1 | reg_act_regs_data_1_11_2_enexo_1 | reg_act_regs_data_0_11_3_enexo_1
      | reg_act_regs_data_0_11_2_enexo_1);
  assign Tanh_for_y_and_40_enex5 = Tanh_for_y_and_ssc & (reg_act_regs_data_1_11_2_enexo_2
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_57 | reg_act_regs_data_1_11_3_enexo_2
      | reg_act_regs_data_2_11_enexo_1 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_57
      | reg_act_regs_data_3_11_2_enexo_2 | reg_act_regs_data_2_11_3_enexo_2 | reg_act_regs_data_3_11_3_enexo_2
      | reg_act_regs_data_0_11_2_enexo_2 | reg_act_regs_data_3_11_1_enexo_2 | reg_act_regs_data_2_11_1_enexo_2
      | reg_act_config_inst_counter_enexo_57 | reg_act_regs_data_2_11_2_enexo_2 |
      reg_act_regs_data_0_11_1_enexo_2 | reg_act_regs_data_0_11_3_enexo_2 | reg_act_regs_data_1_11_1_enexo_2);
  assign Tanh_for_and_69_ssc = ($signed({1'b0, 25'b1000000000000000000000000}) <
      $signed(({nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm})))
      & (~ Tanh_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1);
  assign Tanh_for_y_and_41_enex5 = Tanh_for_y_and_ssc & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_58
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_58 | reg_act_regs_data_0_10_2_enexo_1
      | reg_act_regs_data_1_10_3_enexo_1 | reg_act_regs_data_0_10_3_enexo_1 | reg_act_regs_data_0_10_enexo
      | reg_act_regs_data_2_10_1_enexo_1 | reg_act_regs_data_3_10_3_enexo_1 | reg_act_regs_data_1_10_1_enexo_1
      | reg_act_regs_data_3_10_2_enexo_1 | reg_act_regs_data_0_10_1_enexo_1 | reg_act_regs_data_2_10_2_enexo_1
      | reg_act_regs_data_3_10_1_enexo_1 | reg_act_regs_data_2_10_3_enexo_1 | reg_act_regs_data_1_10_2_enexo_1
      | reg_act_config_inst_counter_enexo_58);
  assign Tanh_for_y_and_42_enex5 = Tanh_for_y_and_ssc & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_59
      | reg_act_regs_data_1_10_1_enexo_2 | reg_act_regs_data_0_10_2_enexo_2 | reg_act_regs_data_0_10_3_enexo_2
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_59 | reg_act_regs_data_1_10_2_enexo_2
      | reg_act_regs_data_0_10_1_enexo_2 | reg_act_regs_data_2_10_3_enexo_2 | reg_act_regs_data_3_10_2_enexo_2
      | reg_act_config_inst_counter_enexo_59 | reg_act_regs_data_0_10_enexo_1 | reg_act_regs_data_1_10_3_enexo_2
      | reg_act_regs_data_3_10_3_enexo_2 | reg_act_regs_data_2_10_1_enexo_2 | reg_act_regs_data_3_10_1_enexo_2
      | reg_act_regs_data_2_10_2_enexo_2);
  assign Tanh_for_and_67_ssc = ($signed({1'b0, 25'b1000000000000000000000000}) <
      $signed(({nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm})))
      & (~ Tanh_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1);
  assign Tanh_for_y_and_43_enex5 = Tanh_for_y_and_ssc & (reg_act_regs_data_3_9_3_enexo_1
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_60 | reg_act_regs_data_2_9_2_enexo_1
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_60 | reg_act_regs_data_2_9_3_enexo_1
      | reg_act_regs_data_1_9_2_enexo_1 | reg_act_regs_data_0_9_2_enexo_1 | reg_act_config_inst_counter_enexo_60
      | reg_act_regs_data_1_9_1_enexo_1 | reg_act_regs_data_0_9_3_enexo_1 | reg_act_regs_data_1_9_enexo
      | reg_act_regs_data_2_9_1_enexo_1 | reg_act_regs_data_1_9_3_enexo_1 | reg_act_regs_data_0_9_1_enexo_1
      | reg_act_regs_data_3_9_1_enexo_1 | reg_act_regs_data_3_9_2_enexo_1);
  assign Tanh_for_y_and_44_enex5 = Tanh_for_y_and_ssc & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_61
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_61 | reg_act_regs_data_2_9_3_enexo_2
      | reg_act_regs_data_0_9_1_enexo_2 | reg_act_regs_data_3_9_1_enexo_2 | reg_act_regs_data_2_9_1_enexo_2
      | reg_act_regs_data_1_9_3_enexo_2 | reg_act_regs_data_1_9_enexo_1 | reg_act_regs_data_0_9_2_enexo_2
      | reg_act_regs_data_0_9_3_enexo_2 | reg_act_regs_data_3_9_2_enexo_2 | reg_act_regs_data_3_9_3_enexo_2
      | reg_act_regs_data_1_9_2_enexo_2 | reg_act_regs_data_2_9_2_enexo_2 | reg_act_regs_data_1_9_1_enexo_2
      | reg_act_config_inst_counter_enexo_61);
  assign Tanh_for_and_65_ssc = ($signed({1'b0, 25'b1000000000000000000000000}) <
      $signed(({nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm})))
      & (~ Tanh_for_9_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1);
  assign Tanh_for_y_and_45_enex5 = Tanh_for_y_and_ssc & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_62
      | reg_act_regs_data_2_8_enexo | reg_act_regs_data_0_8_2_enexo_1 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_62
      | reg_act_regs_data_0_8_3_enexo_1 | reg_act_regs_data_0_8_1_enexo_1 | reg_act_regs_data_3_8_1_enexo_1
      | reg_act_regs_data_2_8_1_enexo_1 | reg_act_regs_data_3_8_2_enexo_1 | reg_act_regs_data_2_8_3_enexo_1
      | reg_act_config_inst_counter_enexo_62 | reg_act_regs_data_1_8_1_enexo_1 |
      reg_act_regs_data_1_8_3_enexo_1 | reg_act_regs_data_2_8_2_enexo_1 | reg_act_regs_data_3_8_3_enexo_1
      | reg_act_regs_data_1_8_2_enexo_1);
  assign Tanh_for_y_and_46_enex5 = Tanh_for_y_and_ssc & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_63
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_63 | reg_act_regs_data_0_8_1_enexo_2
      | reg_act_regs_data_1_8_2_enexo_2 | reg_act_regs_data_3_8_3_enexo_2 | reg_act_regs_data_0_8_3_enexo_2
      | reg_act_regs_data_2_8_enexo_1 | reg_act_regs_data_2_8_1_enexo_2 | reg_act_config_inst_counter_enexo_63
      | reg_act_regs_data_3_8_1_enexo_2 | reg_act_regs_data_0_8_2_enexo_2 | reg_act_regs_data_3_8_2_enexo_2
      | reg_act_regs_data_2_8_3_enexo_2 | reg_act_regs_data_2_8_2_enexo_2 | reg_act_regs_data_1_8_1_enexo_2
      | reg_act_regs_data_1_8_3_enexo_2);
  assign Tanh_for_and_63_ssc = ($signed({1'b0, 25'b1000000000000000000000000}) <
      $signed(({nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm})))
      & (~ Tanh_for_8_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1);
  assign Tanh_for_y_and_47_enex5 = Tanh_for_y_and_ssc & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_64
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_64 | reg_act_regs_data_2_7_2_enexo_1
      | reg_act_regs_data_2_7_1_enexo_1 | reg_act_regs_data_1_7_enexo | reg_act_regs_data_2_7_3_enexo_1
      | reg_act_regs_data_1_7_2_enexo_1 | reg_act_regs_data_3_7_1_enexo_1 | reg_act_regs_data_1_7_1_enexo_1
      | reg_act_regs_data_0_7_1_enexo_1 | reg_act_regs_data_0_7_2_enexo_1 | reg_act_regs_data_3_7_2_enexo_1
      | reg_act_regs_data_3_7_3_enexo_1 | reg_act_regs_data_1_7_3_enexo_1 | reg_act_config_inst_counter_enexo_64
      | reg_act_regs_data_0_7_3_enexo_1);
  assign Tanh_for_y_and_48_enex5 = Tanh_for_y_and_ssc & (reg_act_config_inst_counter_enexo_65
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_65 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_65
      | reg_act_regs_data_2_7_1_enexo_2 | reg_act_regs_data_3_7_3_enexo_2 | reg_act_regs_data_0_7_1_enexo_2
      | reg_act_regs_data_2_7_3_enexo_2 | reg_act_regs_data_1_7_2_enexo_2 | reg_act_regs_data_1_7_enexo_1
      | reg_act_regs_data_1_7_3_enexo_2 | reg_act_regs_data_3_7_2_enexo_2 | reg_act_regs_data_3_7_1_enexo_2
      | reg_act_regs_data_0_7_2_enexo_2 | reg_act_regs_data_2_7_2_enexo_2 | reg_act_regs_data_0_7_3_enexo_2
      | reg_act_regs_data_1_7_1_enexo_2);
  assign Tanh_for_and_61_ssc = ($signed({1'b0, 25'b1000000000000000000000000}) <
      $signed(({nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm})))
      & (~ Tanh_for_7_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1);
  assign Tanh_for_y_and_49_enex5 = Tanh_for_y_and_ssc & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_66
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_66 | reg_act_regs_data_3_6_1_enexo_1
      | reg_act_config_inst_counter_enexo_66 | reg_act_regs_data_3_6_enexo | reg_act_regs_data_0_6_1_enexo_1
      | reg_act_regs_data_1_6_1_enexo_1 | reg_act_regs_data_2_6_1_enexo_1 | reg_act_regs_data_1_6_3_enexo_1
      | reg_act_regs_data_2_6_2_enexo_1 | reg_act_regs_data_1_6_2_enexo_1 | reg_act_regs_data_2_6_3_enexo_1
      | reg_act_regs_data_0_6_3_enexo_1 | reg_act_regs_data_3_6_3_enexo_1 | reg_act_regs_data_0_6_2_enexo_1
      | reg_act_regs_data_3_6_2_enexo_1);
  assign Tanh_for_y_and_50_enex5 = Tanh_for_y_and_ssc & (reg_act_regs_data_3_6_enexo_1
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_67 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_67
      | reg_act_regs_data_0_6_1_enexo_2 | reg_act_regs_data_1_6_2_enexo_2 | reg_act_regs_data_2_6_2_enexo_2
      | reg_act_regs_data_0_6_3_enexo_2 | reg_act_regs_data_1_6_3_enexo_2 | reg_act_config_inst_counter_enexo_67
      | reg_act_regs_data_2_6_1_enexo_2 | reg_act_regs_data_3_6_2_enexo_2 | reg_act_regs_data_0_6_2_enexo_2
      | reg_act_regs_data_3_6_3_enexo_2 | reg_act_regs_data_3_6_1_enexo_2 | reg_act_regs_data_1_6_1_enexo_2
      | reg_act_regs_data_2_6_3_enexo_2);
  assign Tanh_for_and_59_ssc = ($signed({1'b0, 25'b1000000000000000000000000}) <
      $signed(({nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm})))
      & (~ Tanh_for_6_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1);
  assign Tanh_for_y_and_51_enex5 = Tanh_for_y_and_ssc & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_68
      | reg_act_regs_data_3_5_2_enexo_1 | reg_act_regs_data_3_5_1_enexo_1 | reg_act_regs_data_2_5_1_enexo_1
      | reg_act_regs_data_3_5_3_enexo_1 | reg_act_regs_data_1_5_enexo | reg_act_config_inst_regs_20_sva_dfm_6_enexo_68
      | reg_act_regs_data_0_5_3_enexo_1 | reg_act_regs_data_1_5_2_enexo_1 | reg_act_regs_data_2_5_2_enexo_1
      | reg_act_regs_data_2_5_3_enexo_1 | reg_act_regs_data_0_5_1_enexo_1 | reg_act_config_inst_counter_enexo_68
      | reg_act_regs_data_0_5_2_enexo_1 | reg_act_regs_data_1_5_1_enexo_1 | reg_act_regs_data_1_5_3_enexo_1);
  assign Tanh_for_y_and_52_enex5 = Tanh_for_y_and_ssc & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_69
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_69 | reg_act_regs_data_1_5_enexo_1
      | reg_act_regs_data_1_5_3_enexo_2 | reg_act_regs_data_3_5_1_enexo_2 | reg_act_regs_data_0_5_2_enexo_2
      | reg_act_regs_data_1_5_2_enexo_2 | reg_act_regs_data_2_5_2_enexo_2 | reg_act_regs_data_2_5_3_enexo_2
      | reg_act_regs_data_0_5_3_enexo_2 | reg_act_config_inst_counter_enexo_69 |
      reg_act_regs_data_2_5_1_enexo_2 | reg_act_regs_data_3_5_3_enexo_2 | reg_act_regs_data_3_5_2_enexo_2
      | reg_act_regs_data_0_5_1_enexo_2 | reg_act_regs_data_1_5_1_enexo_2);
  assign Tanh_for_and_57_ssc = ($signed({1'b0, 25'b1000000000000000000000000}) <
      $signed(({nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm})))
      & (~ Tanh_for_5_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1);
  assign Tanh_for_y_and_53_enex5 = Tanh_for_y_and_ssc & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_70
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_70 | reg_act_regs_data_3_4_enexo
      | reg_act_regs_data_0_4_2_enexo_1 | reg_act_regs_data_2_4_3_enexo_1 | reg_act_regs_data_1_4_2_enexo_1
      | reg_act_regs_data_3_4_2_enexo_1 | reg_act_regs_data_2_4_2_enexo_1 | reg_act_regs_data_0_4_1_enexo_1
      | reg_act_regs_data_3_4_3_enexo_1 | reg_act_regs_data_1_4_1_enexo_1 | reg_act_regs_data_0_4_3_enexo_1
      | reg_act_regs_data_1_4_3_enexo_1 | reg_act_regs_data_2_4_1_enexo_1 | reg_act_regs_data_3_4_1_enexo_1
      | reg_act_config_inst_counter_enexo_70);
  assign Tanh_for_y_and_54_enex5 = Tanh_for_y_and_ssc & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_71
      | reg_act_regs_data_3_4_enexo_1 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_71
      | reg_act_regs_data_2_4_1_enexo_2 | reg_act_regs_data_2_4_3_enexo_2 | reg_act_config_inst_counter_enexo_71
      | reg_act_regs_data_1_4_1_enexo_2 | reg_act_regs_data_3_4_1_enexo_2 | reg_act_regs_data_1_4_2_enexo_2
      | reg_act_regs_data_1_4_3_enexo_2 | reg_act_regs_data_0_4_3_enexo_2 | reg_act_regs_data_0_4_2_enexo_2
      | reg_act_regs_data_3_4_3_enexo_2 | reg_act_regs_data_3_4_2_enexo_2 | reg_act_regs_data_2_4_2_enexo_2
      | reg_act_regs_data_0_4_1_enexo_2);
  assign Tanh_for_and_55_ssc = ($signed({1'b0, 25'b1000000000000000000000000}) <
      $signed(({nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm})))
      & (~ Tanh_for_4_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1);
  assign Tanh_for_y_and_55_enex5 = Tanh_for_y_and_ssc & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_72
      | reg_act_regs_data_2_3_3_enexo_1 | reg_act_regs_data_0_3_3_enexo_1 | reg_act_regs_data_3_3_enexo
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_72 | reg_act_regs_data_2_3_1_enexo_1
      | reg_act_regs_data_0_3_2_enexo_1 | reg_act_config_inst_counter_enexo_72 |
      reg_act_regs_data_3_3_2_enexo_1 | reg_act_regs_data_0_3_1_enexo_1 | reg_act_regs_data_2_3_2_enexo_1
      | reg_act_regs_data_1_3_3_enexo_1 | reg_act_regs_data_1_3_2_enexo_1 | reg_act_regs_data_3_3_1_enexo_1
      | reg_act_regs_data_1_3_1_enexo_1 | reg_act_regs_data_3_3_3_enexo_1);
  assign Tanh_for_y_and_56_enex5 = Tanh_for_y_and_ssc & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_73
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_73 | reg_act_config_inst_counter_enexo_73
      | reg_act_regs_data_3_3_2_enexo_2 | reg_act_regs_data_2_3_2_enexo_2 | reg_act_regs_data_1_3_3_enexo_2
      | reg_act_regs_data_3_3_enexo_1 | reg_act_regs_data_0_3_2_enexo_2 | reg_act_regs_data_2_3_3_enexo_2
      | reg_act_regs_data_3_3_3_enexo_2 | reg_act_regs_data_1_3_2_enexo_2 | reg_act_regs_data_3_3_1_enexo_2
      | reg_act_regs_data_0_3_1_enexo_2 | reg_act_regs_data_0_3_3_enexo_2 | reg_act_regs_data_1_3_1_enexo_2
      | reg_act_regs_data_2_3_1_enexo_2);
  assign Tanh_for_and_53_ssc = ($signed({1'b0, 25'b1000000000000000000000000}) <
      $signed(({nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm})))
      & (~ Tanh_for_3_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1);
  assign Tanh_for_y_and_57_enex5 = Tanh_for_y_and_ssc & (reg_act_regs_data_0_2_3_enexo_1
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_74 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_74
      | reg_act_config_inst_counter_enexo_74 | reg_act_regs_data_3_2_enexo | reg_act_regs_data_1_2_2_enexo_1
      | reg_act_regs_data_2_2_2_enexo_1 | reg_act_regs_data_0_2_1_enexo_1 | reg_act_regs_data_2_2_1_enexo_1
      | reg_act_regs_data_0_2_2_enexo_1 | reg_act_regs_data_2_2_3_enexo_1 | reg_act_regs_data_3_2_2_enexo_1
      | reg_act_regs_data_1_2_3_enexo_1 | reg_act_regs_data_3_2_1_enexo_1 | reg_act_regs_data_3_2_3_enexo_1
      | reg_act_regs_data_1_2_1_enexo_1);
  assign Tanh_for_y_and_58_enex5 = Tanh_for_y_and_ssc & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_75
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_75 | reg_act_config_inst_counter_enexo_75
      | reg_act_regs_data_3_2_enexo_1 | reg_act_regs_data_3_2_2_enexo_2 | reg_act_regs_data_2_2_2_enexo_2
      | reg_act_regs_data_1_2_1_enexo_2 | reg_act_regs_data_3_2_3_enexo_2 | reg_act_regs_data_2_2_1_enexo_2
      | reg_act_regs_data_0_2_2_enexo_2 | reg_act_regs_data_1_2_3_enexo_2 | reg_act_regs_data_0_2_3_enexo_2
      | reg_act_regs_data_0_2_1_enexo_2 | reg_act_regs_data_2_2_3_enexo_2 | reg_act_regs_data_1_2_2_enexo_2
      | reg_act_regs_data_3_2_1_enexo_2);
  assign Tanh_for_and_51_ssc = ($signed({1'b0, 25'b1000000000000000000000000}) <
      $signed(({nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm})))
      & (~ Tanh_for_2_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1);
  assign Tanh_for_y_and_59_enex5 = Tanh_for_y_and_ssc & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_76
      | reg_act_regs_data_1_1_2_enexo_1 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_76
      | reg_act_regs_data_2_1_enexo | reg_act_regs_data_3_1_2_enexo_1 | reg_act_regs_data_1_1_1_enexo_1
      | reg_act_regs_data_0_1_2_enexo_1 | reg_act_config_inst_counter_enexo_76 |
      reg_act_regs_data_2_1_1_enexo_1 | reg_act_regs_data_0_1_3_enexo_1 | reg_act_regs_data_3_1_1_enexo_1
      | reg_act_regs_data_3_1_3_enexo_1 | reg_act_regs_data_1_1_3_enexo_1 | reg_act_regs_data_0_1_1_enexo_1
      | reg_act_regs_data_2_1_3_enexo_1 | reg_act_regs_data_2_1_2_enexo_1);
  assign Tanh_for_y_and_60_enex5 = Tanh_for_y_and_ssc & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_77
      | reg_act_regs_data_1_1_2_enexo_2 | reg_act_regs_data_2_1_3_enexo_2 | reg_act_regs_data_1_1_3_enexo_2
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_77 | reg_act_regs_data_2_1_2_enexo_2
      | reg_act_regs_data_0_1_1_enexo_2 | reg_act_regs_data_0_1_3_enexo_2 | reg_act_regs_data_3_1_2_enexo_2
      | reg_act_regs_data_2_1_1_enexo_2 | reg_act_regs_data_1_1_1_enexo_2 | reg_act_regs_data_0_1_2_enexo_2
      | reg_act_config_inst_counter_enexo_77 | reg_act_regs_data_2_1_enexo_1 | reg_act_regs_data_3_1_1_enexo_2
      | reg_act_regs_data_3_1_3_enexo_2);
  assign Tanh_for_and_49_ssc = ($signed({1'b0, 25'b1000000000000000000000000}) <
      $signed(({nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm})))
      & (~ Tanh_for_1_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1);
  assign Tanh_for_y_and_61_enex5 = Tanh_for_y_and_ssc & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_78
      | reg_act_regs_data_2_0_2_enexo_1 | reg_act_regs_data_3_0_2_enexo_1 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_78
      | reg_act_regs_data_3_0_enexo | reg_act_regs_data_1_0_1_enexo_1 | reg_act_regs_data_0_0_1_enexo_1
      | reg_act_regs_data_2_0_3_enexo_1 | reg_act_regs_data_3_0_3_enexo_1 | reg_act_regs_data_1_0_2_enexo_1
      | reg_act_regs_data_1_0_3_enexo_1 | reg_act_regs_data_2_0_1_enexo_1 | reg_act_regs_data_3_0_1_enexo_1
      | reg_act_regs_data_0_0_3_enexo_1 | reg_act_config_inst_counter_enexo_78 |
      reg_act_regs_data_0_0_2_enexo_1);
  assign Tanh_for_y_and_62_enex5 = Tanh_for_y_and_ssc & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_79
      | reg_act_regs_data_3_0_1_enexo_2 | reg_act_regs_data_2_0_1_enexo_2 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_79
      | reg_act_regs_data_2_0_3_enexo_2 | reg_act_regs_data_1_0_1_enexo_2 | reg_act_regs_data_3_0_enexo_1
      | reg_act_config_inst_counter_enexo_79 | reg_act_regs_data_1_0_3_enexo_2 |
      reg_act_regs_data_3_0_2_enexo_2 | reg_act_regs_data_1_0_2_enexo_2 | reg_act_regs_data_0_0_1_enexo_2
      | reg_act_regs_data_0_0_3_enexo_2 | reg_act_regs_data_0_0_2_enexo_2 | reg_act_regs_data_2_0_2_enexo_2
      | reg_act_regs_data_3_0_3_enexo_2);
  assign Relu_for_y_qelse_and_ssc = ActUnit_RunInst_switch_lp_and_802_cse & and_dcpl_83
      & (~ (act_config_in_InstFetch_mux_tmp[5])) & and_dcpl_86;
  assign Relu_for_y_qelse_and_31_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_regs_data_1_15_enexo_2
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_80 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_80
      | reg_act_regs_data_2_15_1_enexo_3 | reg_act_regs_data_3_15_1_enexo_3 | reg_act_config_inst_counter_enexo_80
      | reg_act_regs_data_1_15_1_enexo_3 | reg_act_regs_data_0_15_1_enexo_3);
  assign Relu_for_y_qelse_and_32_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_81
      | reg_act_config_inst_counter_enexo_81 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_81
      | reg_act_regs_data_1_15_2_enexo_3 | reg_act_regs_data_1_15_enexo_3 | reg_act_regs_data_3_15_2_enexo_3
      | reg_act_regs_data_0_15_2_enexo_3 | reg_act_regs_data_2_15_2_enexo_3);
  assign Relu_for_y_qelse_and_33_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_82
      | reg_act_regs_data_1_15_enexo_4 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_82
      | reg_act_regs_data_1_15_3_enexo_3 | reg_act_regs_data_3_15_3_enexo_3 | reg_act_regs_data_0_15_3_enexo_3
      | reg_act_config_inst_counter_enexo_82 | reg_act_regs_data_2_15_3_enexo_3);
  assign Relu_for_y_qelse_and_34_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_83
      | reg_act_regs_data_0_14_enexo_2 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_83
      | reg_act_regs_data_3_14_1_enexo_3 | reg_act_regs_data_0_14_1_enexo_3 | reg_act_regs_data_2_14_1_enexo_3
      | reg_act_regs_data_1_14_1_enexo_3 | reg_act_config_inst_counter_enexo_83);
  assign Relu_for_y_qelse_and_35_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_84
      | reg_act_config_inst_counter_enexo_84 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_84
      | reg_act_regs_data_0_14_enexo_3 | reg_act_regs_data_0_14_2_enexo_3 | reg_act_regs_data_1_14_2_enexo_3
      | reg_act_regs_data_2_14_2_enexo_3 | reg_act_regs_data_3_14_2_enexo_3);
  assign Relu_for_y_qelse_and_36_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_regs_data_0_14_3_enexo_3
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_85 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_85
      | reg_act_regs_data_0_14_enexo_4 | reg_act_config_inst_counter_enexo_85 | reg_act_regs_data_1_14_3_enexo_3
      | reg_act_regs_data_2_14_3_enexo_3 | reg_act_regs_data_3_14_3_enexo_3);
  assign Relu_for_y_qelse_and_37_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_config_inst_counter_enexo_86
      | reg_act_regs_data_2_13_1_enexo_3 | reg_act_regs_data_3_13_enexo_2 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_86
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_86 | reg_act_regs_data_0_13_1_enexo_3
      | reg_act_regs_data_3_13_1_enexo_3 | reg_act_regs_data_1_13_1_enexo_3);
  assign Relu_for_y_qelse_and_38_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_87
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_87 | reg_act_regs_data_3_13_enexo_3
      | reg_act_config_inst_counter_enexo_87 | reg_act_regs_data_3_13_2_enexo_3 |
      reg_act_regs_data_0_13_2_enexo_3 | reg_act_regs_data_2_13_2_enexo_3 | reg_act_regs_data_1_13_2_enexo_3);
  assign Relu_for_y_qelse_and_39_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_88
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_88 | reg_act_regs_data_3_13_3_enexo_3
      | reg_act_regs_data_3_13_enexo_4 | reg_act_regs_data_2_13_3_enexo_3 | reg_act_config_inst_counter_enexo_88
      | reg_act_regs_data_0_13_3_enexo_3 | reg_act_regs_data_1_13_3_enexo_3);
  assign Relu_for_y_qelse_and_40_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_89
      | reg_act_config_inst_counter_enexo_89 | reg_act_regs_data_0_12_1_enexo_3 |
      reg_act_regs_data_0_12_enexo_2 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_89
      | reg_act_regs_data_3_12_1_enexo_3 | reg_act_regs_data_2_12_1_enexo_3 | reg_act_regs_data_1_12_1_enexo_3);
  assign Relu_for_y_qelse_and_41_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_90
      | reg_act_regs_data_2_12_2_enexo_3 | reg_act_regs_data_0_12_enexo_3 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_90
      | reg_act_regs_data_0_12_2_enexo_3 | reg_act_regs_data_3_12_2_enexo_3 | reg_act_regs_data_1_12_2_enexo_3
      | reg_act_config_inst_counter_enexo_90);
  assign Relu_for_y_qelse_and_42_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_91
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_91 | reg_act_regs_data_0_12_enexo_4
      | reg_act_regs_data_2_12_3_enexo_3 | reg_act_regs_data_3_12_3_enexo_3 | reg_act_config_inst_counter_enexo_91
      | reg_act_regs_data_0_12_3_enexo_3 | reg_act_regs_data_1_12_3_enexo_3);
  assign Relu_for_y_qelse_and_43_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_regs_data_2_11_enexo_2
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_92 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_92
      | reg_act_config_inst_counter_enexo_92 | reg_act_regs_data_1_11_1_enexo_3 |
      reg_act_regs_data_3_11_1_enexo_3 | reg_act_regs_data_0_11_1_enexo_3 | reg_act_regs_data_2_11_1_enexo_3);
  assign Relu_for_y_qelse_and_44_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_93
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_93 | reg_act_regs_data_2_11_enexo_3
      | reg_act_config_inst_counter_enexo_93 | reg_act_regs_data_2_11_2_enexo_3 |
      reg_act_regs_data_0_11_2_enexo_3 | reg_act_regs_data_3_11_2_enexo_3 | reg_act_regs_data_1_11_2_enexo_3);
  assign Relu_for_y_qelse_and_45_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_regs_data_0_11_3_enexo_3
      | reg_act_regs_data_2_11_enexo_4 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_94
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_94 | reg_act_config_inst_counter_enexo_94
      | reg_act_regs_data_2_11_3_enexo_3 | reg_act_regs_data_1_11_3_enexo_3 | reg_act_regs_data_3_11_3_enexo_3);
  assign Relu_for_y_qelse_and_46_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_config_inst_counter_enexo_95
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_95 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_95
      | reg_act_regs_data_0_10_enexo_2 | reg_act_regs_data_3_10_1_enexo_3 | reg_act_regs_data_1_10_1_enexo_3
      | reg_act_regs_data_2_10_1_enexo_3 | reg_act_regs_data_0_10_1_enexo_3);
  assign Relu_for_y_qelse_and_47_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_96
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_96 | reg_act_regs_data_0_10_enexo_3
      | reg_act_config_inst_counter_enexo_96 | reg_act_regs_data_0_10_2_enexo_3 |
      reg_act_regs_data_2_10_2_enexo_3 | reg_act_regs_data_3_10_2_enexo_3 | reg_act_regs_data_1_10_2_enexo_3);
  assign Relu_for_y_qelse_and_48_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_97
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_97 | reg_act_regs_data_2_10_3_enexo_3
      | reg_act_regs_data_3_10_3_enexo_3 | reg_act_regs_data_0_10_3_enexo_3 | reg_act_regs_data_0_10_enexo_4
      | reg_act_config_inst_counter_enexo_97 | reg_act_regs_data_1_10_3_enexo_3);
  assign Relu_for_y_qelse_and_49_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_98
      | reg_act_regs_data_2_9_1_enexo_3 | reg_act_regs_data_1_9_enexo_2 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_98
      | reg_act_regs_data_1_9_1_enexo_3 | reg_act_regs_data_3_9_1_enexo_3 | reg_act_config_inst_counter_enexo_98
      | reg_act_regs_data_0_9_1_enexo_3);
  assign Relu_for_y_qelse_and_50_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_99
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_99 | reg_act_regs_data_3_9_2_enexo_3
      | reg_act_regs_data_0_9_2_enexo_3 | reg_act_regs_data_1_9_2_enexo_3 | reg_act_regs_data_2_9_2_enexo_3
      | reg_act_regs_data_1_9_enexo_3 | reg_act_config_inst_counter_enexo_99);
  assign Relu_for_y_qelse_and_51_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_100
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_100 | reg_act_regs_data_0_9_3_enexo_3
      | reg_act_regs_data_3_9_3_enexo_3 | reg_act_regs_data_1_9_3_enexo_3 | reg_act_regs_data_1_9_enexo_4
      | reg_act_regs_data_2_9_3_enexo_3 | reg_act_config_inst_counter_enexo_100);
  assign Relu_for_y_qelse_and_52_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_101
      | reg_act_regs_data_2_8_enexo_2 | reg_act_regs_data_1_8_1_enexo_3 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_101
      | reg_act_regs_data_3_8_1_enexo_3 | reg_act_regs_data_0_8_1_enexo_3 | reg_act_config_inst_counter_enexo_101
      | reg_act_regs_data_2_8_1_enexo_3);
  assign Relu_for_y_qelse_and_53_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_102
      | reg_act_regs_data_3_8_2_enexo_3 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_102
      | reg_act_config_inst_counter_enexo_102 | reg_act_regs_data_2_8_enexo_3 | reg_act_regs_data_2_8_2_enexo_3
      | reg_act_regs_data_1_8_2_enexo_3 | reg_act_regs_data_0_8_2_enexo_3);
  assign Relu_for_y_qelse_and_54_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_regs_data_0_8_3_enexo_3
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_103 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_103
      | reg_act_regs_data_2_8_enexo_4 | reg_act_regs_data_3_8_3_enexo_3 | reg_act_regs_data_2_8_3_enexo_3
      | reg_act_regs_data_1_8_3_enexo_3 | reg_act_config_inst_counter_enexo_103);
  assign Relu_for_y_qelse_and_55_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_104
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_104 | reg_act_regs_data_1_7_1_enexo_3
      | reg_act_regs_data_1_7_enexo_2 | reg_act_regs_data_2_7_1_enexo_3 | reg_act_regs_data_3_7_1_enexo_3
      | reg_act_config_inst_counter_enexo_104 | reg_act_regs_data_0_7_1_enexo_3);
  assign Relu_for_y_qelse_and_56_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_105
      | reg_act_regs_data_1_7_enexo_3 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_105
      | reg_act_regs_data_1_7_2_enexo_3 | reg_act_regs_data_3_7_2_enexo_3 | reg_act_config_inst_counter_enexo_105
      | reg_act_regs_data_2_7_2_enexo_3 | reg_act_regs_data_0_7_2_enexo_3);
  assign Relu_for_y_qelse_and_57_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_regs_data_1_7_enexo_4
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_106 | reg_act_regs_data_0_7_3_enexo_3
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_106 | reg_act_regs_data_3_7_3_enexo_3
      | reg_act_regs_data_2_7_3_enexo_3 | reg_act_config_inst_counter_enexo_106 |
      reg_act_regs_data_1_7_3_enexo_3);
  assign Relu_for_y_qelse_and_58_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_regs_data_0_6_1_enexo_3
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_107 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_107
      | reg_act_regs_data_3_6_enexo_2 | reg_act_config_inst_counter_enexo_107 | reg_act_regs_data_2_6_1_enexo_3
      | reg_act_regs_data_1_6_1_enexo_3 | reg_act_regs_data_3_6_1_enexo_3);
  assign Relu_for_y_qelse_and_59_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_108
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_108 | reg_act_regs_data_3_6_enexo_3
      | reg_act_config_inst_counter_enexo_108 | reg_act_regs_data_0_6_2_enexo_3 |
      reg_act_regs_data_3_6_2_enexo_3 | reg_act_regs_data_2_6_2_enexo_3 | reg_act_regs_data_1_6_2_enexo_3);
  assign Relu_for_y_qelse_and_60_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_regs_data_3_6_enexo_4
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_109 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_109
      | reg_act_regs_data_0_6_3_enexo_3 | reg_act_config_inst_counter_enexo_109 |
      reg_act_regs_data_1_6_3_enexo_3 | reg_act_regs_data_3_6_3_enexo_3 | reg_act_regs_data_2_6_3_enexo_3);
  assign Relu_for_y_qelse_and_61_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_110
      | reg_act_config_inst_counter_enexo_110 | reg_act_regs_data_1_5_enexo_2 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_110
      | reg_act_regs_data_3_5_1_enexo_3 | reg_act_regs_data_1_5_1_enexo_3 | reg_act_regs_data_2_5_1_enexo_3
      | reg_act_regs_data_0_5_1_enexo_3);
  assign Relu_for_y_qelse_and_62_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_111
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_111 | reg_act_config_inst_counter_enexo_111
      | reg_act_regs_data_0_5_2_enexo_3 | reg_act_regs_data_3_5_2_enexo_3 | reg_act_regs_data_1_5_enexo_3
      | reg_act_regs_data_1_5_2_enexo_3 | reg_act_regs_data_2_5_2_enexo_3);
  assign Relu_for_y_qelse_and_63_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_112
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_112 | reg_act_regs_data_1_5_enexo_4
      | reg_act_regs_data_0_5_3_enexo_3 | reg_act_regs_data_3_5_3_enexo_3 | reg_act_config_inst_counter_enexo_112
      | reg_act_regs_data_2_5_3_enexo_3 | reg_act_regs_data_1_5_3_enexo_3);
  assign Relu_for_y_qelse_and_64_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_113
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_113 | reg_act_regs_data_3_4_enexo_2
      | reg_act_regs_data_1_4_1_enexo_3 | reg_act_regs_data_3_4_1_enexo_3 | reg_act_regs_data_2_4_1_enexo_3
      | reg_act_config_inst_counter_enexo_113 | reg_act_regs_data_0_4_1_enexo_3);
  assign Relu_for_y_qelse_and_65_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_regs_data_3_4_enexo_3
      | reg_act_regs_data_2_4_2_enexo_3 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_114
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_114 | reg_act_regs_data_3_4_2_enexo_3
      | reg_act_config_inst_counter_enexo_114 | reg_act_regs_data_1_4_2_enexo_3 |
      reg_act_regs_data_0_4_2_enexo_3);
  assign Relu_for_y_qelse_and_66_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_regs_data_0_4_3_enexo_3
      | reg_act_regs_data_3_4_enexo_4 | reg_act_config_inst_counter_enexo_115 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_115
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_115 | reg_act_regs_data_3_4_3_enexo_3
      | reg_act_regs_data_2_4_3_enexo_3 | reg_act_regs_data_1_4_3_enexo_3);
  assign Relu_for_y_qelse_and_67_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_116
      | reg_act_config_inst_counter_enexo_116 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_116
      | reg_act_regs_data_3_3_enexo_2 | reg_act_regs_data_0_3_1_enexo_3 | reg_act_regs_data_3_3_1_enexo_3
      | reg_act_regs_data_2_3_1_enexo_3 | reg_act_regs_data_1_3_1_enexo_3);
  assign Relu_for_y_qelse_and_68_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_regs_data_3_3_enexo_3
      | reg_act_regs_data_2_3_2_enexo_3 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_117
      | reg_act_regs_data_3_3_2_enexo_3 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_117
      | reg_act_regs_data_0_3_2_enexo_3 | reg_act_config_inst_counter_enexo_117 |
      reg_act_regs_data_1_3_2_enexo_3);
  assign Relu_for_y_qelse_and_69_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_118
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_118 | reg_act_regs_data_3_3_enexo_4
      | reg_act_config_inst_counter_enexo_118 | reg_act_regs_data_1_3_3_enexo_3 |
      reg_act_regs_data_0_3_3_enexo_3 | reg_act_regs_data_3_3_3_enexo_3 | reg_act_regs_data_2_3_3_enexo_3);
  assign Relu_for_y_qelse_and_70_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_119
      | reg_act_regs_data_3_2_enexo_2 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_119
      | reg_act_regs_data_3_2_1_enexo_3 | reg_act_regs_data_1_2_1_enexo_3 | reg_act_regs_data_2_2_1_enexo_3
      | reg_act_config_inst_counter_enexo_119 | reg_act_regs_data_0_2_1_enexo_3);
  assign Relu_for_y_qelse_and_71_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_120
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_120 | reg_act_regs_data_0_2_2_enexo_3
      | reg_act_regs_data_2_2_2_enexo_3 | reg_act_regs_data_3_2_enexo_3 | reg_act_regs_data_1_2_2_enexo_3
      | reg_act_regs_data_3_2_2_enexo_3 | reg_act_config_inst_counter_enexo_120);
  assign Relu_for_y_qelse_and_72_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_121
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_121 | reg_act_regs_data_0_2_3_enexo_3
      | reg_act_regs_data_2_2_3_enexo_3 | reg_act_regs_data_3_2_enexo_4 | reg_act_regs_data_3_2_3_enexo_3
      | reg_act_config_inst_counter_enexo_121 | reg_act_regs_data_1_2_3_enexo_3);
  assign Relu_for_y_qelse_and_73_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_122
      | reg_act_regs_data_2_1_enexo_2 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_122
      | reg_act_regs_data_0_1_1_enexo_3 | reg_act_regs_data_1_1_1_enexo_3 | reg_act_regs_data_3_1_1_enexo_3
      | reg_act_regs_data_2_1_1_enexo_3 | reg_act_config_inst_counter_enexo_122);
  assign Relu_for_y_qelse_and_74_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_123
      | reg_act_regs_data_0_1_2_enexo_3 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_123
      | reg_act_regs_data_3_1_2_enexo_3 | reg_act_regs_data_2_1_2_enexo_3 | reg_act_regs_data_2_1_enexo_3
      | reg_act_config_inst_counter_enexo_123 | reg_act_regs_data_1_1_2_enexo_3);
  assign Relu_for_y_qelse_and_75_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_124
      | reg_act_config_inst_counter_enexo_124 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_124
      | reg_act_regs_data_1_1_3_enexo_3 | reg_act_regs_data_0_1_3_enexo_3 | reg_act_regs_data_2_1_3_enexo_3
      | reg_act_regs_data_3_1_3_enexo_3 | reg_act_regs_data_2_1_enexo_4);
  assign Relu_for_y_qelse_and_76_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_125
      | reg_act_regs_data_1_0_1_enexo_3 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_125
      | reg_act_regs_data_0_0_1_enexo_3 | reg_act_config_inst_counter_enexo_125 |
      reg_act_regs_data_2_0_1_enexo_3 | reg_act_regs_data_3_0_enexo_2 | reg_act_regs_data_3_0_1_enexo_3);
  assign Relu_for_y_qelse_and_77_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_126
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_126 | reg_act_regs_data_0_0_2_enexo_3
      | reg_act_regs_data_3_0_2_enexo_3 | reg_act_regs_data_3_0_enexo_3 | reg_act_regs_data_2_0_2_enexo_3
      | reg_act_regs_data_1_0_2_enexo_3 | reg_act_config_inst_counter_enexo_126);
  assign Relu_for_y_qelse_and_78_enex5 = Relu_for_y_qelse_and_ssc & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_127
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_127 | reg_act_regs_data_2_0_3_enexo_3
      | reg_act_config_inst_counter_enexo_127 | reg_act_regs_data_3_0_3_enexo_3 |
      reg_act_regs_data_3_0_enexo_4 | reg_act_regs_data_0_0_3_enexo_3 | reg_act_regs_data_1_0_3_enexo_3);
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_and_cse = ActUnitRun_wen & (~ and_dcpl_1228);
  assign operator_32_8_true_AC_TRN_AC_WRAP_2_and_16_cse = ActUnit_RunInst_switch_lp_and_802_cse
      & and_dcpl_83 & (act_config_in_InstFetch_mux_tmp[6:5]==2'b11);
  assign ActUnit_RunInst_curr_inst_and_enex5 = ActUnit_RunInst_switch_lp_and_802_cse
      & is_start_sva & (reg_act_config_inst_counter_enexo_128 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_128
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_128);
  assign operator_32_8_true_AC_TRN_AC_WRAP_and_cse = ActUnit_RunInst_switch_lp_and_802_cse
      & and_dcpl_117;
  assign operator_32_8_true_AC_TRN_AC_WRAP_and_23_cse = operator_32_8_true_AC_TRN_AC_WRAP_2_and_cse
      & and_dcpl_117;
  assign ActUnit_RunInst_switch_lp_and_811_cse = ActUnitRun_wen & (~ and_dcpl_849);
  assign ActUnit_RunInst_switch_lp_and_813_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_129 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_129
      | reg_act_regs_data_3_0_2_enexo_4 | reg_act_config_inst_counter_enexo_129 |
      reg_act_regs_data_0_0_2_enexo_4 | reg_act_regs_data_1_0_2_enexo_4 | reg_act_regs_data_2_0_2_enexo_4);
  assign ActUnit_RunInst_switch_lp_and_814_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_130 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_130
      | reg_act_config_inst_counter_enexo_130 | reg_act_regs_data_1_0_3_enexo_4 |
      reg_act_regs_data_3_0_3_enexo_4 | reg_act_regs_data_2_0_3_enexo_4 | reg_act_regs_data_0_0_3_enexo_4);
  assign ActUnit_RunInst_switch_lp_and_815_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_131 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_131
      | reg_act_regs_data_2_0_1_enexo_4 | reg_act_regs_data_1_0_1_enexo_4 | reg_act_regs_data_0_0_1_enexo_4
      | reg_act_config_inst_counter_enexo_131 | reg_act_regs_data_3_0_1_enexo_4);
  assign nv_scvector_cctor_nv_scvector_6_for_and_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_132 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_132
      | reg_act_config_inst_counter_enexo_132 | reg_act_regs_data_1_1_2_enexo_4 |
      reg_act_regs_data_3_1_2_enexo_4 | reg_act_regs_data_0_1_2_enexo_4 | reg_act_regs_data_2_1_2_enexo_4);
  assign nv_scvector_cctor_nv_scvector_6_for_and_15_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_regs_data_1_1_3_enexo_4 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_133
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_133 | reg_act_config_inst_counter_enexo_133
      | reg_act_regs_data_0_1_3_enexo_4 | reg_act_regs_data_2_1_3_enexo_4 | reg_act_regs_data_3_1_3_enexo_4);
  assign nv_scvector_cctor_nv_scvector_6_for_and_16_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_134 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_134
      | reg_act_regs_data_3_1_1_enexo_4 | reg_act_regs_data_2_1_1_enexo_4 | reg_act_regs_data_1_1_1_enexo_4
      | reg_act_regs_data_0_1_1_enexo_4 | reg_act_config_inst_counter_enexo_134);
  assign nv_scvector_cctor_nv_scvector_6_for_and_17_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_135 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_135
      | reg_act_regs_data_0_2_2_enexo_4 | reg_act_config_inst_counter_enexo_135 |
      reg_act_regs_data_1_2_2_enexo_4 | reg_act_regs_data_2_2_2_enexo_4 | reg_act_regs_data_3_2_2_enexo_4);
  assign nv_scvector_cctor_nv_scvector_6_for_and_18_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_136 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_136
      | reg_act_config_inst_counter_enexo_136 | reg_act_regs_data_1_2_3_enexo_4 |
      reg_act_regs_data_2_2_3_enexo_4 | reg_act_regs_data_3_2_3_enexo_4 | reg_act_regs_data_0_2_3_enexo_4);
  assign nv_scvector_cctor_nv_scvector_6_for_and_19_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_137 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_137
      | reg_act_regs_data_1_2_1_enexo_4 | reg_act_regs_data_3_2_1_enexo_4 | reg_act_config_inst_counter_enexo_137
      | reg_act_regs_data_0_2_1_enexo_4 | reg_act_regs_data_2_2_1_enexo_4);
  assign nv_scvector_cctor_nv_scvector_6_for_and_20_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_138 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_138
      | reg_act_regs_data_1_3_2_enexo_4 | reg_act_regs_data_0_3_2_enexo_4 | reg_act_config_inst_counter_enexo_138
      | reg_act_regs_data_2_3_2_enexo_4 | reg_act_regs_data_3_3_2_enexo_4);
  assign nv_scvector_cctor_nv_scvector_6_for_and_21_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_139 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_139
      | reg_act_regs_data_0_3_3_enexo_4 | reg_act_config_inst_counter_enexo_139 |
      reg_act_regs_data_2_3_3_enexo_4 | reg_act_regs_data_1_3_3_enexo_4 | reg_act_regs_data_3_3_3_enexo_4);
  assign nv_scvector_cctor_nv_scvector_6_for_and_22_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_140 | reg_act_regs_data_0_3_1_enexo_4
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_140 | reg_act_config_inst_counter_enexo_140
      | reg_act_regs_data_3_3_1_enexo_4 | reg_act_regs_data_2_3_1_enexo_4 | reg_act_regs_data_1_3_1_enexo_4);
  assign nv_scvector_cctor_nv_scvector_6_for_and_23_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_regs_data_3_4_2_enexo_4 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_141
      | reg_act_regs_data_2_4_2_enexo_4 | reg_act_config_inst_counter_enexo_141 |
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_141 | reg_act_regs_data_1_4_2_enexo_4
      | reg_act_regs_data_0_4_2_enexo_4);
  assign nv_scvector_cctor_nv_scvector_6_for_and_24_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_regs_data_3_4_3_enexo_4 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_142
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_142 | reg_act_regs_data_2_4_3_enexo_4
      | reg_act_regs_data_1_4_3_enexo_4 | reg_act_config_inst_counter_enexo_142 |
      reg_act_regs_data_0_4_3_enexo_4);
  assign nv_scvector_cctor_nv_scvector_6_for_and_25_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_143 | reg_act_regs_data_2_4_1_enexo_4
      | reg_act_regs_data_0_4_1_enexo_4 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_143
      | reg_act_regs_data_1_4_1_enexo_4 | reg_act_config_inst_counter_enexo_143 |
      reg_act_regs_data_3_4_1_enexo_4);
  assign nv_scvector_cctor_nv_scvector_6_for_and_26_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_144 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_144
      | reg_act_regs_data_1_5_2_enexo_4 | reg_act_regs_data_2_5_2_enexo_4 | reg_act_config_inst_counter_enexo_144
      | reg_act_regs_data_3_5_2_enexo_4 | reg_act_regs_data_0_5_2_enexo_4);
  assign nv_scvector_cctor_nv_scvector_6_for_and_27_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_145 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_145
      | reg_act_regs_data_0_5_3_enexo_4 | reg_act_regs_data_1_5_3_enexo_4 | reg_act_regs_data_3_5_3_enexo_4
      | reg_act_regs_data_2_5_3_enexo_4 | reg_act_config_inst_counter_enexo_145);
  assign nv_scvector_cctor_nv_scvector_6_for_and_28_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_regs_data_2_5_1_enexo_4 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_146
      | reg_act_regs_data_3_5_1_enexo_4 | reg_act_config_inst_counter_enexo_146 |
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_146 | reg_act_regs_data_0_5_1_enexo_4
      | reg_act_regs_data_1_5_1_enexo_4);
  assign nv_scvector_cctor_nv_scvector_6_for_and_29_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_147 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_147
      | reg_act_config_inst_counter_enexo_147 | reg_act_regs_data_2_6_2_enexo_4 |
      reg_act_regs_data_1_6_2_enexo_4 | reg_act_regs_data_3_6_2_enexo_4 | reg_act_regs_data_0_6_2_enexo_4);
  assign nv_scvector_cctor_nv_scvector_6_for_and_30_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_148 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_148
      | reg_act_regs_data_1_6_3_enexo_4 | reg_act_config_inst_counter_enexo_148 |
      reg_act_regs_data_2_6_3_enexo_4 | reg_act_regs_data_3_6_3_enexo_4 | reg_act_regs_data_0_6_3_enexo_4);
  assign nv_scvector_cctor_nv_scvector_6_for_and_31_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_149 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_149
      | reg_act_config_inst_counter_enexo_149 | reg_act_regs_data_0_6_1_enexo_4 |
      reg_act_regs_data_2_6_1_enexo_4 | reg_act_regs_data_1_6_1_enexo_4 | reg_act_regs_data_3_6_1_enexo_4);
  assign nv_scvector_cctor_nv_scvector_6_for_and_32_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_150 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_150
      | reg_act_regs_data_3_7_2_enexo_4 | reg_act_regs_data_1_7_2_enexo_4 | reg_act_regs_data_0_7_2_enexo_4
      | reg_act_regs_data_2_7_2_enexo_4 | reg_act_config_inst_counter_enexo_150);
  assign nv_scvector_cctor_nv_scvector_6_for_and_33_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_151 | reg_act_regs_data_1_7_3_enexo_4
      | reg_act_regs_data_2_7_3_enexo_4 | reg_act_regs_data_0_7_3_enexo_4 | reg_act_config_inst_counter_enexo_151
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_151 | reg_act_regs_data_3_7_3_enexo_4);
  assign nv_scvector_cctor_nv_scvector_6_for_and_34_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_152 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_152
      | reg_act_regs_data_0_7_1_enexo_4 | reg_act_config_inst_counter_enexo_152 |
      reg_act_regs_data_3_7_1_enexo_4 | reg_act_regs_data_2_7_1_enexo_4 | reg_act_regs_data_1_7_1_enexo_4);
  assign nv_scvector_cctor_nv_scvector_6_for_and_35_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_153 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_153
      | reg_act_regs_data_2_8_2_enexo_4 | reg_act_regs_data_1_8_2_enexo_4 | reg_act_config_inst_counter_enexo_153
      | reg_act_regs_data_0_8_2_enexo_4 | reg_act_regs_data_3_8_2_enexo_4);
  assign nv_scvector_cctor_nv_scvector_6_for_and_36_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_154 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_154
      | reg_act_regs_data_3_8_3_enexo_4 | reg_act_regs_data_1_8_3_enexo_4 | reg_act_regs_data_0_8_3_enexo_4
      | reg_act_config_inst_counter_enexo_154 | reg_act_regs_data_2_8_3_enexo_4);
  assign nv_scvector_cctor_nv_scvector_6_for_and_37_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_155 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_155
      | reg_act_regs_data_3_8_1_enexo_4 | reg_act_regs_data_1_8_1_enexo_4 | reg_act_regs_data_2_8_1_enexo_4
      | reg_act_config_inst_counter_enexo_155 | reg_act_regs_data_0_8_1_enexo_4);
  assign nv_scvector_cctor_nv_scvector_6_for_and_38_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_156 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_156
      | reg_act_config_inst_counter_enexo_156 | reg_act_regs_data_3_9_2_enexo_4 |
      reg_act_regs_data_2_9_2_enexo_4 | reg_act_regs_data_0_9_2_enexo_4 | reg_act_regs_data_1_9_2_enexo_4);
  assign nv_scvector_cctor_nv_scvector_6_for_and_39_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_157 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_157
      | reg_act_regs_data_0_9_3_enexo_4 | reg_act_regs_data_1_9_3_enexo_4 | reg_act_regs_data_3_9_3_enexo_4
      | reg_act_regs_data_2_9_3_enexo_4 | reg_act_config_inst_counter_enexo_157);
  assign nv_scvector_cctor_nv_scvector_6_for_and_40_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_158 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_158
      | reg_act_regs_data_1_9_1_enexo_4 | reg_act_regs_data_3_9_1_enexo_4 | reg_act_regs_data_0_9_1_enexo_4
      | reg_act_regs_data_2_9_1_enexo_4 | reg_act_config_inst_counter_enexo_158);
  assign nv_scvector_cctor_nv_scvector_6_for_and_41_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_159 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_159
      | reg_act_regs_data_3_10_2_enexo_4 | reg_act_regs_data_0_10_2_enexo_4 | reg_act_regs_data_2_10_2_enexo_4
      | reg_act_config_inst_counter_enexo_159 | reg_act_regs_data_1_10_2_enexo_4);
  assign nv_scvector_cctor_nv_scvector_6_for_and_42_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_160 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_160
      | reg_act_config_inst_counter_enexo_160 | reg_act_regs_data_2_10_3_enexo_4
      | reg_act_regs_data_0_10_3_enexo_4 | reg_act_regs_data_3_10_3_enexo_4 | reg_act_regs_data_1_10_3_enexo_4);
  assign nv_scvector_cctor_nv_scvector_6_for_and_43_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_161 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_161
      | reg_act_regs_data_0_10_1_enexo_4 | reg_act_config_inst_counter_enexo_161
      | reg_act_regs_data_1_10_1_enexo_4 | reg_act_regs_data_3_10_1_enexo_4 | reg_act_regs_data_2_10_1_enexo_4);
  assign nv_scvector_cctor_nv_scvector_6_for_and_44_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_162 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_162
      | reg_act_config_inst_counter_enexo_162 | reg_act_regs_data_0_11_2_enexo_4
      | reg_act_regs_data_2_11_2_enexo_4 | reg_act_regs_data_3_11_2_enexo_4 | reg_act_regs_data_1_11_2_enexo_4);
  assign nv_scvector_cctor_nv_scvector_6_for_and_45_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_163 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_163
      | reg_act_regs_data_1_11_3_enexo_4 | reg_act_regs_data_3_11_3_enexo_4 | reg_act_regs_data_0_11_3_enexo_4
      | reg_act_regs_data_2_11_3_enexo_4 | reg_act_config_inst_counter_enexo_163);
  assign nv_scvector_cctor_nv_scvector_6_for_and_46_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_164 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_164
      | reg_act_regs_data_2_11_1_enexo_4 | reg_act_regs_data_1_11_1_enexo_4 | reg_act_config_inst_counter_enexo_164
      | reg_act_regs_data_3_11_1_enexo_4 | reg_act_regs_data_0_11_1_enexo_4);
  assign nv_scvector_cctor_nv_scvector_6_for_and_47_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_165 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_165
      | reg_act_regs_data_0_12_2_enexo_4 | reg_act_config_inst_counter_enexo_165
      | reg_act_regs_data_1_12_2_enexo_4 | reg_act_regs_data_3_12_2_enexo_4 | reg_act_regs_data_2_12_2_enexo_4);
  assign nv_scvector_cctor_nv_scvector_6_for_and_48_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_166 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_166
      | reg_act_config_inst_counter_enexo_166 | reg_act_regs_data_3_12_3_enexo_4
      | reg_act_regs_data_2_12_3_enexo_4 | reg_act_regs_data_1_12_3_enexo_4 | reg_act_regs_data_0_12_3_enexo_4);
  assign nv_scvector_cctor_nv_scvector_6_for_and_49_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_167 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_167
      | reg_act_regs_data_3_12_1_enexo_4 | reg_act_config_inst_counter_enexo_167
      | reg_act_regs_data_2_12_1_enexo_4 | reg_act_regs_data_0_12_1_enexo_4 | reg_act_regs_data_1_12_1_enexo_4);
  assign nv_scvector_cctor_nv_scvector_6_for_and_50_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_168 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_168
      | reg_act_regs_data_3_13_2_enexo_4 | reg_act_regs_data_1_13_2_enexo_4 | reg_act_config_inst_counter_enexo_168
      | reg_act_regs_data_0_13_2_enexo_4 | reg_act_regs_data_2_13_2_enexo_4);
  assign nv_scvector_cctor_nv_scvector_6_for_and_51_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_169 | reg_act_regs_data_2_13_3_enexo_4
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_169 | reg_act_regs_data_0_13_3_enexo_4
      | reg_act_regs_data_3_13_3_enexo_4 | reg_act_regs_data_1_13_3_enexo_4 | reg_act_config_inst_counter_enexo_169);
  assign nv_scvector_cctor_nv_scvector_6_for_and_52_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_170 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_170
      | reg_act_regs_data_0_13_1_enexo_4 | reg_act_regs_data_1_13_1_enexo_4 | reg_act_config_inst_counter_enexo_170
      | reg_act_regs_data_2_13_1_enexo_4 | reg_act_regs_data_3_13_1_enexo_4);
  assign nv_scvector_cctor_nv_scvector_6_for_and_53_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_171 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_171
      | reg_act_regs_data_0_14_2_enexo_4 | reg_act_regs_data_3_14_2_enexo_4 | reg_act_regs_data_2_14_2_enexo_4
      | reg_act_config_inst_counter_enexo_171 | reg_act_regs_data_1_14_2_enexo_4);
  assign nv_scvector_cctor_nv_scvector_6_for_and_54_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_172 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_172
      | reg_act_config_inst_counter_enexo_172 | reg_act_regs_data_3_14_3_enexo_4
      | reg_act_regs_data_2_14_3_enexo_4 | reg_act_regs_data_0_14_3_enexo_4 | reg_act_regs_data_1_14_3_enexo_4);
  assign nv_scvector_cctor_nv_scvector_6_for_and_55_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_173 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_173
      | reg_act_regs_data_3_14_1_enexo_4 | reg_act_regs_data_0_14_1_enexo_4 | reg_act_regs_data_2_14_1_enexo_4
      | reg_act_regs_data_1_14_1_enexo_4 | reg_act_config_inst_counter_enexo_173);
  assign nv_scvector_cctor_nv_scvector_6_for_and_56_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_174 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_174
      | reg_act_config_inst_counter_enexo_174 | reg_act_regs_data_1_15_2_enexo_4
      | reg_act_regs_data_3_15_2_enexo_4 | reg_act_regs_data_2_15_2_enexo_4 | reg_act_regs_data_0_15_2_enexo_4);
  assign nv_scvector_cctor_nv_scvector_6_for_and_57_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_175 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_175
      | reg_act_regs_data_3_15_3_enexo_4 | reg_act_regs_data_2_15_3_enexo_4 | reg_act_regs_data_1_15_3_enexo_4
      | reg_act_config_inst_counter_enexo_175 | reg_act_regs_data_0_15_3_enexo_4);
  assign nv_scvector_cctor_nv_scvector_6_for_and_58_enex5 = ActUnit_RunInst_switch_lp_and_811_cse
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_176 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_176
      | reg_act_regs_data_0_15_1_enexo_4 | reg_act_regs_data_3_15_1_enexo_4 | reg_act_regs_data_2_15_1_enexo_4
      | reg_act_regs_data_1_15_1_enexo_4 | reg_act_config_inst_counter_enexo_176);
  assign Gelu_for_if_and_cse = ActUnit_RunInst_switch_lp_and_802_cse & and_dcpl_84
      & and_dcpl_78;
  assign or_243_cse = (~ is_start_sva) | (act_config_in_InstFetch_mux_tmp[7:4]!=4'b0010)
      | (z_out[4]);
  assign ActUnit_RunInst_case_2_for_and_27_seb = and_2350_cse & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign act_write_data_data_and_15_cse = ActUnitRun_wen & (~ and_dcpl_1112);
  assign act_write_data_data_and_ssc = ActUnitRun_wen & ((~ or_dcpl_817) | and_dcpl_1240);
  assign act_write_data_data_and_16_ssc = act_write_data_data_and_ssc & (~ and_dcpl_1112);
  assign act_write_data_data_act_write_data_data_and_26_cse = ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_31
      & (~ and_dcpl_847);
  assign act_write_data_data_and_96_cse = (~ and_dcpl_1112) & and_dcpl_1240;
  assign or_3396_cse = (fsm_output!=4'b0100);
  assign nor_1479_cse = ~((~ (fsm_output[0])) | (fsm_output[3]) | (fsm_output[2]));
  assign nand_cse = ~((ActUnit_PushOutput_if_for_i_4_0_sva_3_0==4'b1110));
  assign mux_665_nl = MUX_s_1_2_2(or_3396_cse, nor_1479_cse, nand_cse);
  assign and_1821_cse = mux_665_nl & ActUnitRun_wen;
  assign nor_1484_cse = ~((fsm_output!=4'b0100));
  assign mux_668_nl = MUX_s_1_2_2(or_tmp_653, nor_1484_cse, ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]);
  assign or_1678_nl = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3:1]!=3'b000);
  assign mux_669_nl = MUX_s_1_2_2(mux_668_nl, or_tmp_653, or_1678_nl);
  assign and_1824_cse = (~ mux_669_nl) & ActUnitRun_wen;
  assign mux_674_nl = MUX_s_1_2_2(or_tmp_653, nor_1484_cse, ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]);
  assign or_1690_nl = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3:1]!=3'b110);
  assign mux_675_nl = MUX_s_1_2_2(mux_674_nl, or_tmp_653, or_1690_nl);
  assign and_1827_cse = (~ mux_675_nl) & ActUnitRun_wen;
  assign or_1702_cse = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0!=4'b0010);
  assign mux_680_nl = MUX_s_1_2_2(or_3396_cse, nor_1479_cse, or_1702_cse);
  assign and_1830_cse = mux_680_nl & ActUnitRun_wen;
  assign or_1714_cse = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0!=4'b1100);
  assign mux_683_nl = MUX_s_1_2_2(or_3396_cse, nor_1479_cse, or_1714_cse);
  assign and_1833_cse = mux_683_nl & ActUnitRun_wen;
  assign and_2344_cse = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1:0]==2'b11);
  assign or_1726_cse = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3:2]!=2'b00);
  assign mux_1529_nl = MUX_s_1_2_2(or_tmp_653, nor_1484_cse, and_2344_cse);
  assign mux_687_nl = MUX_s_1_2_2(mux_1529_nl, or_tmp_653, or_1726_cse);
  assign and_1836_cse = (~ mux_687_nl) & ActUnitRun_wen;
  assign or_1738_cse = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3:2]!=2'b10);
  assign mux_686_nl = MUX_s_1_2_2(or_tmp_653, nor_1484_cse, and_2344_cse);
  assign mux_693_nl = MUX_s_1_2_2(mux_686_nl, or_tmp_653, or_1738_cse);
  assign and_1839_cse = (~ mux_693_nl) & ActUnitRun_wen;
  assign or_1750_cse = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0!=4'b0100);
  assign mux_698_nl = MUX_s_1_2_2(or_3396_cse, nor_1479_cse, or_1750_cse);
  assign and_1842_cse = mux_698_nl & ActUnitRun_wen;
  assign or_1762_cse = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0!=4'b1010);
  assign mux_701_nl = MUX_s_1_2_2(or_3396_cse, nor_1479_cse, or_1762_cse);
  assign and_1845_cse = mux_701_nl & ActUnitRun_wen;
  assign mux_704_nl = MUX_s_1_2_2(or_tmp_653, nor_1484_cse, ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]);
  assign or_1774_nl = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3:1]!=3'b010);
  assign mux_705_nl = MUX_s_1_2_2(mux_704_nl, or_tmp_653, or_1774_nl);
  assign and_1848_cse = (~ mux_705_nl) & ActUnitRun_wen;
  assign mux_710_nl = MUX_s_1_2_2(or_tmp_653, nor_1484_cse, ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]);
  assign or_1786_nl = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3:1]!=3'b100);
  assign mux_711_nl = MUX_s_1_2_2(mux_710_nl, or_tmp_653, or_1786_nl);
  assign and_1851_cse = (~ mux_711_nl) & ActUnitRun_wen;
  assign or_1798_cse = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0!=4'b0110);
  assign mux_716_nl = MUX_s_1_2_2(or_3396_cse, nor_1479_cse, or_1798_cse);
  assign and_1854_cse = mux_716_nl & ActUnitRun_wen;
  assign or_1810_cse = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0!=4'b1000);
  assign mux_719_nl = MUX_s_1_2_2(or_3396_cse, nor_1479_cse, or_1810_cse);
  assign and_1857_cse = mux_719_nl & ActUnitRun_wen;
  assign and_2350_cse = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2:0]==3'b111);
  assign mux_722_nl = MUX_s_1_2_2(or_tmp_653, nor_1484_cse, and_2350_cse);
  assign mux_723_nl = MUX_s_1_2_2(mux_722_nl, or_tmp_653, ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign and_1860_cse = (~ mux_723_nl) & ActUnitRun_wen;
  assign act_mem_banks_read_for_and_cse = ActUnitRun_wen & not_tmp_237;
  assign rva_out_reg_data_and_62_cse = ActUnitRun_wen & (~ not_tmp_495) & or_tmp_146;
  assign while_and_282_cse = (~ and_dcpl_1257) & while_asn_2039;
  assign while_and_283_cse = and_dcpl_1257 & while_asn_2039;
  assign act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_20_itm
      = MUX_v_6_2_2(6'b000000, (act_config_inst_regs_19_sva_dfm_6[5:0]), act_config_ActConfigRead_else_else_not_21);
  assign act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_21_itm
      = MUX_v_8_2_2(8'b00000000, act_config_inst_regs_20_sva_dfm_6, act_config_ActConfigRead_else_else_not_21);
  assign act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_23_itm
      = MUX_v_8_2_2(8'b00000000, act_config_inst_regs_24_sva_dfm_6, act_config_ActConfigRead_else_else_not_21);
  assign mux_433_nl = MUX_s_1_2_2((~ (fsm_output[2])), or_tmp_485, fsm_output[3]);
  assign act_config_output_counter_and_1_cse = ActUnitRun_wen & mux_433_nl;
  assign nl_Silu_for_1_else_else_else_if_acc_nl = conv_u2u_25_26({reg_ActUnit_RunInst_case_14_nv_scvector_cctor_data_0_1_ftd_rsp_0
      , reg_ActUnit_RunInst_case_14_nv_scvector_cctor_data_0_1_ftd_rsp_1 , (reg_ActUnit_RunInst_case_14_nv_scvector_cctor_data_0_1_ftd_1[21:1])})
      + ({reg_ActUnit_RunInst_case_14_nv_scvector_cctor_data_0_1_ftd_rsp_0 , reg_ActUnit_RunInst_case_14_nv_scvector_cctor_data_0_1_ftd_rsp_1
      , reg_ActUnit_RunInst_case_14_nv_scvector_cctor_data_0_1_ftd_1});
  assign Silu_for_1_else_else_else_if_acc_nl = nl_Silu_for_1_else_else_else_if_acc_nl[25:0];
  assign Silu_for_1_else_else_else_if_acc_itm_25_1_1 = readslicef_26_25_1(Silu_for_1_else_else_else_if_acc_nl);
  assign and_1751_cse = and_dcpl_1236 & (~ or_dcpl_1015);
  assign or_1831_cse = (fsm_output[3:1]!=3'b100);
  assign nl_Silu_for_2_else_else_else_if_acc_nl = conv_u2u_25_26({reg_nv_scvector_cctor_nv_scvector_5_for_2_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_2_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , (reg_nv_scvector_cctor_nv_scvector_5_for_2_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:1])})
      + ({reg_nv_scvector_cctor_nv_scvector_5_for_2_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_2_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_5_for_2_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1});
  assign Silu_for_2_else_else_else_if_acc_nl = nl_Silu_for_2_else_else_else_if_acc_nl[25:0];
  assign Silu_for_2_else_else_else_if_acc_itm_25_1_1 = readslicef_26_25_1(Silu_for_2_else_else_else_if_acc_nl);
  assign and_2354_cse = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0==4'b1110);
  assign nl_Silu_for_3_else_else_else_if_acc_nl = conv_u2u_25_26({reg_nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , (reg_nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:1])})
      + ({reg_nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1});
  assign Silu_for_3_else_else_else_if_acc_nl = nl_Silu_for_3_else_else_else_if_acc_nl[25:0];
  assign Silu_for_3_else_else_else_if_acc_itm_25_1_1 = readslicef_26_25_1(Silu_for_3_else_else_else_if_acc_nl);
  assign nl_Silu_for_4_else_else_else_if_acc_nl = conv_u2u_25_26({reg_nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , (reg_nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:1])})
      + ({reg_nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1});
  assign Silu_for_4_else_else_else_if_acc_nl = nl_Silu_for_4_else_else_else_if_acc_nl[25:0];
  assign Silu_for_4_else_else_else_if_acc_itm_25_1_1 = readslicef_26_25_1(Silu_for_4_else_else_else_if_acc_nl);
  assign nand_533_cse = ~((ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1:0]==2'b11));
  assign nl_Silu_for_5_else_else_else_if_acc_nl = conv_u2u_25_26({reg_nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , (reg_nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:1])})
      + ({reg_nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1});
  assign Silu_for_5_else_else_else_if_acc_nl = nl_Silu_for_5_else_else_else_if_acc_nl[25:0];
  assign Silu_for_5_else_else_else_if_acc_itm_25_1_1 = readslicef_26_25_1(Silu_for_5_else_else_else_if_acc_nl);
  assign nl_Silu_for_6_else_else_else_if_acc_nl = conv_u2u_25_26({reg_nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , (reg_nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:1])})
      + ({reg_nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1});
  assign Silu_for_6_else_else_else_if_acc_nl = nl_Silu_for_6_else_else_else_if_acc_nl[25:0];
  assign Silu_for_6_else_else_else_if_acc_itm_25_1_1 = readslicef_26_25_1(Silu_for_6_else_else_else_if_acc_nl);
  assign nl_Silu_for_7_else_else_else_if_acc_nl = conv_u2u_25_26({reg_nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , (reg_nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:1])})
      + ({reg_nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1});
  assign Silu_for_7_else_else_else_if_acc_nl = nl_Silu_for_7_else_else_else_if_acc_nl[25:0];
  assign Silu_for_7_else_else_else_if_acc_itm_25_1_1 = readslicef_26_25_1(Silu_for_7_else_else_else_if_acc_nl);
  assign nl_Silu_for_8_else_else_else_if_acc_nl = conv_u2u_25_26({reg_nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , (reg_nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:1])})
      + ({reg_nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1});
  assign Silu_for_8_else_else_else_if_acc_nl = nl_Silu_for_8_else_else_else_if_acc_nl[25:0];
  assign Silu_for_8_else_else_else_if_acc_itm_25_1_1 = readslicef_26_25_1(Silu_for_8_else_else_else_if_acc_nl);
  assign nl_Silu_for_9_else_else_else_if_acc_nl = conv_u2u_25_26({reg_nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , (reg_nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:1])})
      + ({reg_nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1});
  assign Silu_for_9_else_else_else_if_acc_nl = nl_Silu_for_9_else_else_else_if_acc_nl[25:0];
  assign Silu_for_9_else_else_else_if_acc_itm_25_1_1 = readslicef_26_25_1(Silu_for_9_else_else_else_if_acc_nl);
  assign act_regs_data_and_832_cse = ActUnitRun_wen & and_dcpl_1246 & and_dcpl_333
      & (~ act_config_is_zero_first_sva_dfm_4) & (z_out[4]);
  assign act_regs_data_and_2704_enex5 = act_regs_data_and_832_cse & (reg_act_port_read_out_data_0_14_sva_dfm_enexo
      | reg_act_port_read_out_data_0_6_sva_dfm_enexo | reg_act_port_read_out_data_0_13_sva_dfm_enexo
      | reg_act_port_read_out_data_0_0_sva_dfm_enexo | reg_act_port_read_out_data_0_5_sva_dfm_enexo
      | reg_act_port_read_out_data_0_15_sva_dfm_enexo | reg_act_port_read_out_data_0_1_sva_dfm_enexo
      | reg_act_port_read_out_data_0_4_sva_dfm_enexo | reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo
      | reg_act_port_read_out_data_0_8_sva_dfm_enexo | reg_act_port_read_out_data_0_11_sva_dfm_enexo
      | reg_act_regs_data_3_15_sva_dfm_2_30_26_enexo_1 | reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo
      | reg_act_port_read_out_data_0_3_sva_dfm_enexo | reg_act_port_read_out_data_0_7_sva_dfm_enexo
      | reg_act_port_read_out_data_0_12_sva_dfm_enexo | reg_act_port_read_out_data_0_2_sva_dfm_enexo
      | reg_act_port_read_out_data_0_10_sva_dfm_enexo | reg_act_port_read_out_data_0_9_sva_dfm_enexo);
  assign act_regs_data_and_2705_enex5 = act_regs_data_and_832_cse & (reg_act_port_read_out_data_0_3_sva_dfm_enexo_1
      | reg_act_port_read_out_data_0_10_sva_dfm_enexo_1 | reg_act_port_read_out_data_0_6_sva_dfm_enexo_1
      | reg_act_port_read_out_data_0_7_sva_dfm_enexo_1 | reg_act_port_read_out_data_0_11_sva_dfm_enexo_1
      | reg_act_regs_data_3_15_sva_dfm_2_25_22_enexo_1 | reg_act_port_read_out_data_0_1_sva_dfm_enexo_1
      | reg_act_port_read_out_data_0_5_sva_dfm_enexo_1 | reg_act_port_read_out_data_0_8_sva_dfm_enexo_1
      | reg_act_port_read_out_data_0_15_sva_dfm_enexo_1 | reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_1
      | reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_1 | reg_act_port_read_out_data_0_4_sva_dfm_enexo_1
      | reg_act_port_read_out_data_0_14_sva_dfm_enexo_1 | reg_act_port_read_out_data_0_0_sva_dfm_enexo_1
      | reg_act_port_read_out_data_0_12_sva_dfm_enexo_1 | reg_act_port_read_out_data_0_9_sva_dfm_enexo_1
      | reg_act_port_read_out_data_0_2_sva_dfm_enexo_1 | reg_act_port_read_out_data_0_13_sva_dfm_enexo_1);
  assign act_regs_data_and_2706_enex5 = act_regs_data_and_832_cse & (reg_act_port_read_out_data_0_0_sva_dfm_enexo_2
      | reg_act_port_read_out_data_0_11_sva_dfm_enexo_2 | reg_act_port_read_out_data_0_9_sva_dfm_enexo_2
      | reg_act_port_read_out_data_0_14_sva_dfm_enexo_2 | reg_act_port_read_out_data_0_8_sva_dfm_enexo_2
      | reg_act_port_read_out_data_0_15_sva_dfm_enexo_2 | reg_act_regs_data_3_15_sva_dfm_2_21_0_enexo_1
      | reg_act_port_read_out_data_0_13_sva_dfm_enexo_2 | reg_act_port_read_out_data_0_4_sva_dfm_enexo_2
      | reg_act_port_read_out_data_0_3_sva_dfm_enexo_2 | reg_act_port_read_out_data_0_10_sva_dfm_enexo_2
      | reg_act_port_read_out_data_0_1_sva_dfm_enexo_2 | reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_2
      | reg_act_port_read_out_data_0_2_sva_dfm_enexo_2 | reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_2
      | reg_act_port_read_out_data_0_12_sva_dfm_enexo_2 | reg_act_port_read_out_data_0_7_sva_dfm_enexo_2
      | reg_act_port_read_out_data_0_6_sva_dfm_enexo_2 | reg_act_port_read_out_data_0_5_sva_dfm_enexo_2);
  assign act_regs_data_and_2707_enex5 = act_regs_data_and_832_cse & (reg_act_port_read_out_data_0_1_sva_dfm_enexo_3
      | reg_act_port_read_out_data_0_9_sva_dfm_enexo_3 | reg_act_port_read_out_data_0_3_sva_dfm_enexo_3
      | reg_act_port_read_out_data_0_12_sva_dfm_enexo_3 | reg_act_port_read_out_data_0_4_sva_dfm_enexo_3
      | reg_act_regs_data_3_14_sva_dfm_2_30_26_enexo_1 | reg_act_port_read_out_data_0_14_sva_dfm_enexo_3
      | reg_act_port_read_out_data_0_2_sva_dfm_enexo_3 | reg_act_port_read_out_data_0_0_sva_dfm_enexo_3
      | reg_act_port_read_out_data_0_8_sva_dfm_enexo_3 | reg_act_port_read_out_data_0_7_sva_dfm_enexo_3
      | reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_3 | reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_3
      | reg_act_port_read_out_data_0_5_sva_dfm_enexo_3 | reg_act_port_read_out_data_0_13_sva_dfm_enexo_3
      | reg_act_port_read_out_data_0_6_sva_dfm_enexo_3 | reg_act_port_read_out_data_0_15_sva_dfm_enexo_3
      | reg_act_port_read_out_data_0_11_sva_dfm_enexo_3 | reg_act_port_read_out_data_0_10_sva_dfm_enexo_3);
  assign act_regs_data_and_2708_enex5 = act_regs_data_and_832_cse & (reg_act_port_read_out_data_0_8_sva_dfm_enexo_4
      | reg_act_port_read_out_data_0_5_sva_dfm_enexo_4 | reg_act_port_read_out_data_0_2_sva_dfm_enexo_4
      | reg_act_port_read_out_data_0_14_sva_dfm_enexo_4 | reg_act_port_read_out_data_0_7_sva_dfm_enexo_4
      | reg_act_port_read_out_data_0_15_sva_dfm_enexo_4 | reg_act_port_read_out_data_0_10_sva_dfm_enexo_4
      | reg_act_regs_data_3_14_sva_dfm_2_25_22_enexo_1 | reg_act_port_read_out_data_0_13_sva_dfm_enexo_4
      | reg_act_port_read_out_data_0_6_sva_dfm_enexo_4 | reg_act_port_read_out_data_0_11_sva_dfm_enexo_4
      | reg_act_port_read_out_data_0_4_sva_dfm_enexo_4 | reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_4
      | reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_4 | reg_act_port_read_out_data_0_12_sva_dfm_enexo_4
      | reg_act_port_read_out_data_0_0_sva_dfm_enexo_4 | reg_act_port_read_out_data_0_3_sva_dfm_enexo_4
      | reg_act_port_read_out_data_0_1_sva_dfm_enexo_4 | reg_act_port_read_out_data_0_9_sva_dfm_enexo_4);
  assign act_regs_data_and_2709_enex5 = act_regs_data_and_832_cse & (reg_act_port_read_out_data_0_11_sva_dfm_enexo_5
      | reg_act_port_read_out_data_0_5_sva_dfm_enexo_5 | reg_act_port_read_out_data_0_10_sva_dfm_enexo_5
      | reg_act_port_read_out_data_0_14_sva_dfm_enexo_5 | reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_5
      | reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_5 | reg_act_port_read_out_data_0_1_sva_dfm_enexo_5
      | reg_act_port_read_out_data_0_9_sva_dfm_enexo_5 | reg_act_port_read_out_data_0_3_sva_dfm_enexo_5
      | reg_act_port_read_out_data_0_12_sva_dfm_enexo_5 | reg_act_port_read_out_data_0_6_sva_dfm_enexo_5
      | reg_act_port_read_out_data_0_0_sva_dfm_enexo_5 | reg_act_port_read_out_data_0_8_sva_dfm_enexo_5
      | reg_act_port_read_out_data_0_2_sva_dfm_enexo_5 | reg_act_regs_data_3_14_sva_dfm_2_21_0_enexo_1
      | reg_act_port_read_out_data_0_4_sva_dfm_enexo_5 | reg_act_port_read_out_data_0_13_sva_dfm_enexo_5
      | reg_act_port_read_out_data_0_7_sva_dfm_enexo_5 | reg_act_port_read_out_data_0_15_sva_dfm_enexo_5);
  assign act_regs_data_and_2710_enex5 = act_regs_data_and_832_cse & (reg_act_port_read_out_data_0_3_sva_dfm_enexo_6
      | reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_6 | reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_6
      | reg_act_port_read_out_data_0_7_sva_dfm_enexo_6 | reg_act_port_read_out_data_0_15_sva_dfm_enexo_6
      | reg_act_port_read_out_data_0_0_sva_dfm_enexo_6 | reg_act_port_read_out_data_0_4_sva_dfm_enexo_6
      | reg_act_port_read_out_data_0_11_sva_dfm_enexo_6 | reg_act_regs_data_3_13_sva_dfm_2_30_26_enexo_1
      | reg_act_port_read_out_data_0_13_sva_dfm_enexo_6 | reg_act_port_read_out_data_0_6_sva_dfm_enexo_6
      | reg_act_port_read_out_data_0_5_sva_dfm_enexo_6 | reg_act_port_read_out_data_0_14_sva_dfm_enexo_6
      | reg_act_port_read_out_data_0_8_sva_dfm_enexo_6 | reg_act_port_read_out_data_0_12_sva_dfm_enexo_6
      | reg_act_port_read_out_data_0_2_sva_dfm_enexo_6 | reg_act_port_read_out_data_0_10_sva_dfm_enexo_6
      | reg_act_port_read_out_data_0_1_sva_dfm_enexo_6 | reg_act_port_read_out_data_0_9_sva_dfm_enexo_6);
  assign act_regs_data_and_2711_enex5 = act_regs_data_and_832_cse & (reg_act_port_read_out_data_0_10_sva_dfm_enexo_7
      | reg_act_regs_data_3_13_sva_dfm_2_25_22_enexo_1 | reg_act_port_read_out_data_0_15_sva_dfm_enexo_7
      | reg_act_port_read_out_data_0_2_sva_dfm_enexo_7 | reg_act_port_read_out_data_0_7_sva_dfm_enexo_7
      | reg_act_port_read_out_data_0_8_sva_dfm_enexo_7 | reg_act_port_read_out_data_0_6_sva_dfm_enexo_7
      | reg_act_port_read_out_data_0_13_sva_dfm_enexo_7 | reg_act_port_read_out_data_0_14_sva_dfm_enexo_7
      | reg_act_port_read_out_data_0_9_sva_dfm_enexo_7 | reg_act_port_read_out_data_0_4_sva_dfm_enexo_7
      | reg_act_port_read_out_data_0_11_sva_dfm_enexo_7 | reg_act_port_read_out_data_0_0_sva_dfm_enexo_7
      | reg_act_port_read_out_data_0_3_sva_dfm_enexo_7 | reg_act_port_read_out_data_0_12_sva_dfm_enexo_7
      | reg_act_port_read_out_data_0_5_sva_dfm_enexo_7 | reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_7
      | reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_7 | reg_act_port_read_out_data_0_1_sva_dfm_enexo_7);
  assign act_regs_data_and_2712_enex5 = act_regs_data_and_832_cse & (reg_act_port_read_out_data_0_8_sva_dfm_enexo_8
      | reg_act_port_read_out_data_0_12_sva_dfm_enexo_8 | reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_8
      | reg_act_port_read_out_data_0_7_sva_dfm_enexo_8 | reg_act_port_read_out_data_0_15_sva_dfm_enexo_8
      | reg_act_regs_data_3_13_sva_dfm_2_21_0_enexo_1 | reg_act_port_read_out_data_0_10_sva_dfm_enexo_8
      | reg_act_port_read_out_data_0_0_sva_dfm_enexo_8 | reg_act_port_read_out_data_0_2_sva_dfm_enexo_8
      | reg_act_port_read_out_data_0_3_sva_dfm_enexo_8 | reg_act_port_read_out_data_0_14_sva_dfm_enexo_8
      | reg_act_port_read_out_data_0_9_sva_dfm_enexo_8 | reg_act_port_read_out_data_0_5_sva_dfm_enexo_8
      | reg_act_port_read_out_data_0_4_sva_dfm_enexo_8 | reg_act_port_read_out_data_0_11_sva_dfm_enexo_8
      | reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_8 | reg_act_port_read_out_data_0_13_sva_dfm_enexo_8
      | reg_act_port_read_out_data_0_6_sva_dfm_enexo_8 | reg_act_port_read_out_data_0_1_sva_dfm_enexo_8);
  assign act_regs_data_and_2713_enex5 = act_regs_data_and_832_cse & (reg_act_port_read_out_data_0_8_sva_dfm_enexo_9
      | reg_act_port_read_out_data_0_6_sva_dfm_enexo_9 | reg_act_port_read_out_data_0_13_sva_dfm_enexo_9
      | reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_9 | reg_act_port_read_out_data_0_4_sva_dfm_enexo_9
      | reg_act_port_read_out_data_0_2_sva_dfm_enexo_9 | reg_act_port_read_out_data_0_7_sva_dfm_enexo_9
      | reg_act_port_read_out_data_0_5_sva_dfm_enexo_9 | reg_act_port_read_out_data_0_11_sva_dfm_enexo_9
      | reg_act_port_read_out_data_0_1_sva_dfm_enexo_9 | reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_9
      | reg_act_port_read_out_data_0_10_sva_dfm_enexo_9 | reg_act_port_read_out_data_0_15_sva_dfm_enexo_9
      | reg_act_port_read_out_data_0_9_sva_dfm_enexo_9 | reg_act_port_read_out_data_0_3_sva_dfm_enexo_9
      | reg_act_regs_data_3_12_sva_dfm_2_30_26_enexo_1 | reg_act_port_read_out_data_0_0_sva_dfm_enexo_9
      | reg_act_port_read_out_data_0_12_sva_dfm_enexo_9 | reg_act_port_read_out_data_0_14_sva_dfm_enexo_9);
  assign act_regs_data_and_2714_enex5 = act_regs_data_and_832_cse & (reg_act_port_read_out_data_0_13_sva_dfm_enexo_10
      | reg_act_port_read_out_data_0_10_sva_dfm_enexo_10 | reg_act_port_read_out_data_0_11_sva_dfm_enexo_10
      | reg_act_port_read_out_data_0_9_sva_dfm_enexo_10 | reg_act_port_read_out_data_0_0_sva_dfm_enexo_10
      | reg_act_port_read_out_data_0_5_sva_dfm_enexo_10 | reg_act_port_read_out_data_0_6_sva_dfm_enexo_10
      | reg_act_regs_data_3_12_sva_dfm_2_25_22_enexo_1 | reg_act_port_read_out_data_0_12_sva_dfm_enexo_10
      | reg_act_port_read_out_data_0_15_sva_dfm_enexo_10 | reg_act_port_read_out_data_0_7_sva_dfm_enexo_10
      | reg_act_port_read_out_data_0_2_sva_dfm_enexo_10 | reg_act_port_read_out_data_0_8_sva_dfm_enexo_10
      | reg_act_port_read_out_data_0_4_sva_dfm_enexo_10 | reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_10
      | reg_act_port_read_out_data_0_3_sva_dfm_enexo_10 | reg_act_port_read_out_data_0_1_sva_dfm_enexo_10
      | reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_10 | reg_act_port_read_out_data_0_14_sva_dfm_enexo_10);
  assign act_regs_data_and_2715_enex5 = act_regs_data_and_832_cse & (reg_act_port_read_out_data_0_8_sva_dfm_enexo_11
      | reg_act_port_read_out_data_0_7_sva_dfm_enexo_11 | reg_act_port_read_out_data_0_5_sva_dfm_enexo_11
      | reg_act_port_read_out_data_0_3_sva_dfm_enexo_11 | reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_11
      | reg_act_port_read_out_data_0_13_sva_dfm_enexo_11 | reg_act_port_read_out_data_0_10_sva_dfm_enexo_11
      | reg_act_port_read_out_data_0_6_sva_dfm_enexo_11 | reg_act_port_read_out_data_0_4_sva_dfm_enexo_11
      | reg_act_port_read_out_data_0_0_sva_dfm_enexo_11 | reg_act_regs_data_3_12_sva_dfm_2_21_0_enexo_1
      | reg_act_port_read_out_data_0_15_sva_dfm_enexo_11 | reg_act_port_read_out_data_0_11_sva_dfm_enexo_11
      | reg_act_port_read_out_data_0_9_sva_dfm_enexo_11 | reg_act_port_read_out_data_0_1_sva_dfm_enexo_11
      | reg_act_port_read_out_data_0_14_sva_dfm_enexo_11 | reg_act_port_read_out_data_0_12_sva_dfm_enexo_11
      | reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_11 | reg_act_port_read_out_data_0_2_sva_dfm_enexo_11);
  assign act_regs_data_and_2716_enex5 = act_regs_data_and_832_cse & (reg_act_port_read_out_data_0_12_sva_dfm_enexo_12
      | reg_act_port_read_out_data_0_3_sva_dfm_enexo_12 | reg_act_port_read_out_data_0_2_sva_dfm_enexo_12
      | reg_act_regs_data_3_11_sva_dfm_2_30_26_enexo_1 | reg_act_port_read_out_data_0_4_sva_dfm_enexo_12
      | reg_act_port_read_out_data_0_10_sva_dfm_enexo_12 | reg_act_port_read_out_data_0_9_sva_dfm_enexo_12
      | reg_act_port_read_out_data_0_1_sva_dfm_enexo_12 | reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_12
      | reg_act_port_read_out_data_0_14_sva_dfm_enexo_12 | reg_act_port_read_out_data_0_13_sva_dfm_enexo_12
      | reg_act_port_read_out_data_0_11_sva_dfm_enexo_12 | reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_12
      | reg_act_port_read_out_data_0_6_sva_dfm_enexo_12 | reg_act_port_read_out_data_0_0_sva_dfm_enexo_12
      | reg_act_port_read_out_data_0_8_sva_dfm_enexo_12 | reg_act_port_read_out_data_0_5_sva_dfm_enexo_12
      | reg_act_port_read_out_data_0_15_sva_dfm_enexo_12 | reg_act_port_read_out_data_0_7_sva_dfm_enexo_12);
  assign act_regs_data_and_2717_enex5 = act_regs_data_and_832_cse & (reg_act_port_read_out_data_0_11_sva_dfm_enexo_13
      | reg_act_port_read_out_data_0_5_sva_dfm_enexo_13 | reg_act_port_read_out_data_0_13_sva_dfm_enexo_13
      | reg_act_port_read_out_data_0_1_sva_dfm_enexo_13 | reg_act_port_read_out_data_0_4_sva_dfm_enexo_13
      | reg_act_port_read_out_data_0_2_sva_dfm_enexo_13 | reg_act_port_read_out_data_0_15_sva_dfm_enexo_13
      | reg_act_port_read_out_data_0_7_sva_dfm_enexo_13 | reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_13
      | reg_act_regs_data_3_11_sva_dfm_2_25_22_enexo_1 | reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_13
      | reg_act_port_read_out_data_0_3_sva_dfm_enexo_13 | reg_act_port_read_out_data_0_6_sva_dfm_enexo_13
      | reg_act_port_read_out_data_0_10_sva_dfm_enexo_13 | reg_act_port_read_out_data_0_8_sva_dfm_enexo_13
      | reg_act_port_read_out_data_0_9_sva_dfm_enexo_13 | reg_act_port_read_out_data_0_0_sva_dfm_enexo_13
      | reg_act_port_read_out_data_0_12_sva_dfm_enexo_13 | reg_act_port_read_out_data_0_14_sva_dfm_enexo_13);
  assign act_regs_data_and_2718_enex5 = act_regs_data_and_832_cse & (reg_act_port_read_out_data_0_2_sva_dfm_enexo_14
      | reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_14 | reg_act_port_read_out_data_0_1_sva_dfm_enexo_14
      | reg_act_port_read_out_data_0_9_sva_dfm_enexo_14 | reg_act_port_read_out_data_0_5_sva_dfm_enexo_14
      | reg_act_port_read_out_data_0_12_sva_dfm_enexo_14 | reg_act_port_read_out_data_0_3_sva_dfm_enexo_14
      | reg_act_port_read_out_data_0_14_sva_dfm_enexo_14 | reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_14
      | reg_act_port_read_out_data_0_0_sva_dfm_enexo_14 | reg_act_port_read_out_data_0_13_sva_dfm_enexo_14
      | reg_act_port_read_out_data_0_6_sva_dfm_enexo_14 | reg_act_port_read_out_data_0_10_sva_dfm_enexo_14
      | reg_act_port_read_out_data_0_15_sva_dfm_enexo_14 | reg_act_regs_data_3_11_sva_dfm_2_21_0_enexo_1
      | reg_act_port_read_out_data_0_7_sva_dfm_enexo_14 | reg_act_port_read_out_data_0_11_sva_dfm_enexo_14
      | reg_act_port_read_out_data_0_4_sva_dfm_enexo_14 | reg_act_port_read_out_data_0_8_sva_dfm_enexo_14);
  assign act_regs_data_and_2719_enex5 = act_regs_data_and_832_cse & (reg_act_port_read_out_data_0_5_sva_dfm_enexo_15
      | reg_act_port_read_out_data_0_13_sva_dfm_enexo_15 | reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_15
      | reg_act_port_read_out_data_0_15_sva_dfm_enexo_15 | reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_15
      | reg_act_port_read_out_data_0_11_sva_dfm_enexo_15 | reg_act_port_read_out_data_0_14_sva_dfm_enexo_15
      | reg_act_regs_data_3_10_sva_dfm_2_30_26_enexo_1 | reg_act_port_read_out_data_0_10_sva_dfm_enexo_15
      | reg_act_port_read_out_data_0_0_sva_dfm_enexo_15 | reg_act_port_read_out_data_0_4_sva_dfm_enexo_15
      | reg_act_port_read_out_data_0_12_sva_dfm_enexo_15 | reg_act_port_read_out_data_0_3_sva_dfm_enexo_15
      | reg_act_port_read_out_data_0_2_sva_dfm_enexo_15 | reg_act_port_read_out_data_0_7_sva_dfm_enexo_15
      | reg_act_port_read_out_data_0_6_sva_dfm_enexo_15 | reg_act_port_read_out_data_0_1_sva_dfm_enexo_15
      | reg_act_port_read_out_data_0_9_sva_dfm_enexo_15 | reg_act_port_read_out_data_0_8_sva_dfm_enexo_15);
  assign act_regs_data_and_2720_enex5 = act_regs_data_and_832_cse & (reg_act_port_read_out_data_0_12_sva_dfm_enexo_16
      | reg_act_port_read_out_data_0_4_sva_dfm_enexo_16 | reg_act_port_read_out_data_0_2_sva_dfm_enexo_16
      | reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_16 | reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_16
      | reg_act_port_read_out_data_0_14_sva_dfm_enexo_16 | reg_act_port_read_out_data_0_10_sva_dfm_enexo_16
      | reg_act_port_read_out_data_0_0_sva_dfm_enexo_16 | reg_act_port_read_out_data_0_6_sva_dfm_enexo_16
      | reg_act_port_read_out_data_0_11_sva_dfm_enexo_16 | reg_act_port_read_out_data_0_1_sva_dfm_enexo_16
      | reg_act_port_read_out_data_0_3_sva_dfm_enexo_16 | reg_act_port_read_out_data_0_5_sva_dfm_enexo_16
      | reg_act_port_read_out_data_0_15_sva_dfm_enexo_16 | reg_act_port_read_out_data_0_8_sva_dfm_enexo_16
      | reg_act_port_read_out_data_0_9_sva_dfm_enexo_16 | reg_act_port_read_out_data_0_13_sva_dfm_enexo_16
      | reg_act_regs_data_3_10_sva_dfm_2_25_22_enexo_1 | reg_act_port_read_out_data_0_7_sva_dfm_enexo_16);
  assign act_regs_data_and_2721_enex5 = act_regs_data_and_832_cse & (reg_act_port_read_out_data_0_14_sva_dfm_enexo_17
      | reg_act_port_read_out_data_0_4_sva_dfm_enexo_17 | reg_act_port_read_out_data_0_5_sva_dfm_enexo_17
      | reg_act_port_read_out_data_0_8_sva_dfm_enexo_17 | reg_act_port_read_out_data_0_10_sva_dfm_enexo_17
      | reg_act_regs_data_3_10_sva_dfm_2_21_0_enexo_1 | reg_act_port_read_out_data_0_15_sva_dfm_enexo_17
      | reg_act_port_read_out_data_0_13_sva_dfm_enexo_17 | reg_act_port_read_out_data_0_12_sva_dfm_enexo_17
      | reg_act_port_read_out_data_0_9_sva_dfm_enexo_17 | reg_act_port_read_out_data_0_7_sva_dfm_enexo_17
      | reg_act_port_read_out_data_0_3_sva_dfm_enexo_17 | reg_act_port_read_out_data_0_11_sva_dfm_enexo_17
      | reg_act_port_read_out_data_0_0_sva_dfm_enexo_17 | reg_act_port_read_out_data_0_6_sva_dfm_enexo_17
      | reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_17 | reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_17
      | reg_act_port_read_out_data_0_2_sva_dfm_enexo_17 | reg_act_port_read_out_data_0_1_sva_dfm_enexo_17);
  assign act_regs_data_and_2722_enex5 = act_regs_data_and_832_cse & (reg_act_port_read_out_data_0_14_sva_dfm_enexo_18
      | reg_act_port_read_out_data_0_2_sva_dfm_enexo_18 | reg_act_port_read_out_data_0_8_sva_dfm_enexo_18
      | reg_act_port_read_out_data_0_10_sva_dfm_enexo_18 | reg_act_port_read_out_data_0_6_sva_dfm_enexo_18
      | reg_act_port_read_out_data_0_4_sva_dfm_enexo_18 | reg_act_port_read_out_data_0_11_sva_dfm_enexo_18
      | reg_act_port_read_out_data_0_12_sva_dfm_enexo_18 | reg_act_port_read_out_data_0_13_sva_dfm_enexo_18
      | reg_act_port_read_out_data_0_0_sva_dfm_enexo_18 | reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_18
      | reg_act_port_read_out_data_0_5_sva_dfm_enexo_18 | reg_act_port_read_out_data_0_15_sva_dfm_enexo_18
      | reg_act_port_read_out_data_0_9_sva_dfm_enexo_18 | reg_act_port_read_out_data_0_1_sva_dfm_enexo_18
      | reg_act_port_read_out_data_0_7_sva_dfm_enexo_18 | reg_act_port_read_out_data_0_3_sva_dfm_enexo_18
      | reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_18 | reg_act_regs_data_3_9_sva_dfm_2_30_26_enexo_1);
  assign act_regs_data_and_2723_enex5 = act_regs_data_and_832_cse & (reg_act_port_read_out_data_0_14_sva_dfm_enexo_19
      | reg_act_port_read_out_data_0_11_sva_dfm_enexo_19 | reg_act_port_read_out_data_0_12_sva_dfm_enexo_19
      | reg_act_port_read_out_data_0_2_sva_dfm_enexo_19 | reg_act_port_read_out_data_0_13_sva_dfm_enexo_19
      | reg_act_port_read_out_data_0_8_sva_dfm_enexo_19 | reg_act_port_read_out_data_0_15_sva_dfm_enexo_19
      | reg_act_port_read_out_data_0_7_sva_dfm_enexo_19 | reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_19
      | reg_act_port_read_out_data_0_4_sva_dfm_enexo_19 | reg_act_port_read_out_data_0_0_sva_dfm_enexo_19
      | reg_act_port_read_out_data_0_6_sva_dfm_enexo_19 | reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_19
      | reg_act_port_read_out_data_0_9_sva_dfm_enexo_19 | reg_act_port_read_out_data_0_1_sva_dfm_enexo_19
      | reg_act_regs_data_3_9_sva_dfm_2_25_22_enexo_1 | reg_act_port_read_out_data_0_5_sva_dfm_enexo_19
      | reg_act_port_read_out_data_0_10_sva_dfm_enexo_19 | reg_act_port_read_out_data_0_3_sva_dfm_enexo_19);
  assign act_regs_data_and_2724_enex5 = act_regs_data_and_832_cse & (reg_act_port_read_out_data_0_6_sva_dfm_enexo_20
      | reg_act_port_read_out_data_0_7_sva_dfm_enexo_20 | reg_act_port_read_out_data_0_15_sva_dfm_enexo_20
      | reg_act_port_read_out_data_0_3_sva_dfm_enexo_20 | reg_act_port_read_out_data_0_10_sva_dfm_enexo_20
      | reg_act_port_read_out_data_0_11_sva_dfm_enexo_20 | reg_act_port_read_out_data_0_4_sva_dfm_enexo_20
      | reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_20 | reg_act_port_read_out_data_0_14_sva_dfm_enexo_20
      | reg_act_port_read_out_data_0_0_sva_dfm_enexo_20 | reg_act_port_read_out_data_0_8_sva_dfm_enexo_20
      | reg_act_regs_data_3_9_sva_dfm_2_21_0_enexo_1 | reg_act_port_read_out_data_0_2_sva_dfm_enexo_20
      | reg_act_port_read_out_data_0_5_sva_dfm_enexo_20 | reg_act_port_read_out_data_0_12_sva_dfm_enexo_20
      | reg_act_port_read_out_data_0_13_sva_dfm_enexo_20 | reg_act_port_read_out_data_0_1_sva_dfm_enexo_20
      | reg_act_port_read_out_data_0_9_sva_dfm_enexo_20 | reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_20);
  assign act_regs_data_and_2725_enex5 = act_regs_data_and_832_cse & (reg_act_port_read_out_data_0_11_sva_dfm_enexo_21
      | reg_act_port_read_out_data_0_8_sva_dfm_enexo_21 | reg_act_port_read_out_data_0_12_sva_dfm_enexo_21
      | reg_act_port_read_out_data_0_9_sva_dfm_enexo_21 | reg_act_port_read_out_data_0_13_sva_dfm_enexo_21
      | reg_act_port_read_out_data_0_2_sva_dfm_enexo_21 | reg_act_port_read_out_data_0_4_sva_dfm_enexo_21
      | reg_act_port_read_out_data_0_15_sva_dfm_enexo_21 | reg_act_port_read_out_data_0_6_sva_dfm_enexo_21
      | reg_act_port_read_out_data_0_10_sva_dfm_enexo_21 | reg_act_port_read_out_data_0_0_sva_dfm_enexo_21
      | reg_act_port_read_out_data_0_1_sva_dfm_enexo_21 | reg_act_port_read_out_data_0_3_sva_dfm_enexo_21
      | reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_21 | reg_act_port_read_out_data_0_14_sva_dfm_enexo_21
      | reg_act_regs_data_3_8_sva_dfm_2_30_26_enexo_1 | reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_21
      | reg_act_port_read_out_data_0_5_sva_dfm_enexo_21 | reg_act_port_read_out_data_0_7_sva_dfm_enexo_21);
  assign act_regs_data_and_2726_enex5 = act_regs_data_and_832_cse & (reg_act_port_read_out_data_0_11_sva_dfm_enexo_22
      | reg_act_port_read_out_data_0_10_sva_dfm_enexo_22 | reg_act_port_read_out_data_0_6_sva_dfm_enexo_22
      | reg_act_port_read_out_data_0_1_sva_dfm_enexo_22 | reg_act_port_read_out_data_0_9_sva_dfm_enexo_22
      | reg_act_port_read_out_data_0_3_sva_dfm_enexo_22 | reg_act_port_read_out_data_0_12_sva_dfm_enexo_22
      | reg_act_port_read_out_data_0_0_sva_dfm_enexo_22 | reg_act_port_read_out_data_0_8_sva_dfm_enexo_22
      | reg_act_port_read_out_data_0_15_sva_dfm_enexo_22 | reg_act_port_read_out_data_0_7_sva_dfm_enexo_22
      | reg_act_port_read_out_data_0_5_sva_dfm_enexo_22 | reg_act_port_read_out_data_0_2_sva_dfm_enexo_22
      | reg_act_port_read_out_data_0_14_sva_dfm_enexo_22 | reg_act_port_read_out_data_0_4_sva_dfm_enexo_22
      | reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_22 | reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_22
      | reg_act_regs_data_3_8_sva_dfm_2_25_22_enexo_1 | reg_act_port_read_out_data_0_13_sva_dfm_enexo_22);
  assign act_regs_data_and_2727_enex5 = act_regs_data_and_832_cse & (reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_23
      | reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_23 | reg_act_port_read_out_data_0_1_sva_dfm_enexo_23
      | reg_act_port_read_out_data_0_9_sva_dfm_enexo_23 | reg_act_port_read_out_data_0_3_sva_dfm_enexo_23
      | reg_act_port_read_out_data_0_12_sva_dfm_enexo_23 | reg_act_port_read_out_data_0_0_sva_dfm_enexo_23
      | reg_act_port_read_out_data_0_8_sva_dfm_enexo_23 | reg_act_port_read_out_data_0_7_sva_dfm_enexo_23
      | reg_act_port_read_out_data_0_15_sva_dfm_enexo_23 | reg_act_port_read_out_data_0_2_sva_dfm_enexo_23
      | reg_act_regs_data_3_8_sva_dfm_2_21_0_enexo_1 | reg_act_port_read_out_data_0_4_sva_dfm_enexo_23
      | reg_act_port_read_out_data_0_14_sva_dfm_enexo_23 | reg_act_port_read_out_data_0_11_sva_dfm_enexo_23
      | reg_act_port_read_out_data_0_10_sva_dfm_enexo_23 | reg_act_port_read_out_data_0_13_sva_dfm_enexo_23
      | reg_act_port_read_out_data_0_6_sva_dfm_enexo_23 | reg_act_port_read_out_data_0_5_sva_dfm_enexo_23);
  assign act_regs_data_and_2728_enex5 = act_regs_data_and_832_cse & (reg_act_port_read_out_data_0_4_sva_dfm_enexo_24
      | reg_act_port_read_out_data_0_12_sva_dfm_enexo_24 | reg_act_port_read_out_data_0_14_sva_dfm_enexo_24
      | reg_act_port_read_out_data_0_2_sva_dfm_enexo_24 | reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_24
      | reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_24 | reg_act_port_read_out_data_0_0_sva_dfm_enexo_24
      | reg_act_port_read_out_data_0_8_sva_dfm_enexo_24 | reg_act_port_read_out_data_0_7_sva_dfm_enexo_24
      | reg_act_port_read_out_data_0_15_sva_dfm_enexo_24 | reg_act_port_read_out_data_0_11_sva_dfm_enexo_24
      | reg_act_port_read_out_data_0_10_sva_dfm_enexo_24 | reg_act_port_read_out_data_0_13_sva_dfm_enexo_24
      | reg_act_port_read_out_data_0_6_sva_dfm_enexo_24 | reg_act_port_read_out_data_0_5_sva_dfm_enexo_24
      | reg_act_port_read_out_data_0_3_sva_dfm_enexo_24 | reg_act_regs_data_3_7_sva_dfm_2_30_26_enexo_1
      | reg_act_port_read_out_data_0_1_sva_dfm_enexo_24 | reg_act_port_read_out_data_0_9_sva_dfm_enexo_24);
  assign act_regs_data_and_2729_enex5 = act_regs_data_and_832_cse & (reg_act_port_read_out_data_0_2_sva_dfm_enexo_25
      | reg_act_port_read_out_data_0_5_sva_dfm_enexo_25 | reg_act_port_read_out_data_0_3_sva_dfm_enexo_25
      | reg_act_port_read_out_data_0_10_sva_dfm_enexo_25 | reg_act_port_read_out_data_0_11_sva_dfm_enexo_25
      | reg_act_port_read_out_data_0_1_sva_dfm_enexo_25 | reg_act_port_read_out_data_0_15_sva_dfm_enexo_25
      | reg_act_port_read_out_data_0_7_sva_dfm_enexo_25 | reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_25
      | reg_act_port_read_out_data_0_14_sva_dfm_enexo_25 | reg_act_port_read_out_data_0_4_sva_dfm_enexo_25
      | reg_act_port_read_out_data_0_12_sva_dfm_enexo_25 | reg_act_regs_data_3_7_sva_dfm_2_25_22_enexo_1
      | reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_25 | reg_act_port_read_out_data_0_8_sva_dfm_enexo_25
      | reg_act_port_read_out_data_0_9_sva_dfm_enexo_25 | reg_act_port_read_out_data_0_0_sva_dfm_enexo_25
      | reg_act_port_read_out_data_0_6_sva_dfm_enexo_25 | reg_act_port_read_out_data_0_13_sva_dfm_enexo_25);
  assign act_regs_data_and_2730_enex5 = act_regs_data_and_832_cse & (reg_act_port_read_out_data_0_14_sva_dfm_enexo_26
      | reg_act_port_read_out_data_0_4_sva_dfm_enexo_26 | reg_act_port_read_out_data_0_1_sva_dfm_enexo_26
      | reg_act_port_read_out_data_0_3_sva_dfm_enexo_26 | reg_act_port_read_out_data_0_15_sva_dfm_enexo_26
      | reg_act_port_read_out_data_0_2_sva_dfm_enexo_26 | reg_act_port_read_out_data_0_7_sva_dfm_enexo_26
      | reg_act_port_read_out_data_0_8_sva_dfm_enexo_26 | reg_act_port_read_out_data_0_9_sva_dfm_enexo_26
      | reg_act_port_read_out_data_0_11_sva_dfm_enexo_26 | reg_act_port_read_out_data_0_0_sva_dfm_enexo_26
      | reg_act_port_read_out_data_0_5_sva_dfm_enexo_26 | reg_act_regs_data_3_7_sva_dfm_2_21_0_enexo_1
      | reg_act_port_read_out_data_0_10_sva_dfm_enexo_26 | reg_act_port_read_out_data_0_12_sva_dfm_enexo_26
      | reg_act_port_read_out_data_0_13_sva_dfm_enexo_26 | reg_act_port_read_out_data_0_6_sva_dfm_enexo_26
      | reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_26 | reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_26);
  assign act_regs_data_and_2731_enex5 = act_regs_data_and_832_cse & (reg_act_port_read_out_data_0_13_sva_dfm_enexo_27
      | reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_27 | reg_act_port_read_out_data_0_1_sva_dfm_enexo_27
      | reg_act_port_read_out_data_0_6_sva_dfm_enexo_27 | reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_27
      | reg_act_port_read_out_data_0_12_sva_dfm_enexo_27 | reg_act_port_read_out_data_0_3_sva_dfm_enexo_27
      | reg_act_port_read_out_data_0_4_sva_dfm_enexo_27 | reg_act_port_read_out_data_0_2_sva_dfm_enexo_27
      | reg_act_port_read_out_data_0_10_sva_dfm_enexo_27 | reg_act_port_read_out_data_0_9_sva_dfm_enexo_27
      | reg_act_port_read_out_data_0_8_sva_dfm_enexo_27 | reg_act_port_read_out_data_0_0_sva_dfm_enexo_27
      | reg_act_port_read_out_data_0_7_sva_dfm_enexo_27 | reg_act_port_read_out_data_0_11_sva_dfm_enexo_27
      | reg_act_port_read_out_data_0_15_sva_dfm_enexo_27 | reg_act_port_read_out_data_0_14_sva_dfm_enexo_27
      | reg_act_regs_data_3_6_sva_dfm_2_30_26_enexo_1 | reg_act_port_read_out_data_0_5_sva_dfm_enexo_27);
  assign act_regs_data_and_2732_enex5 = act_regs_data_and_832_cse & (reg_act_port_read_out_data_0_4_sva_dfm_enexo_28
      | reg_act_port_read_out_data_0_2_sva_dfm_enexo_28 | reg_act_port_read_out_data_0_9_sva_dfm_enexo_28
      | reg_act_port_read_out_data_0_11_sva_dfm_enexo_28 | reg_act_port_read_out_data_0_12_sva_dfm_enexo_28
      | reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_28 | reg_act_port_read_out_data_0_3_sva_dfm_enexo_28
      | reg_act_port_read_out_data_0_8_sva_dfm_enexo_28 | reg_act_regs_data_3_6_sva_dfm_2_25_22_enexo_1
      | reg_act_port_read_out_data_0_6_sva_dfm_enexo_28 | reg_act_port_read_out_data_0_0_sva_dfm_enexo_28
      | reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_28 | reg_act_port_read_out_data_0_15_sva_dfm_enexo_28
      | reg_act_port_read_out_data_0_7_sva_dfm_enexo_28 | reg_act_port_read_out_data_0_10_sva_dfm_enexo_28
      | reg_act_port_read_out_data_0_14_sva_dfm_enexo_28 | reg_act_port_read_out_data_0_5_sva_dfm_enexo_28
      | reg_act_port_read_out_data_0_1_sva_dfm_enexo_28 | reg_act_port_read_out_data_0_13_sva_dfm_enexo_28);
  assign act_regs_data_and_2733_enex5 = act_regs_data_and_832_cse & (reg_act_port_read_out_data_0_0_sva_dfm_enexo_29
      | reg_act_regs_data_3_6_sva_dfm_2_21_0_enexo_1 | reg_act_port_read_out_data_0_9_sva_dfm_enexo_29
      | reg_act_port_read_out_data_0_5_sva_dfm_enexo_29 | reg_act_port_read_out_data_0_10_sva_dfm_enexo_29
      | reg_act_port_read_out_data_0_14_sva_dfm_enexo_29 | reg_act_port_read_out_data_0_4_sva_dfm_enexo_29
      | reg_act_port_read_out_data_0_2_sva_dfm_enexo_29 | reg_act_port_read_out_data_0_15_sva_dfm_enexo_29
      | reg_act_port_read_out_data_0_11_sva_dfm_enexo_29 | reg_act_port_read_out_data_0_3_sva_dfm_enexo_29
      | reg_act_port_read_out_data_0_13_sva_dfm_enexo_29 | reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_29
      | reg_act_port_read_out_data_0_8_sva_dfm_enexo_29 | reg_act_port_read_out_data_0_12_sva_dfm_enexo_29
      | reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_29 | reg_act_port_read_out_data_0_1_sva_dfm_enexo_29
      | reg_act_port_read_out_data_0_6_sva_dfm_enexo_29 | reg_act_port_read_out_data_0_7_sva_dfm_enexo_29);
  assign act_regs_data_and_2734_enex5 = act_regs_data_and_832_cse & (reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_30
      | reg_act_port_read_out_data_0_14_sva_dfm_enexo_30 | reg_act_port_read_out_data_0_7_sva_dfm_enexo_30
      | reg_act_port_read_out_data_0_4_sva_dfm_enexo_30 | reg_act_port_read_out_data_0_8_sva_dfm_enexo_30
      | reg_act_port_read_out_data_0_10_sva_dfm_enexo_30 | reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_30
      | reg_act_port_read_out_data_0_11_sva_dfm_enexo_30 | reg_act_port_read_out_data_0_6_sva_dfm_enexo_30
      | reg_act_port_read_out_data_0_5_sva_dfm_enexo_30 | reg_act_port_read_out_data_0_3_sva_dfm_enexo_30
      | reg_act_port_read_out_data_0_13_sva_dfm_enexo_30 | reg_act_port_read_out_data_0_12_sva_dfm_enexo_30
      | reg_act_regs_data_3_5_sva_dfm_2_30_26_enexo_1 | reg_act_port_read_out_data_0_15_sva_dfm_enexo_30
      | reg_act_port_read_out_data_0_9_sva_dfm_enexo_30 | reg_act_port_read_out_data_0_1_sva_dfm_enexo_30
      | reg_act_port_read_out_data_0_0_sva_dfm_enexo_30 | reg_act_port_read_out_data_0_2_sva_dfm_enexo_30);
  assign act_regs_data_and_2735_enex5 = act_regs_data_and_832_cse & (reg_act_port_read_out_data_0_4_sva_dfm_enexo_31
      | reg_act_port_read_out_data_0_11_sva_dfm_enexo_31 | reg_act_port_read_out_data_0_3_sva_dfm_enexo_31
      | reg_act_port_read_out_data_0_1_sva_dfm_enexo_31 | reg_act_port_read_out_data_0_5_sva_dfm_enexo_31
      | reg_act_port_read_out_data_0_7_sva_dfm_enexo_31 | reg_act_port_read_out_data_0_8_sva_dfm_enexo_31
      | reg_act_port_read_out_data_0_13_sva_dfm_enexo_31 | reg_act_port_read_out_data_0_6_sva_dfm_enexo_31
      | reg_act_port_read_out_data_0_15_sva_dfm_enexo_31 | reg_act_regs_data_3_5_sva_dfm_2_25_22_enexo_1
      | reg_act_port_read_out_data_0_10_sva_dfm_enexo_31 | reg_act_port_read_out_data_0_9_sva_dfm_enexo_31
      | reg_act_port_read_out_data_0_12_sva_dfm_enexo_31 | reg_act_port_read_out_data_0_0_sva_dfm_enexo_31
      | reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_31 | reg_act_port_read_out_data_0_14_sva_dfm_enexo_31
      | reg_act_port_read_out_data_0_2_sva_dfm_enexo_31 | reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_31);
  assign act_regs_data_and_2736_enex5 = act_regs_data_and_832_cse & (reg_act_port_read_out_data_0_8_sva_dfm_enexo_32
      | reg_act_port_read_out_data_0_13_sva_dfm_enexo_32 | reg_act_port_read_out_data_0_6_sva_dfm_enexo_32
      | reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_32 | reg_act_port_read_out_data_0_12_sva_dfm_enexo_32
      | reg_act_port_read_out_data_0_9_sva_dfm_enexo_32 | reg_act_port_read_out_data_0_1_sva_dfm_enexo_32
      | reg_act_port_read_out_data_0_5_sva_dfm_enexo_32 | reg_act_port_read_out_data_0_7_sva_dfm_enexo_32
      | reg_act_port_read_out_data_0_3_sva_dfm_enexo_32 | reg_act_port_read_out_data_0_2_sva_dfm_enexo_32
      | reg_act_port_read_out_data_0_0_sva_dfm_enexo_32 | reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_32
      | reg_act_port_read_out_data_0_4_sva_dfm_enexo_32 | reg_act_regs_data_3_5_sva_dfm_2_21_0_enexo_1
      | reg_act_port_read_out_data_0_11_sva_dfm_enexo_32 | reg_act_port_read_out_data_0_10_sva_dfm_enexo_32
      | reg_act_port_read_out_data_0_15_sva_dfm_enexo_32 | reg_act_port_read_out_data_0_14_sva_dfm_enexo_32);
  assign act_regs_data_and_2737_enex5 = act_regs_data_and_832_cse & (reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_33
      | reg_act_port_read_out_data_0_5_sva_dfm_enexo_33 | reg_act_port_read_out_data_0_10_sva_dfm_enexo_33
      | reg_act_port_read_out_data_0_6_sva_dfm_enexo_33 | reg_act_port_read_out_data_0_0_sva_dfm_enexo_33
      | reg_act_port_read_out_data_0_14_sva_dfm_enexo_33 | reg_act_port_read_out_data_0_7_sva_dfm_enexo_33
      | reg_act_port_read_out_data_0_15_sva_dfm_enexo_33 | reg_act_port_read_out_data_0_11_sva_dfm_enexo_33
      | reg_act_port_read_out_data_0_4_sva_dfm_enexo_33 | reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_33
      | reg_act_port_read_out_data_0_8_sva_dfm_enexo_33 | reg_act_port_read_out_data_0_1_sva_dfm_enexo_33
      | reg_act_port_read_out_data_0_12_sva_dfm_enexo_33 | reg_act_port_read_out_data_0_3_sva_dfm_enexo_33
      | reg_act_port_read_out_data_0_2_sva_dfm_enexo_33 | reg_act_port_read_out_data_0_13_sva_dfm_enexo_33
      | reg_act_port_read_out_data_0_9_sva_dfm_enexo_33 | reg_act_regs_data_3_4_sva_dfm_2_30_26_enexo_1);
  assign act_regs_data_and_2738_enex5 = act_regs_data_and_832_cse & (reg_act_port_read_out_data_0_14_sva_dfm_enexo_34
      | reg_act_port_read_out_data_0_4_sva_dfm_enexo_34 | reg_act_port_read_out_data_0_9_sva_dfm_enexo_34
      | reg_act_port_read_out_data_0_2_sva_dfm_enexo_34 | reg_act_port_read_out_data_0_15_sva_dfm_enexo_34
      | reg_act_port_read_out_data_0_11_sva_dfm_enexo_34 | reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_34
      | reg_act_port_read_out_data_0_1_sva_dfm_enexo_34 | reg_act_port_read_out_data_0_0_sva_dfm_enexo_34
      | reg_act_port_read_out_data_0_8_sva_dfm_enexo_34 | reg_act_regs_data_3_4_sva_dfm_2_25_22_enexo_1
      | reg_act_port_read_out_data_0_12_sva_dfm_enexo_34 | reg_act_port_read_out_data_0_10_sva_dfm_enexo_34
      | reg_act_port_read_out_data_0_6_sva_dfm_enexo_34 | reg_act_port_read_out_data_0_7_sva_dfm_enexo_34
      | reg_act_port_read_out_data_0_3_sva_dfm_enexo_34 | reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_34
      | reg_act_port_read_out_data_0_5_sva_dfm_enexo_34 | reg_act_port_read_out_data_0_13_sva_dfm_enexo_34);
  assign act_regs_data_and_2739_enex5 = act_regs_data_and_832_cse & (reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_35
      | reg_act_port_read_out_data_0_10_sva_dfm_enexo_35 | reg_act_port_read_out_data_0_4_sva_dfm_enexo_35
      | reg_act_port_read_out_data_0_14_sva_dfm_enexo_35 | reg_act_port_read_out_data_0_13_sva_dfm_enexo_35
      | reg_act_port_read_out_data_0_15_sva_dfm_enexo_35 | reg_act_port_read_out_data_0_12_sva_dfm_enexo_35
      | reg_act_port_read_out_data_0_0_sva_dfm_enexo_35 | reg_act_port_read_out_data_0_8_sva_dfm_enexo_35
      | reg_act_port_read_out_data_0_1_sva_dfm_enexo_35 | reg_act_port_read_out_data_0_7_sva_dfm_enexo_35
      | reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_35 | reg_act_port_read_out_data_0_11_sva_dfm_enexo_35
      | reg_act_port_read_out_data_0_2_sva_dfm_enexo_35 | reg_act_regs_data_3_4_sva_dfm_2_21_0_enexo_1
      | reg_act_port_read_out_data_0_6_sva_dfm_enexo_35 | reg_act_port_read_out_data_0_9_sva_dfm_enexo_35
      | reg_act_port_read_out_data_0_3_sva_dfm_enexo_35 | reg_act_port_read_out_data_0_5_sva_dfm_enexo_35);
  assign act_regs_data_and_2740_enex5 = act_regs_data_and_832_cse & (reg_act_regs_data_3_3_sva_dfm_2_30_26_enexo_1
      | reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_36 | reg_act_port_read_out_data_0_6_sva_dfm_enexo_36
      | reg_act_port_read_out_data_0_2_sva_dfm_enexo_36 | reg_act_port_read_out_data_0_3_sva_dfm_enexo_36
      | reg_act_port_read_out_data_0_4_sva_dfm_enexo_36 | reg_act_port_read_out_data_0_5_sva_dfm_enexo_36
      | reg_act_port_read_out_data_0_9_sva_dfm_enexo_36 | reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_36
      | reg_act_port_read_out_data_0_1_sva_dfm_enexo_36 | reg_act_port_read_out_data_0_14_sva_dfm_enexo_36
      | reg_act_port_read_out_data_0_15_sva_dfm_enexo_36 | reg_act_port_read_out_data_0_11_sva_dfm_enexo_36
      | reg_act_port_read_out_data_0_13_sva_dfm_enexo_36 | reg_act_port_read_out_data_0_10_sva_dfm_enexo_36
      | reg_act_port_read_out_data_0_12_sva_dfm_enexo_36 | reg_act_port_read_out_data_0_7_sva_dfm_enexo_36
      | reg_act_port_read_out_data_0_0_sva_dfm_enexo_36 | reg_act_port_read_out_data_0_8_sva_dfm_enexo_36);
  assign act_regs_data_and_2741_enex5 = act_regs_data_and_832_cse & (reg_act_port_read_out_data_0_14_sva_dfm_enexo_37
      | reg_act_port_read_out_data_0_2_sva_dfm_enexo_37 | reg_act_port_read_out_data_0_4_sva_dfm_enexo_37
      | reg_act_regs_data_3_3_sva_dfm_2_25_22_enexo_1 | reg_act_port_read_out_data_0_13_sva_dfm_enexo_37
      | reg_act_port_read_out_data_0_11_sva_dfm_enexo_37 | reg_act_port_read_out_data_0_10_sva_dfm_enexo_37
      | reg_act_port_read_out_data_0_6_sva_dfm_enexo_37 | reg_act_port_read_out_data_0_5_sva_dfm_enexo_37
      | reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_37 | reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_37
      | reg_act_port_read_out_data_0_1_sva_dfm_enexo_37 | reg_act_port_read_out_data_0_3_sva_dfm_enexo_37
      | reg_act_port_read_out_data_0_15_sva_dfm_enexo_37 | reg_act_port_read_out_data_0_9_sva_dfm_enexo_37
      | reg_act_port_read_out_data_0_12_sva_dfm_enexo_37 | reg_act_port_read_out_data_0_8_sva_dfm_enexo_37
      | reg_act_port_read_out_data_0_0_sva_dfm_enexo_37 | reg_act_port_read_out_data_0_7_sva_dfm_enexo_37);
  assign act_regs_data_and_2742_enex5 = act_regs_data_and_832_cse & (reg_act_port_read_out_data_0_11_sva_dfm_enexo_38
      | reg_act_regs_data_3_3_sva_dfm_2_21_0_enexo_1 | reg_act_port_read_out_data_0_10_sva_dfm_enexo_38
      | reg_act_port_read_out_data_0_4_sva_dfm_enexo_38 | reg_act_port_read_out_data_0_9_sva_dfm_enexo_38
      | reg_act_port_read_out_data_0_7_sva_dfm_enexo_38 | reg_act_port_read_out_data_0_13_sva_dfm_enexo_38
      | reg_act_port_read_out_data_0_8_sva_dfm_enexo_38 | reg_act_port_read_out_data_0_3_sva_dfm_enexo_38
      | reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_38 | reg_act_port_read_out_data_0_12_sva_dfm_enexo_38
      | reg_act_port_read_out_data_0_14_sva_dfm_enexo_38 | reg_act_port_read_out_data_0_6_sva_dfm_enexo_38
      | reg_act_port_read_out_data_0_0_sva_dfm_enexo_38 | reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_38
      | reg_act_port_read_out_data_0_5_sva_dfm_enexo_38 | reg_act_port_read_out_data_0_15_sva_dfm_enexo_38
      | reg_act_port_read_out_data_0_1_sva_dfm_enexo_38 | reg_act_port_read_out_data_0_2_sva_dfm_enexo_38);
  assign act_regs_data_and_2743_enex5 = act_regs_data_and_832_cse & (reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_39
      | reg_act_port_read_out_data_0_0_sva_dfm_enexo_39 | reg_act_port_read_out_data_0_5_sva_dfm_enexo_39
      | reg_act_port_read_out_data_0_14_sva_dfm_enexo_39 | reg_act_port_read_out_data_0_13_sva_dfm_enexo_39
      | reg_act_port_read_out_data_0_7_sva_dfm_enexo_39 | reg_act_port_read_out_data_0_3_sva_dfm_enexo_39
      | reg_act_port_read_out_data_0_11_sva_dfm_enexo_39 | reg_act_port_read_out_data_0_9_sva_dfm_enexo_39
      | reg_act_port_read_out_data_0_6_sva_dfm_enexo_39 | reg_act_port_read_out_data_0_12_sva_dfm_enexo_39
      | reg_act_port_read_out_data_0_2_sva_dfm_enexo_39 | reg_act_port_read_out_data_0_15_sva_dfm_enexo_39
      | reg_act_port_read_out_data_0_8_sva_dfm_enexo_39 | reg_act_regs_data_3_2_sva_dfm_2_30_26_enexo_1
      | reg_act_port_read_out_data_0_1_sva_dfm_enexo_39 | reg_act_port_read_out_data_0_4_sva_dfm_enexo_39
      | reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_39 | reg_act_port_read_out_data_0_10_sva_dfm_enexo_39);
  assign act_regs_data_and_2744_enex5 = act_regs_data_and_832_cse & (reg_act_port_read_out_data_0_9_sva_dfm_enexo_40
      | reg_act_port_read_out_data_0_1_sva_dfm_enexo_40 | reg_act_regs_data_3_2_sva_dfm_2_25_22_enexo_1
      | reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_40 | reg_act_port_read_out_data_0_5_sva_dfm_enexo_40
      | reg_act_port_read_out_data_0_11_sva_dfm_enexo_40 | reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_40
      | reg_act_port_read_out_data_0_14_sva_dfm_enexo_40 | reg_act_port_read_out_data_0_15_sva_dfm_enexo_40
      | reg_act_port_read_out_data_0_7_sva_dfm_enexo_40 | reg_act_port_read_out_data_0_0_sva_dfm_enexo_40
      | reg_act_port_read_out_data_0_12_sva_dfm_enexo_40 | reg_act_port_read_out_data_0_3_sva_dfm_enexo_40
      | reg_act_port_read_out_data_0_6_sva_dfm_enexo_40 | reg_act_port_read_out_data_0_8_sva_dfm_enexo_40
      | reg_act_port_read_out_data_0_4_sva_dfm_enexo_40 | reg_act_port_read_out_data_0_13_sva_dfm_enexo_40
      | reg_act_port_read_out_data_0_2_sva_dfm_enexo_40 | reg_act_port_read_out_data_0_10_sva_dfm_enexo_40);
  assign act_regs_data_and_2745_enex5 = act_regs_data_and_832_cse & (reg_act_port_read_out_data_0_11_sva_dfm_enexo_41
      | reg_act_port_read_out_data_0_12_sva_dfm_enexo_41 | reg_act_port_read_out_data_0_0_sva_dfm_enexo_41
      | reg_act_port_read_out_data_0_6_sva_dfm_enexo_41 | reg_act_port_read_out_data_0_5_sva_dfm_enexo_41
      | reg_act_port_read_out_data_0_9_sva_dfm_enexo_41 | reg_act_port_read_out_data_0_13_sva_dfm_enexo_41
      | reg_act_regs_data_3_2_sva_dfm_2_21_0_enexo_1 | reg_act_port_read_out_data_0_10_sva_dfm_enexo_41
      | reg_act_port_read_out_data_0_15_sva_dfm_enexo_41 | reg_act_port_read_out_data_0_14_sva_dfm_enexo_41
      | reg_act_port_read_out_data_0_8_sva_dfm_enexo_41 | reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_41
      | reg_act_port_read_out_data_0_2_sva_dfm_enexo_41 | reg_act_port_read_out_data_0_4_sva_dfm_enexo_41
      | reg_act_port_read_out_data_0_3_sva_dfm_enexo_41 | reg_act_port_read_out_data_0_7_sva_dfm_enexo_41
      | reg_act_port_read_out_data_0_1_sva_dfm_enexo_41 | reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_41);
  assign act_regs_data_and_2746_enex5 = act_regs_data_and_832_cse & (reg_act_port_read_out_data_0_5_sva_dfm_enexo_42
      | reg_act_port_read_out_data_0_10_sva_dfm_enexo_42 | reg_act_regs_data_3_1_sva_dfm_2_30_26_enexo_1
      | reg_act_port_read_out_data_0_4_sva_dfm_enexo_42 | reg_act_port_read_out_data_0_2_sva_dfm_enexo_42
      | reg_act_port_read_out_data_0_14_sva_dfm_enexo_42 | reg_act_port_read_out_data_0_13_sva_dfm_enexo_42
      | reg_act_port_read_out_data_0_8_sva_dfm_enexo_42 | reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_42
      | reg_act_port_read_out_data_0_9_sva_dfm_enexo_42 | reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_42
      | reg_act_port_read_out_data_0_0_sva_dfm_enexo_42 | reg_act_port_read_out_data_0_3_sva_dfm_enexo_42
      | reg_act_port_read_out_data_0_7_sva_dfm_enexo_42 | reg_act_port_read_out_data_0_12_sva_dfm_enexo_42
      | reg_act_port_read_out_data_0_6_sva_dfm_enexo_42 | reg_act_port_read_out_data_0_11_sva_dfm_enexo_42
      | reg_act_port_read_out_data_0_1_sva_dfm_enexo_42 | reg_act_port_read_out_data_0_15_sva_dfm_enexo_42);
  assign act_regs_data_and_2747_enex5 = act_regs_data_and_832_cse & (reg_act_port_read_out_data_0_9_sva_dfm_enexo_43
      | reg_act_port_read_out_data_0_3_sva_dfm_enexo_43 | reg_act_port_read_out_data_0_12_sva_dfm_enexo_43
      | reg_act_port_read_out_data_0_0_sva_dfm_enexo_43 | reg_act_port_read_out_data_0_8_sva_dfm_enexo_43
      | reg_act_port_read_out_data_0_5_sva_dfm_enexo_43 | reg_act_port_read_out_data_0_4_sva_dfm_enexo_43
      | reg_act_port_read_out_data_0_7_sva_dfm_enexo_43 | reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_43
      | reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_43 | reg_act_port_read_out_data_0_1_sva_dfm_enexo_43
      | reg_act_port_read_out_data_0_2_sva_dfm_enexo_43 | reg_act_port_read_out_data_0_13_sva_dfm_enexo_43
      | reg_act_port_read_out_data_0_14_sva_dfm_enexo_43 | reg_act_port_read_out_data_0_15_sva_dfm_enexo_43
      | reg_act_regs_data_3_1_sva_dfm_2_25_22_enexo_1 | reg_act_port_read_out_data_0_10_sva_dfm_enexo_43
      | reg_act_port_read_out_data_0_6_sva_dfm_enexo_43 | reg_act_port_read_out_data_0_11_sva_dfm_enexo_43);
  assign act_regs_data_and_2748_enex5 = act_regs_data_and_832_cse & (reg_act_port_read_out_data_0_14_sva_dfm_enexo_44
      | reg_act_port_read_out_data_0_8_sva_dfm_enexo_44 | reg_act_port_read_out_data_0_2_sva_dfm_enexo_44
      | reg_act_port_read_out_data_0_9_sva_dfm_enexo_44 | reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_44
      | reg_act_port_read_out_data_0_0_sva_dfm_enexo_44 | reg_act_port_read_out_data_0_5_sva_dfm_enexo_44
      | reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_44 | reg_act_port_read_out_data_0_6_sva_dfm_enexo_44
      | reg_act_port_read_out_data_0_3_sva_dfm_enexo_44 | reg_act_port_read_out_data_0_13_sva_dfm_enexo_44
      | reg_act_regs_data_3_1_sva_dfm_2_21_0_enexo_1 | reg_act_port_read_out_data_0_12_sva_dfm_enexo_44
      | reg_act_port_read_out_data_0_10_sva_dfm_enexo_44 | reg_act_port_read_out_data_0_11_sva_dfm_enexo_44
      | reg_act_port_read_out_data_0_4_sva_dfm_enexo_44 | reg_act_port_read_out_data_0_7_sva_dfm_enexo_44
      | reg_act_port_read_out_data_0_1_sva_dfm_enexo_44 | reg_act_port_read_out_data_0_15_sva_dfm_enexo_44);
  assign act_regs_data_or_64_nl = (and_dcpl_1267 & and_dcpl_1266 & and_dcpl_1265)
      | and_dcpl_1270;
  assign act_regs_data_mux_320_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_64_nl, and_dcpl_1246);
  assign act_regs_data_and_124_cse = ActUnitRun_wen & act_regs_data_mux_320_nl &
      mux_450_itm;
  assign act_regs_data_and_892_cse = (~ and_dcpl_1270) & and_dcpl_1246;
  assign act_regs_data_and_893_cse = and_dcpl_1270 & and_dcpl_1246;
  assign act_regs_data_or_65_nl = (and_dcpl_1275 & and_dcpl_1272) | and_dcpl_1277;
  assign act_regs_data_mux_324_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_65_nl, and_dcpl_1246);
  assign act_regs_data_and_128_cse = ActUnitRun_wen & act_regs_data_mux_324_nl &
      mux_450_itm;
  assign act_regs_data_and_898_cse = (~ and_dcpl_1277) & and_dcpl_1246;
  assign act_regs_data_and_899_cse = and_dcpl_1277 & and_dcpl_1246;
  assign act_regs_data_or_66_nl = (and_dcpl_1275 & and_dcpl_1278) | and_dcpl_1280;
  assign act_regs_data_mux_328_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_66_nl, and_dcpl_1246);
  assign act_regs_data_and_132_cse = ActUnitRun_wen & act_regs_data_mux_328_nl &
      mux_450_itm;
  assign act_regs_data_and_904_cse = (~ and_dcpl_1280) & and_dcpl_1246;
  assign act_regs_data_and_905_cse = and_dcpl_1280 & and_dcpl_1246;
  assign act_regs_data_or_67_nl = (and_dcpl_1275 & and_dcpl_1282) | and_dcpl_1284;
  assign act_regs_data_mux_332_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_67_nl, and_dcpl_1246);
  assign act_regs_data_and_136_cse = ActUnitRun_wen & act_regs_data_mux_332_nl &
      mux_450_itm;
  assign act_regs_data_and_910_cse = (~ and_dcpl_1284) & and_dcpl_1246;
  assign act_regs_data_and_911_cse = and_dcpl_1284 & and_dcpl_1246;
  assign act_regs_data_or_68_nl = (and_dcpl_1275 & and_dcpl_1285) | and_dcpl_1287;
  assign act_regs_data_mux_336_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_68_nl, and_dcpl_1246);
  assign act_regs_data_and_140_cse = ActUnitRun_wen & act_regs_data_mux_336_nl &
      mux_450_itm;
  assign act_regs_data_and_916_cse = (~ and_dcpl_1287) & and_dcpl_1246;
  assign act_regs_data_and_917_cse = and_dcpl_1287 & and_dcpl_1246;
  assign act_regs_data_or_69_nl = (and_dcpl_1275 & and_dcpl_1289) | and_dcpl_1291;
  assign act_regs_data_mux_340_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_69_nl, and_dcpl_1246);
  assign act_regs_data_and_144_cse = ActUnitRun_wen & act_regs_data_mux_340_nl &
      mux_450_itm;
  assign act_regs_data_and_922_cse = (~ and_dcpl_1291) & and_dcpl_1246;
  assign act_regs_data_and_923_cse = and_dcpl_1291 & and_dcpl_1246;
  assign act_regs_data_or_70_nl = (and_dcpl_1275 & and_dcpl_1292) | and_dcpl_1294;
  assign act_regs_data_mux_344_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_70_nl, and_dcpl_1246);
  assign act_regs_data_and_148_cse = ActUnitRun_wen & act_regs_data_mux_344_nl &
      mux_450_itm;
  assign act_regs_data_and_928_cse = (~ and_dcpl_1294) & and_dcpl_1246;
  assign act_regs_data_and_929_cse = and_dcpl_1294 & and_dcpl_1246;
  assign act_regs_data_or_71_nl = (and_dcpl_1275 & and_dcpl_1295) | and_dcpl_1297;
  assign act_regs_data_mux_348_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_71_nl, and_dcpl_1246);
  assign act_regs_data_and_152_cse = ActUnitRun_wen & act_regs_data_mux_348_nl &
      mux_450_itm;
  assign act_regs_data_and_934_cse = (~ and_dcpl_1297) & and_dcpl_1246;
  assign act_regs_data_and_935_cse = and_dcpl_1297 & and_dcpl_1246;
  assign act_regs_data_or_72_nl = (and_dcpl_1275 & and_dcpl_1265) | and_dcpl_1299;
  assign act_regs_data_mux_352_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_72_nl, and_dcpl_1246);
  assign act_regs_data_and_156_cse = ActUnitRun_wen & act_regs_data_mux_352_nl &
      mux_450_itm;
  assign act_regs_data_and_940_cse = (~ and_dcpl_1299) & and_dcpl_1246;
  assign act_regs_data_and_941_cse = and_dcpl_1299 & and_dcpl_1246;
  assign act_regs_data_or_73_nl = (and_dcpl_1300 & and_dcpl_1272) | and_dcpl_1302;
  assign act_regs_data_mux_356_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_73_nl, and_dcpl_1246);
  assign act_regs_data_and_160_cse = ActUnitRun_wen & act_regs_data_mux_356_nl &
      mux_450_itm;
  assign act_regs_data_and_946_cse = (~ and_dcpl_1302) & and_dcpl_1246;
  assign act_regs_data_and_947_cse = and_dcpl_1302 & and_dcpl_1246;
  assign act_regs_data_or_74_nl = (and_dcpl_1300 & and_dcpl_1278) | and_dcpl_1304;
  assign act_regs_data_mux_360_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_74_nl, and_dcpl_1246);
  assign act_regs_data_and_164_cse = ActUnitRun_wen & act_regs_data_mux_360_nl &
      mux_450_itm;
  assign act_regs_data_and_952_cse = (~ and_dcpl_1304) & and_dcpl_1246;
  assign act_regs_data_and_953_cse = and_dcpl_1304 & and_dcpl_1246;
  assign act_regs_data_or_75_nl = (and_dcpl_1300 & and_dcpl_1282) | and_dcpl_1306;
  assign act_regs_data_mux_364_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_75_nl, and_dcpl_1246);
  assign act_regs_data_and_168_cse = ActUnitRun_wen & act_regs_data_mux_364_nl &
      mux_450_itm;
  assign act_regs_data_and_958_cse = (~ and_dcpl_1306) & and_dcpl_1246;
  assign act_regs_data_and_959_cse = and_dcpl_1306 & and_dcpl_1246;
  assign act_regs_data_or_76_nl = (and_dcpl_1300 & and_dcpl_1285) | and_dcpl_1308;
  assign act_regs_data_mux_368_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_76_nl, and_dcpl_1246);
  assign act_regs_data_and_172_cse = ActUnitRun_wen & act_regs_data_mux_368_nl &
      mux_450_itm;
  assign act_regs_data_and_964_cse = (~ and_dcpl_1308) & and_dcpl_1246;
  assign act_regs_data_and_965_cse = and_dcpl_1308 & and_dcpl_1246;
  assign act_regs_data_or_77_nl = (and_dcpl_1300 & and_dcpl_1289) | and_dcpl_1310;
  assign act_regs_data_mux_372_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_77_nl, and_dcpl_1246);
  assign act_regs_data_and_176_cse = ActUnitRun_wen & act_regs_data_mux_372_nl &
      mux_450_itm;
  assign act_regs_data_and_970_cse = (~ and_dcpl_1310) & and_dcpl_1246;
  assign act_regs_data_and_971_cse = and_dcpl_1310 & and_dcpl_1246;
  assign act_regs_data_or_78_nl = (and_dcpl_1300 & and_dcpl_1292) | and_dcpl_1312;
  assign act_regs_data_mux_376_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_78_nl, and_dcpl_1246);
  assign act_regs_data_and_180_cse = ActUnitRun_wen & act_regs_data_mux_376_nl &
      mux_450_itm;
  assign act_regs_data_and_976_cse = (~ and_dcpl_1312) & and_dcpl_1246;
  assign act_regs_data_and_977_cse = and_dcpl_1312 & and_dcpl_1246;
  assign act_regs_data_or_79_nl = (and_dcpl_1300 & and_dcpl_1295) | and_dcpl_1314;
  assign act_regs_data_mux_380_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_79_nl, and_dcpl_1246);
  assign act_regs_data_and_184_cse = ActUnitRun_wen & act_regs_data_mux_380_nl &
      mux_450_itm;
  assign act_regs_data_and_982_cse = (~ and_dcpl_1314) & and_dcpl_1246;
  assign act_regs_data_and_983_cse = and_dcpl_1314 & and_dcpl_1246;
  assign act_regs_data_or_80_nl = (and_dcpl_1300 & and_dcpl_1265) | and_dcpl_1316;
  assign act_regs_data_mux_384_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_80_nl, and_dcpl_1246);
  assign act_regs_data_and_188_cse = ActUnitRun_wen & act_regs_data_mux_384_nl &
      mux_450_itm;
  assign act_regs_data_and_988_cse = (~ and_dcpl_1316) & and_dcpl_1246;
  assign act_regs_data_and_989_cse = and_dcpl_1316 & and_dcpl_1246;
  assign act_regs_data_or_81_nl = (and_dcpl_1318 & and_dcpl_1272) | and_dcpl_1320;
  assign act_regs_data_mux_388_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_81_nl, and_dcpl_1246);
  assign act_regs_data_and_192_cse = ActUnitRun_wen & act_regs_data_mux_388_nl &
      mux_450_itm;
  assign act_regs_data_and_994_cse = (~ and_dcpl_1320) & and_dcpl_1246;
  assign act_regs_data_and_995_cse = and_dcpl_1320 & and_dcpl_1246;
  assign act_regs_data_or_82_nl = (and_dcpl_1318 & and_dcpl_1278) | and_dcpl_1322;
  assign act_regs_data_mux_392_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_82_nl, and_dcpl_1246);
  assign act_regs_data_and_196_cse = ActUnitRun_wen & act_regs_data_mux_392_nl &
      mux_450_itm;
  assign act_regs_data_and_1000_cse = (~ and_dcpl_1322) & and_dcpl_1246;
  assign act_regs_data_and_1001_cse = and_dcpl_1322 & and_dcpl_1246;
  assign act_regs_data_or_83_nl = (and_dcpl_1318 & and_dcpl_1282) | and_dcpl_1324;
  assign act_regs_data_mux_396_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_83_nl, and_dcpl_1246);
  assign act_regs_data_and_200_cse = ActUnitRun_wen & act_regs_data_mux_396_nl &
      mux_450_itm;
  assign act_regs_data_and_1006_cse = (~ and_dcpl_1324) & and_dcpl_1246;
  assign act_regs_data_and_1007_cse = and_dcpl_1324 & and_dcpl_1246;
  assign act_regs_data_or_84_nl = (and_dcpl_1318 & and_dcpl_1285) | and_dcpl_1326;
  assign act_regs_data_mux_400_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_84_nl, and_dcpl_1246);
  assign act_regs_data_and_204_cse = ActUnitRun_wen & act_regs_data_mux_400_nl &
      mux_450_itm;
  assign act_regs_data_and_1012_cse = (~ and_dcpl_1326) & and_dcpl_1246;
  assign act_regs_data_and_1013_cse = and_dcpl_1326 & and_dcpl_1246;
  assign act_regs_data_or_85_nl = (and_dcpl_1318 & and_dcpl_1289) | and_dcpl_1328;
  assign act_regs_data_mux_404_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_85_nl, and_dcpl_1246);
  assign act_regs_data_and_208_cse = ActUnitRun_wen & act_regs_data_mux_404_nl &
      mux_450_itm;
  assign act_regs_data_and_1018_cse = (~ and_dcpl_1328) & and_dcpl_1246;
  assign act_regs_data_and_1019_cse = and_dcpl_1328 & and_dcpl_1246;
  assign act_regs_data_or_86_nl = (and_dcpl_1318 & and_dcpl_1292) | and_dcpl_1330;
  assign act_regs_data_mux_408_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_86_nl, and_dcpl_1246);
  assign act_regs_data_and_212_cse = ActUnitRun_wen & act_regs_data_mux_408_nl &
      mux_450_itm;
  assign act_regs_data_and_1024_cse = (~ and_dcpl_1330) & and_dcpl_1246;
  assign act_regs_data_and_1025_cse = and_dcpl_1330 & and_dcpl_1246;
  assign act_regs_data_or_87_nl = (and_dcpl_1318 & and_dcpl_1295) | and_dcpl_1332;
  assign act_regs_data_mux_412_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_87_nl, and_dcpl_1246);
  assign act_regs_data_and_216_cse = ActUnitRun_wen & act_regs_data_mux_412_nl &
      mux_450_itm;
  assign act_regs_data_and_1030_cse = (~ and_dcpl_1332) & and_dcpl_1246;
  assign act_regs_data_and_1031_cse = and_dcpl_1332 & and_dcpl_1246;
  assign act_regs_data_or_88_nl = (and_dcpl_1318 & and_dcpl_1265) | and_dcpl_1334;
  assign act_regs_data_mux_416_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_88_nl, and_dcpl_1246);
  assign act_regs_data_and_220_cse = ActUnitRun_wen & act_regs_data_mux_416_nl &
      mux_450_itm;
  assign act_regs_data_and_1036_cse = (~ and_dcpl_1334) & and_dcpl_1246;
  assign act_regs_data_and_1037_cse = and_dcpl_1334 & and_dcpl_1246;
  assign act_regs_data_or_89_nl = (and_dcpl_1336 & and_dcpl_1272) | and_dcpl_1338;
  assign act_regs_data_mux_420_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_89_nl, and_dcpl_1246);
  assign act_regs_data_and_224_cse = ActUnitRun_wen & act_regs_data_mux_420_nl &
      mux_450_itm;
  assign act_regs_data_and_1042_cse = (~ and_dcpl_1338) & and_dcpl_1246;
  assign act_regs_data_and_1043_cse = and_dcpl_1338 & and_dcpl_1246;
  assign act_regs_data_or_90_nl = (and_dcpl_1336 & and_dcpl_1278) | and_dcpl_1340;
  assign act_regs_data_mux_424_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_90_nl, and_dcpl_1246);
  assign act_regs_data_and_228_cse = ActUnitRun_wen & act_regs_data_mux_424_nl &
      mux_450_itm;
  assign act_regs_data_and_1048_cse = (~ and_dcpl_1340) & and_dcpl_1246;
  assign act_regs_data_and_1049_cse = and_dcpl_1340 & and_dcpl_1246;
  assign act_regs_data_or_91_nl = (and_dcpl_1336 & and_dcpl_1282) | and_dcpl_1342;
  assign act_regs_data_mux_428_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_91_nl, and_dcpl_1246);
  assign act_regs_data_and_232_cse = ActUnitRun_wen & act_regs_data_mux_428_nl &
      mux_450_itm;
  assign act_regs_data_and_1054_cse = (~ and_dcpl_1342) & and_dcpl_1246;
  assign act_regs_data_and_1055_cse = and_dcpl_1342 & and_dcpl_1246;
  assign act_regs_data_or_92_nl = (and_dcpl_1336 & and_dcpl_1285) | and_dcpl_1344;
  assign act_regs_data_mux_432_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_92_nl, and_dcpl_1246);
  assign act_regs_data_and_236_cse = ActUnitRun_wen & act_regs_data_mux_432_nl &
      mux_450_itm;
  assign act_regs_data_and_1060_cse = (~ and_dcpl_1344) & and_dcpl_1246;
  assign act_regs_data_and_1061_cse = and_dcpl_1344 & and_dcpl_1246;
  assign act_regs_data_or_93_nl = (and_dcpl_1336 & and_dcpl_1289) | and_dcpl_1346;
  assign act_regs_data_mux_436_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_93_nl, and_dcpl_1246);
  assign act_regs_data_and_240_cse = ActUnitRun_wen & act_regs_data_mux_436_nl &
      mux_450_itm;
  assign act_regs_data_and_1066_cse = (~ and_dcpl_1346) & and_dcpl_1246;
  assign act_regs_data_and_1067_cse = and_dcpl_1346 & and_dcpl_1246;
  assign act_regs_data_or_94_nl = (and_dcpl_1336 & and_dcpl_1292) | and_dcpl_1348;
  assign act_regs_data_mux_440_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_94_nl, and_dcpl_1246);
  assign act_regs_data_and_244_cse = ActUnitRun_wen & act_regs_data_mux_440_nl &
      mux_450_itm;
  assign act_regs_data_and_1072_cse = (~ and_dcpl_1348) & and_dcpl_1246;
  assign act_regs_data_and_1073_cse = and_dcpl_1348 & and_dcpl_1246;
  assign act_regs_data_or_95_nl = (and_dcpl_1336 & and_dcpl_1295) | and_dcpl_1350;
  assign act_regs_data_mux_444_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_95_nl, and_dcpl_1246);
  assign act_regs_data_and_248_cse = ActUnitRun_wen & act_regs_data_mux_444_nl &
      mux_450_itm;
  assign act_regs_data_and_1078_cse = (~ and_dcpl_1350) & and_dcpl_1246;
  assign act_regs_data_and_1079_cse = and_dcpl_1350 & and_dcpl_1246;
  assign act_regs_data_or_96_nl = (and_dcpl_1336 & and_dcpl_1265) | and_dcpl_1352;
  assign act_regs_data_mux_448_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_96_nl, and_dcpl_1246);
  assign act_regs_data_and_252_cse = ActUnitRun_wen & act_regs_data_mux_448_nl &
      mux_450_itm;
  assign act_regs_data_and_1084_cse = (~ and_dcpl_1352) & and_dcpl_1246;
  assign act_regs_data_and_1085_cse = and_dcpl_1352 & and_dcpl_1246;
  assign act_regs_data_or_97_nl = (and_dcpl_1353 & and_dcpl_1272) | and_dcpl_1355;
  assign act_regs_data_mux_452_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_97_nl, and_dcpl_1246);
  assign act_regs_data_and_256_cse = ActUnitRun_wen & act_regs_data_mux_452_nl &
      mux_450_itm;
  assign act_regs_data_and_1090_cse = (~ and_dcpl_1355) & and_dcpl_1246;
  assign act_regs_data_and_1091_cse = and_dcpl_1355 & and_dcpl_1246;
  assign act_regs_data_or_98_nl = (and_dcpl_1353 & and_dcpl_1278) | and_dcpl_1357;
  assign act_regs_data_mux_456_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_98_nl, and_dcpl_1246);
  assign act_regs_data_and_260_cse = ActUnitRun_wen & act_regs_data_mux_456_nl &
      mux_450_itm;
  assign act_regs_data_and_1096_cse = (~ and_dcpl_1357) & and_dcpl_1246;
  assign act_regs_data_and_1097_cse = and_dcpl_1357 & and_dcpl_1246;
  assign act_regs_data_or_99_nl = (and_dcpl_1353 & and_dcpl_1282) | and_dcpl_1359;
  assign act_regs_data_mux_460_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_99_nl, and_dcpl_1246);
  assign act_regs_data_and_264_cse = ActUnitRun_wen & act_regs_data_mux_460_nl &
      mux_450_itm;
  assign act_regs_data_and_1102_cse = (~ and_dcpl_1359) & and_dcpl_1246;
  assign act_regs_data_and_1103_cse = and_dcpl_1359 & and_dcpl_1246;
  assign act_regs_data_or_100_nl = (and_dcpl_1353 & and_dcpl_1285) | and_dcpl_1361;
  assign act_regs_data_mux_464_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_100_nl, and_dcpl_1246);
  assign act_regs_data_and_268_cse = ActUnitRun_wen & act_regs_data_mux_464_nl &
      mux_450_itm;
  assign act_regs_data_and_1108_cse = (~ and_dcpl_1361) & and_dcpl_1246;
  assign act_regs_data_and_1109_cse = and_dcpl_1361 & and_dcpl_1246;
  assign act_regs_data_or_101_nl = (and_dcpl_1353 & and_dcpl_1289) | and_dcpl_1363;
  assign act_regs_data_mux_468_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_101_nl, and_dcpl_1246);
  assign act_regs_data_and_272_cse = ActUnitRun_wen & act_regs_data_mux_468_nl &
      mux_450_itm;
  assign act_regs_data_and_1114_cse = (~ and_dcpl_1363) & and_dcpl_1246;
  assign act_regs_data_and_1115_cse = and_dcpl_1363 & and_dcpl_1246;
  assign act_regs_data_or_102_nl = (and_dcpl_1353 & and_dcpl_1292) | and_dcpl_1365;
  assign act_regs_data_mux_472_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_102_nl, and_dcpl_1246);
  assign act_regs_data_and_276_cse = ActUnitRun_wen & act_regs_data_mux_472_nl &
      mux_450_itm;
  assign act_regs_data_and_1120_cse = (~ and_dcpl_1365) & and_dcpl_1246;
  assign act_regs_data_and_1121_cse = and_dcpl_1365 & and_dcpl_1246;
  assign act_regs_data_or_103_nl = (and_dcpl_1353 & and_dcpl_1295) | and_dcpl_1367;
  assign act_regs_data_mux_476_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_103_nl, and_dcpl_1246);
  assign act_regs_data_and_280_cse = ActUnitRun_wen & act_regs_data_mux_476_nl &
      mux_450_itm;
  assign act_regs_data_and_1126_cse = (~ and_dcpl_1367) & and_dcpl_1246;
  assign act_regs_data_and_1127_cse = and_dcpl_1367 & and_dcpl_1246;
  assign act_regs_data_or_104_nl = (and_dcpl_1353 & and_dcpl_1265) | and_dcpl_1369;
  assign act_regs_data_mux_480_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_104_nl, and_dcpl_1246);
  assign act_regs_data_and_284_cse = ActUnitRun_wen & act_regs_data_mux_480_nl &
      mux_450_itm;
  assign act_regs_data_and_1132_cse = (~ and_dcpl_1369) & and_dcpl_1246;
  assign act_regs_data_and_1133_cse = and_dcpl_1369 & and_dcpl_1246;
  assign act_regs_data_or_105_nl = (and_dcpl_1370 & and_dcpl_1272) | and_dcpl_1372;
  assign act_regs_data_mux_484_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_105_nl, and_dcpl_1246);
  assign act_regs_data_and_288_cse = ActUnitRun_wen & act_regs_data_mux_484_nl &
      mux_450_itm;
  assign act_regs_data_and_1138_cse = (~ and_dcpl_1372) & and_dcpl_1246;
  assign act_regs_data_and_1139_cse = and_dcpl_1372 & and_dcpl_1246;
  assign act_regs_data_or_106_nl = (and_dcpl_1370 & and_dcpl_1278) | and_dcpl_1374;
  assign act_regs_data_mux_488_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_106_nl, and_dcpl_1246);
  assign act_regs_data_and_292_cse = ActUnitRun_wen & act_regs_data_mux_488_nl &
      mux_450_itm;
  assign act_regs_data_and_1144_cse = (~ and_dcpl_1374) & and_dcpl_1246;
  assign act_regs_data_and_1145_cse = and_dcpl_1374 & and_dcpl_1246;
  assign act_regs_data_or_107_nl = (and_dcpl_1370 & and_dcpl_1282) | and_dcpl_1376;
  assign act_regs_data_mux_492_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_107_nl, and_dcpl_1246);
  assign act_regs_data_and_296_cse = ActUnitRun_wen & act_regs_data_mux_492_nl &
      mux_450_itm;
  assign act_regs_data_and_1150_cse = (~ and_dcpl_1376) & and_dcpl_1246;
  assign act_regs_data_and_1151_cse = and_dcpl_1376 & and_dcpl_1246;
  assign act_regs_data_or_108_nl = (and_dcpl_1370 & and_dcpl_1285) | and_dcpl_1378;
  assign act_regs_data_mux_496_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_108_nl, and_dcpl_1246);
  assign act_regs_data_and_300_cse = ActUnitRun_wen & act_regs_data_mux_496_nl &
      mux_450_itm;
  assign act_regs_data_and_1156_cse = (~ and_dcpl_1378) & and_dcpl_1246;
  assign act_regs_data_and_1157_cse = and_dcpl_1378 & and_dcpl_1246;
  assign act_regs_data_or_109_nl = (and_dcpl_1370 & and_dcpl_1289) | and_dcpl_1380;
  assign act_regs_data_mux_500_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_109_nl, and_dcpl_1246);
  assign act_regs_data_and_304_cse = ActUnitRun_wen & act_regs_data_mux_500_nl &
      mux_450_itm;
  assign act_regs_data_and_1162_cse = (~ and_dcpl_1380) & and_dcpl_1246;
  assign act_regs_data_and_1163_cse = and_dcpl_1380 & and_dcpl_1246;
  assign act_regs_data_or_110_nl = (and_dcpl_1370 & and_dcpl_1292) | and_dcpl_1382;
  assign act_regs_data_mux_504_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_110_nl, and_dcpl_1246);
  assign act_regs_data_and_308_cse = ActUnitRun_wen & act_regs_data_mux_504_nl &
      mux_450_itm;
  assign act_regs_data_and_1168_cse = (~ and_dcpl_1382) & and_dcpl_1246;
  assign act_regs_data_and_1169_cse = and_dcpl_1382 & and_dcpl_1246;
  assign act_regs_data_or_111_nl = (and_dcpl_1370 & and_dcpl_1295) | and_dcpl_1384;
  assign act_regs_data_mux_508_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_111_nl, and_dcpl_1246);
  assign act_regs_data_and_312_cse = ActUnitRun_wen & act_regs_data_mux_508_nl &
      mux_450_itm;
  assign act_regs_data_and_1174_cse = (~ and_dcpl_1384) & and_dcpl_1246;
  assign act_regs_data_and_1175_cse = and_dcpl_1384 & and_dcpl_1246;
  assign act_regs_data_or_112_nl = (and_dcpl_1370 & and_dcpl_1265) | and_dcpl_1386;
  assign act_regs_data_mux_512_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_regs_data_or_112_nl, and_dcpl_1246);
  assign act_regs_data_and_316_cse = ActUnitRun_wen & act_regs_data_mux_512_nl &
      mux_450_itm;
  assign act_regs_data_and_1180_cse = (~ and_dcpl_1386) & and_dcpl_1246;
  assign act_regs_data_and_1181_cse = and_dcpl_1386 & and_dcpl_1246;
  assign and_2363_nl = (fsm_output[2]) & (fsm_output[0]);
  assign or_1866_nl = (fsm_output[2]) | (fsm_output[0]);
  assign mux_746_cse = MUX_s_1_2_2(and_2363_nl, or_1866_nl, fsm_output[1]);
  assign and_2364_cse = or_3395_cse & (fsm_output[0]);
  assign and_2367_cse = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0==4'b1011);
  assign or_1872_cse = (fsm_output[1:0]!=2'b00);
  assign and_2371_cse = (fsm_output[1:0]==2'b11);
  assign and_2372_cse = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0==4'b1101);
  assign and_nl = (~(act_config_is_zero_first_sva & w_load_lpi_1_dfm_1)) & or_tmp;
  assign nor_nl = ~(w_load_lpi_1_dfm_1 | (~ or_tmp));
  assign mux_16_nl = MUX_s_1_2_2(nor_nl, or_tmp, act_config_is_zero_first_sva);
  assign mux_17_nl = MUX_s_1_2_2(and_nl, mux_16_nl, act_config_is_zero_first_sva_dfm_4);
  assign mux_18_nl = MUX_s_1_2_2(mux_17_nl, or_tmp, ActUnit_RunInst_switch_lp_equal_tmp_3);
  assign Silu_for_y_and_2_cse = ActUnitRun_wen & mux_18_nl & is_start_sva & ActUnit_RunInst_switch_lp_equal_tmp_7;
  assign Silu_for_else_or_7_itm = Silu_for_else_else_else_and_14_ssc_1 | Silu_for_else_else_else_and_15_ssc_1;
  assign Silu_for_else_or_6_itm = Silu_for_else_else_else_and_12_ssc_1 | Silu_for_else_else_else_and_13_ssc_1;
  assign Silu_for_else_or_5_itm = Silu_for_else_else_else_and_10_ssc_1 | Silu_for_else_else_else_and_11_ssc_1;
  assign Silu_for_else_or_4_itm = Silu_for_else_else_else_and_8_ssc_1 | Silu_for_else_else_else_and_9_ssc_1;
  assign Silu_for_else_or_3_itm = Silu_for_else_else_else_and_6_ssc_1 | Silu_for_else_else_else_and_7_ssc_1;
  assign Silu_for_else_or_2_itm = Silu_for_else_else_else_and_4_ssc_1 | Silu_for_else_else_else_and_5_ssc_1;
  assign Silu_for_else_or_1_itm = Silu_for_else_else_else_and_2_ssc_1 | Silu_for_else_else_else_and_3_ssc_1;
  assign Silu_for_else_or_itm = Silu_for_else_else_else_and_ssc_1 | Silu_for_else_else_else_and_1_ssc_1;
  assign nor_1553_cse = ~((ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1:0]!=2'b00));
  assign ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_31_3 = MUX_s_1_64_2(act_regs_data_0_0_sva_dfm_2_31,
      act_regs_data_0_1_sva_dfm_2_31, act_regs_data_0_2_sva_dfm_2_31, act_regs_data_0_3_sva_dfm_2_31,
      act_regs_data_0_4_sva_dfm_2_31, act_regs_data_0_5_sva_dfm_2_31, act_regs_data_0_6_sva_dfm_2_31,
      act_regs_data_0_7_sva_dfm_2_31, act_regs_data_0_8_sva_dfm_2_31, act_regs_data_0_9_sva_dfm_2_31,
      act_regs_data_0_10_sva_dfm_2_31, act_regs_data_0_11_sva_dfm_2_31, act_regs_data_0_12_sva_dfm_2_31,
      act_regs_data_0_13_sva_dfm_2_31, act_regs_data_0_14_sva_dfm_2_31, act_regs_data_0_15_sva_dfm_2_31,
      act_regs_data_1_0_sva_dfm_2_31, act_regs_data_1_1_sva_dfm_2_31, act_regs_data_1_2_sva_dfm_2_31,
      act_regs_data_1_3_sva_dfm_2_31, act_regs_data_1_4_sva_dfm_2_31, act_regs_data_1_5_sva_dfm_2_31,
      act_regs_data_1_6_sva_dfm_2_31, act_regs_data_1_7_sva_dfm_2_31, act_regs_data_1_8_sva_dfm_2_31,
      act_regs_data_1_9_sva_dfm_2_31, act_regs_data_1_10_sva_dfm_2_31, act_regs_data_1_11_sva_dfm_2_31,
      act_regs_data_1_12_sva_dfm_2_31, act_regs_data_1_13_sva_dfm_2_31, act_regs_data_1_14_sva_dfm_2_31,
      act_regs_data_1_15_sva_dfm_2_31, act_regs_data_2_0_sva_dfm_2_31, act_regs_data_2_1_sva_dfm_2_31,
      act_regs_data_2_2_sva_dfm_2_31, act_regs_data_2_3_sva_dfm_2_31, act_regs_data_2_4_sva_dfm_2_31,
      act_regs_data_2_5_sva_dfm_2_31, act_regs_data_2_6_sva_dfm_2_31, act_regs_data_2_7_sva_dfm_2_31,
      act_regs_data_2_8_sva_dfm_2_31, act_regs_data_2_9_sva_dfm_2_31, act_regs_data_2_10_sva_dfm_2_31,
      act_regs_data_2_11_sva_dfm_2_31, act_regs_data_2_12_sva_dfm_2_31, act_regs_data_2_13_sva_dfm_2_31,
      act_regs_data_2_14_sva_dfm_2_31, act_regs_data_2_15_sva_dfm_2_31, act_regs_data_3_0_sva_dfm_2_31,
      act_regs_data_3_1_sva_dfm_2_31, act_regs_data_3_2_sva_dfm_2_31, act_regs_data_3_3_sva_dfm_2_31,
      act_regs_data_3_4_sva_dfm_2_31, act_regs_data_3_5_sva_dfm_2_31, act_regs_data_3_6_sva_dfm_2_31,
      act_regs_data_3_7_sva_dfm_2_31, act_regs_data_3_8_sva_dfm_2_31, act_regs_data_3_9_sva_dfm_2_31,
      act_regs_data_3_10_sva_dfm_2_31, act_regs_data_3_11_sva_dfm_2_31, act_regs_data_3_12_sva_dfm_2_31,
      act_regs_data_3_13_sva_dfm_2_31, act_regs_data_3_14_sva_dfm_2_31, act_regs_data_3_15_sva_dfm_2_31,
      {nvhls_get_slc_2U_NVUINT8_return_2_sva , ActUnit_PushOutput_if_for_i_4_0_sva_3_0});
  assign ActUnit_PushOutput_if_output_port_reg_data_data_and_22_cse = ActUnitRun_wen
      & ((~(or_dcpl_830 | and_dcpl_1090)) | and_dcpl_1244 | and_dcpl_1236);
  assign ActUnit_PushOutput_if_output_port_reg_data_data_and_25_cse = ActUnitRun_wen
      & ((~(or_dcpl_833 | and_dcpl_1090)) | and_dcpl_1244 | and_dcpl_1236);
  assign ActUnit_PushOutput_if_output_port_reg_data_data_and_28_cse = ActUnitRun_wen
      & ((~(or_dcpl_837 | and_dcpl_1090)) | and_dcpl_1244 | and_dcpl_1236);
  assign ActUnit_PushOutput_if_output_port_reg_data_data_and_31_cse = ActUnitRun_wen
      & ((~(or_dcpl_839 | and_dcpl_1090)) | and_dcpl_1244 | and_dcpl_1236);
  assign ActUnit_PushOutput_if_output_port_reg_data_data_and_33_cse = ActUnitRun_wen
      & ((~(or_dcpl_840 | and_dcpl_1090)) | and_dcpl_1244 | and_dcpl_1236);
  assign ActUnit_PushOutput_if_output_port_reg_data_data_and_36_cse = ActUnitRun_wen
      & ((~(or_dcpl_841 | and_dcpl_1090)) | and_dcpl_1244 | and_dcpl_1236);
  assign ActUnit_PushOutput_if_output_port_reg_data_data_and_38_cse = ActUnitRun_wen
      & ((~(or_dcpl_842 | and_dcpl_1090)) | and_dcpl_1244 | and_dcpl_1236);
  assign ActUnit_PushOutput_if_output_port_reg_data_data_and_40_cse = ActUnitRun_wen
      & ((~(or_dcpl_843 | and_dcpl_1090)) | and_dcpl_1244 | and_dcpl_1236);
  assign act_regs_data_and_1186_cse = while_nand_64_ssc_1 & (~ and_dcpl_1246);
  assign act_regs_data_and_1187_cse = ActUnit_RunInst_switch_lp_and_704_ssc_1 & (~
      and_dcpl_1246);
  assign act_regs_data_and_1188_cse = ActUnit_RunInst_switch_lp_and_65_ssc_1 & (~
      and_dcpl_1246);
  assign act_regs_data_and_1189_cse = ActUnit_RunInst_switch_lp_and_67_ssc_1 & (~
      and_dcpl_1246);
  assign act_regs_data_and_1190_cse = ActUnit_RunInst_switch_lp_and_69_ssc_1 & (~
      and_dcpl_1246);
  assign act_regs_data_and_1191_cse = ActUnit_RunInst_switch_lp_and_71_ssc_1 & (~
      and_dcpl_1246);
  assign act_regs_data_and_1192_cse = ActUnit_RunInst_switch_lp_and_73_ssc_1 & (~
      and_dcpl_1246);
  assign nand_542_cse = ~((fsm_output[2:1]==2'b11));
  assign or_1905_cse = (z_out[4]) | (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]) |
      (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign and_2391_nl = nand_542_cse & or_tmp_873;
  assign mux_770_nl = MUX_s_1_2_2((fsm_output[0]), or_tmp_873, or_3395_cse);
  assign mux_771_cse = MUX_s_1_2_2(and_2391_nl, mux_770_nl, fsm_output[3]);
  assign nand_543_cse = ~((fsm_output[0]) & or_tmp_873);
  assign nor_1554_cse = ~((fsm_output[3:1]!=3'b010) | nand_543_cse);
  assign mux_772_nl = MUX_s_1_2_2(mux_771_cse, nor_1554_cse, or_1905_cse);
  assign and_1935_cse = mux_772_nl & ActUnitRun_wen;
  assign or_1913_cse = (z_out[4]) | (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]) |
      (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_775_nl = MUX_s_1_2_2(mux_771_cse, nor_1554_cse, or_1913_cse);
  assign and_1937_cse = mux_775_nl & ActUnitRun_wen;
  assign or_1921_cse = (z_out[4]) | (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]) |
      (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_778_nl = MUX_s_1_2_2(mux_771_cse, nor_1554_cse, or_1921_cse);
  assign and_1939_cse = mux_778_nl & ActUnitRun_wen;
  assign or_1929_cse = (z_out[4]) | (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]) |
      (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_781_nl = MUX_s_1_2_2(mux_771_cse, nor_1554_cse, or_1929_cse);
  assign and_1941_cse = mux_781_nl & ActUnitRun_wen;
  assign or_1937_cse = (z_out[4]) | (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]) |
      (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_784_nl = MUX_s_1_2_2(mux_771_cse, nor_1554_cse, or_1937_cse);
  assign and_1943_cse = mux_784_nl & ActUnitRun_wen;
  assign or_1945_cse = (z_out[4]) | (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]) |
      (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_787_nl = MUX_s_1_2_2(mux_771_cse, nor_1554_cse, or_1945_cse);
  assign and_1945_cse = mux_787_nl & ActUnitRun_wen;
  assign or_1953_cse = (z_out[4]) | (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]) |
      (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_790_nl = MUX_s_1_2_2(mux_771_cse, nor_1554_cse, or_1953_cse);
  assign and_1947_cse = mux_790_nl & ActUnitRun_wen;
  assign or_1961_cse = (z_out[4]) | (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]) |
      (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_793_nl = MUX_s_1_2_2(mux_771_cse, nor_1554_cse, or_1961_cse);
  assign and_1949_cse = mux_793_nl & ActUnitRun_wen;
  assign or_1969_cse = (z_out[4]) | (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]) |
      (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]);
  assign mux_796_nl = MUX_s_1_2_2(or_tmp_938, (~ mux_771_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_797_nl = MUX_s_1_2_2(mux_796_nl, or_tmp_938, or_1969_cse);
  assign and_1951_cse = (~ mux_797_nl) & ActUnitRun_wen;
  assign or_1977_cse = (z_out[4]) | (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]) |
      (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]);
  assign mux_800_nl = MUX_s_1_2_2(or_tmp_938, (~ mux_771_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_801_nl = MUX_s_1_2_2(mux_800_nl, or_tmp_938, or_1977_cse);
  assign and_1953_cse = (~ mux_801_nl) & ActUnitRun_wen;
  assign and_2412_cse = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]) & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign or_1985_cse = (z_out[4]) | (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]) |
      (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]);
  assign mux_804_nl = MUX_s_1_2_2(or_tmp_938, (~ mux_771_cse), and_2412_cse);
  assign mux_805_nl = MUX_s_1_2_2(mux_804_nl, or_tmp_938, or_1985_cse);
  assign and_1955_cse = (~ mux_805_nl) & ActUnitRun_wen;
  assign or_1993_cse = (z_out[4]) | (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]) |
      (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]);
  assign mux_808_nl = MUX_s_1_2_2(or_tmp_938, (~ mux_771_cse), and_2412_cse);
  assign mux_809_nl = MUX_s_1_2_2(mux_808_nl, or_tmp_938, or_1993_cse);
  assign and_1957_cse = (~ mux_809_nl) & ActUnitRun_wen;
  assign or_2001_cse = (z_out[4]) | (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]) |
      (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]);
  assign mux_812_nl = MUX_s_1_2_2(or_tmp_938, (~ mux_771_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_813_nl = MUX_s_1_2_2(mux_812_nl, or_tmp_938, or_2001_cse);
  assign and_1959_cse = (~ mux_813_nl) & ActUnitRun_wen;
  assign or_2009_cse = (z_out[4]) | (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]) |
      (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]);
  assign mux_816_nl = MUX_s_1_2_2(or_tmp_938, (~ mux_771_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_817_nl = MUX_s_1_2_2(mux_816_nl, or_tmp_938, or_2009_cse);
  assign and_1961_cse = (~ mux_817_nl) & ActUnitRun_wen;
  assign or_2017_cse = (z_out[4]) | (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]) |
      (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]);
  assign mux_820_nl = MUX_s_1_2_2(or_tmp_938, (~ mux_771_cse), and_2412_cse);
  assign mux_821_nl = MUX_s_1_2_2(mux_820_nl, or_tmp_938, or_2017_cse);
  assign and_1963_cse = (~ mux_821_nl) & ActUnitRun_wen;
  assign or_2025_cse = (z_out[4]) | (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]) |
      (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]);
  assign mux_824_nl = MUX_s_1_2_2(or_tmp_938, (~ mux_771_cse), and_2412_cse);
  assign mux_825_nl = MUX_s_1_2_2(mux_824_nl, or_tmp_938, or_2025_cse);
  assign and_1965_cse = (~ mux_825_nl) & ActUnitRun_wen;
  assign act_regs_data_and_1298_cse = while_nand_80_ssc_1 & (~ and_dcpl_1246);
  assign act_regs_data_and_1299_cse = ActUnit_RunInst_switch_lp_and_737_ssc_1 & (~
      and_dcpl_1246);
  assign act_regs_data_and_1300_cse = ActUnit_RunInst_switch_lp_and_225_ssc_1 & (~
      and_dcpl_1246);
  assign act_regs_data_and_1301_cse = ActUnit_RunInst_switch_lp_and_227_ssc_1 & (~
      and_dcpl_1246);
  assign act_regs_data_and_1302_cse = ActUnit_RunInst_switch_lp_and_229_ssc_1 & (~
      and_dcpl_1246);
  assign act_regs_data_and_1303_cse = ActUnit_RunInst_switch_lp_and_231_ssc_1 & (~
      and_dcpl_1246);
  assign act_regs_data_and_1304_cse = ActUnit_RunInst_switch_lp_and_233_ssc_1 & (~
      and_dcpl_1246);
  assign or_2033_cse = (z_out[4]) | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign and_2427_nl = nand_542_cse & nand_tmp_41;
  assign mux_826_nl = MUX_s_1_2_2((fsm_output[0]), nand_tmp_41, or_3395_cse);
  assign mux_827_cse = MUX_s_1_2_2(and_2427_nl, mux_826_nl, fsm_output[3]);
  assign nand_583_cse = ~((fsm_output[0]) & nand_tmp_41);
  assign nor_1562_cse = ~((fsm_output[3:1]!=3'b010) | nand_583_cse);
  assign mux_828_nl = MUX_s_1_2_2(mux_827_cse, nor_1562_cse, or_2033_cse);
  assign and_1967_cse = mux_828_nl & ActUnitRun_wen;
  assign or_2040_cse = (z_out[4]) | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]))
      | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_831_nl = MUX_s_1_2_2(mux_827_cse, nor_1562_cse, or_2040_cse);
  assign and_1969_cse = mux_831_nl & ActUnitRun_wen;
  assign or_2047_cse = (z_out[4]) | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_834_nl = MUX_s_1_2_2(mux_827_cse, nor_1562_cse, or_2047_cse);
  assign and_1971_cse = mux_834_nl & ActUnitRun_wen;
  assign or_2054_cse = (z_out[4]) | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]))
      | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_837_nl = MUX_s_1_2_2(mux_827_cse, nor_1562_cse, or_2054_cse);
  assign and_1973_cse = mux_837_nl & ActUnitRun_wen;
  assign or_2061_cse = (z_out[4]) | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_840_nl = MUX_s_1_2_2(mux_827_cse, nor_1562_cse, or_2061_cse);
  assign and_1975_cse = mux_840_nl & ActUnitRun_wen;
  assign or_2068_cse = (z_out[4]) | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]))
      | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_843_nl = MUX_s_1_2_2(mux_827_cse, nor_1562_cse, or_2068_cse);
  assign and_1977_cse = mux_843_nl & ActUnitRun_wen;
  assign or_2075_cse = (z_out[4]) | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_846_nl = MUX_s_1_2_2(mux_827_cse, nor_1562_cse, or_2075_cse);
  assign and_1979_cse = mux_846_nl & ActUnitRun_wen;
  assign or_2082_cse = (z_out[4]) | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]))
      | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_849_nl = MUX_s_1_2_2(mux_827_cse, nor_1562_cse, or_2082_cse);
  assign and_1981_cse = mux_849_nl & ActUnitRun_wen;
  assign or_2089_cse = (z_out[4]) | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]);
  assign mux_852_nl = MUX_s_1_2_2(or_tmp_1057, (~ mux_827_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_853_nl = MUX_s_1_2_2(mux_852_nl, or_tmp_1057, or_2089_cse);
  assign and_1983_cse = (~ mux_853_nl) & ActUnitRun_wen;
  assign or_2096_cse = (z_out[4]) | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]))
      | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]);
  assign mux_856_nl = MUX_s_1_2_2(or_tmp_1057, (~ mux_827_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_857_nl = MUX_s_1_2_2(mux_856_nl, or_tmp_1057, or_2096_cse);
  assign and_1985_cse = (~ mux_857_nl) & ActUnitRun_wen;
  assign or_2103_cse = (z_out[4]) | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]);
  assign mux_860_nl = MUX_s_1_2_2(or_tmp_1057, (~ mux_827_cse), and_2412_cse);
  assign mux_861_nl = MUX_s_1_2_2(mux_860_nl, or_tmp_1057, or_2103_cse);
  assign and_1987_cse = (~ mux_861_nl) & ActUnitRun_wen;
  assign or_2110_cse = (z_out[4]) | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]))
      | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2])
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]);
  assign mux_864_nl = MUX_s_1_2_2(or_tmp_1057, (~ mux_827_cse), and_2412_cse);
  assign mux_865_nl = MUX_s_1_2_2(mux_864_nl, or_tmp_1057, or_2110_cse);
  assign and_1989_cse = (~ mux_865_nl) & ActUnitRun_wen;
  assign or_2117_cse = (z_out[4]) | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]);
  assign mux_868_nl = MUX_s_1_2_2(or_tmp_1057, (~ mux_827_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_869_nl = MUX_s_1_2_2(mux_868_nl, or_tmp_1057, or_2117_cse);
  assign and_1991_cse = (~ mux_869_nl) & ActUnitRun_wen;
  assign or_2124_cse = (z_out[4]) | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]))
      | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]);
  assign mux_872_nl = MUX_s_1_2_2(or_tmp_1057, (~ mux_827_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_873_nl = MUX_s_1_2_2(mux_872_nl, or_tmp_1057, or_2124_cse);
  assign and_1993_cse = (~ mux_873_nl) & ActUnitRun_wen;
  assign or_2131_cse = (z_out[4]) | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]);
  assign mux_876_nl = MUX_s_1_2_2(or_tmp_1057, (~ mux_827_cse), and_2412_cse);
  assign mux_877_nl = MUX_s_1_2_2(mux_876_nl, or_tmp_1057, or_2131_cse);
  assign and_1995_cse = (~ mux_877_nl) & ActUnitRun_wen;
  assign or_2138_cse = (z_out[4]) | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]))
      | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]))
      | (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]);
  assign mux_880_nl = MUX_s_1_2_2(or_tmp_1057, (~ mux_827_cse), and_2412_cse);
  assign mux_881_nl = MUX_s_1_2_2(mux_880_nl, or_tmp_1057, or_2138_cse);
  assign and_1997_cse = (~ mux_881_nl) & ActUnitRun_wen;
  assign act_regs_data_and_1410_cse = while_nand_96_ssc_1 & (~ and_dcpl_1246);
  assign act_regs_data_and_1411_cse = ActUnit_RunInst_switch_lp_and_769_ssc_1 & (~
      and_dcpl_1246);
  assign act_regs_data_and_1412_cse = ActUnit_RunInst_switch_lp_and_385_ssc_1 & (~
      and_dcpl_1246);
  assign act_regs_data_and_1413_cse = ActUnit_RunInst_switch_lp_and_387_ssc_1 & (~
      and_dcpl_1246);
  assign act_regs_data_and_1414_cse = ActUnit_RunInst_switch_lp_and_389_ssc_1 & (~
      and_dcpl_1246);
  assign act_regs_data_and_1415_cse = ActUnit_RunInst_switch_lp_and_391_ssc_1 & (~
      and_dcpl_1246);
  assign act_regs_data_and_1416_cse = ActUnit_RunInst_switch_lp_and_393_ssc_1 & (~
      and_dcpl_1246);
  assign or_2145_cse = (z_out[4]) | (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]) |
      (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2])
      | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[1])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign and_2463_nl = nand_542_cse & or_tmp_1113;
  assign mux_882_nl = MUX_s_1_2_2((fsm_output[0]), or_tmp_1113, or_3395_cse);
  assign mux_883_cse = MUX_s_1_2_2(and_2463_nl, mux_882_nl, fsm_output[3]);
  assign nand_623_cse = ~((fsm_output[0]) & or_tmp_1113);
  assign nor_1570_cse = ~((fsm_output[3:1]!=3'b010) | nand_623_cse);
  assign mux_884_nl = MUX_s_1_2_2(mux_883_cse, nor_1570_cse, or_2145_cse);
  assign and_1999_cse = mux_884_nl & ActUnitRun_wen;
  assign or_2153_cse = (z_out[4]) | (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]) |
      (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2])
      | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[1])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_887_nl = MUX_s_1_2_2(mux_883_cse, nor_1570_cse, or_2153_cse);
  assign and_2001_cse = mux_887_nl & ActUnitRun_wen;
  assign or_2161_cse = (z_out[4]) | (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]) |
      (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2])
      | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[1])) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_890_nl = MUX_s_1_2_2(mux_883_cse, nor_1570_cse, or_2161_cse);
  assign and_2003_cse = mux_890_nl & ActUnitRun_wen;
  assign or_2169_cse = (z_out[4]) | (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]) |
      (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2])
      | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[1])) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_893_nl = MUX_s_1_2_2(mux_883_cse, nor_1570_cse, or_2169_cse);
  assign and_2005_cse = mux_893_nl & ActUnitRun_wen;
  assign or_2177_cse = (z_out[4]) | (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]) |
      (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]))
      | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[1])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_896_nl = MUX_s_1_2_2(mux_883_cse, nor_1570_cse, or_2177_cse);
  assign and_2007_cse = mux_896_nl & ActUnitRun_wen;
  assign or_2185_cse = (z_out[4]) | (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]) |
      (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]))
      | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[1])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_899_nl = MUX_s_1_2_2(mux_883_cse, nor_1570_cse, or_2185_cse);
  assign and_2009_cse = mux_899_nl & ActUnitRun_wen;
  assign or_2193_cse = (z_out[4]) | (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]) |
      (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]))
      | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[1])) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_902_nl = MUX_s_1_2_2(mux_883_cse, nor_1570_cse, or_2193_cse);
  assign and_2011_cse = mux_902_nl & ActUnitRun_wen;
  assign or_2201_cse = (z_out[4]) | (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]) |
      (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]))
      | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[1])) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_905_nl = MUX_s_1_2_2(mux_883_cse, nor_1570_cse, or_2201_cse);
  assign and_2013_cse = mux_905_nl & ActUnitRun_wen;
  assign or_2209_cse = (z_out[4]) | (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]) |
      (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2])
      | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[1])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]);
  assign mux_908_nl = MUX_s_1_2_2(or_tmp_1178, (~ mux_883_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_909_nl = MUX_s_1_2_2(mux_908_nl, or_tmp_1178, or_2209_cse);
  assign and_2015_cse = (~ mux_909_nl) & ActUnitRun_wen;
  assign or_2217_cse = (z_out[4]) | (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]) |
      (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2])
      | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[1])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]);
  assign mux_912_nl = MUX_s_1_2_2(or_tmp_1178, (~ mux_883_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_913_nl = MUX_s_1_2_2(mux_912_nl, or_tmp_1178, or_2217_cse);
  assign and_2017_cse = (~ mux_913_nl) & ActUnitRun_wen;
  assign and_2484_cse = (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]) & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign or_2225_cse = (z_out[4]) | (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]) |
      (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign mux_916_nl = MUX_s_1_2_2(or_tmp_1178, (~ mux_883_cse), and_2484_cse);
  assign mux_917_nl = MUX_s_1_2_2(mux_916_nl, or_tmp_1178, or_2225_cse);
  assign and_2019_cse = (~ mux_917_nl) & ActUnitRun_wen;
  assign or_2233_cse = (z_out[4]) | (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]) |
      (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign mux_920_nl = MUX_s_1_2_2(or_tmp_1178, (~ mux_883_cse), and_2484_cse);
  assign mux_921_nl = MUX_s_1_2_2(mux_920_nl, or_tmp_1178, or_2233_cse);
  assign and_2021_cse = (~ mux_921_nl) & ActUnitRun_wen;
  assign or_2241_cse = (z_out[4]) | (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]) |
      (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]))
      | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[1])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]);
  assign mux_924_nl = MUX_s_1_2_2(or_tmp_1178, (~ mux_883_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_925_nl = MUX_s_1_2_2(mux_924_nl, or_tmp_1178, or_2241_cse);
  assign and_2023_cse = (~ mux_925_nl) & ActUnitRun_wen;
  assign or_2249_cse = (z_out[4]) | (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]) |
      (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]))
      | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[1])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]);
  assign mux_928_nl = MUX_s_1_2_2(or_tmp_1178, (~ mux_883_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_929_nl = MUX_s_1_2_2(mux_928_nl, or_tmp_1178, or_2249_cse);
  assign and_2025_cse = (~ mux_929_nl) & ActUnitRun_wen;
  assign and_2494_cse = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]) & (nvhls_get_slc_2U_NVUINT8_return_3_sva[1])
      & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]) & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign or_2257_cse = (z_out[4]) | (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]) |
      (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]);
  assign mux_932_nl = MUX_s_1_2_2(or_tmp_1178, (~ mux_883_cse), and_2494_cse);
  assign mux_933_nl = MUX_s_1_2_2(mux_932_nl, or_tmp_1178, or_2257_cse);
  assign and_2027_cse = (~ mux_933_nl) & ActUnitRun_wen;
  assign and_2497_cse = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]) & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2])
      & (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]) & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign or_2265_cse = (z_out[4]) | (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]);
  assign mux_936_nl = MUX_s_1_2_2(or_tmp_1178, (~ mux_883_cse), and_2497_cse);
  assign mux_937_nl = MUX_s_1_2_2(mux_936_nl, or_tmp_1178, or_2265_cse);
  assign and_2029_cse = (~ mux_937_nl) & ActUnitRun_wen;
  assign act_regs_data_and_1522_cse = while_nand_112_ssc_1 & (~ and_dcpl_1246);
  assign act_regs_data_and_1523_cse = ActUnit_RunInst_switch_lp_and_801_ssc_1 & (~
      and_dcpl_1246);
  assign act_regs_data_and_1524_cse = ActUnit_RunInst_switch_lp_and_545_ssc_1 & (~
      and_dcpl_1246);
  assign act_regs_data_and_1525_cse = ActUnit_RunInst_switch_lp_and_547_ssc_1 & (~
      and_dcpl_1246);
  assign act_regs_data_and_1526_cse = ActUnit_RunInst_switch_lp_and_549_ssc_1 & (~
      and_dcpl_1246);
  assign act_regs_data_and_1527_cse = ActUnit_RunInst_switch_lp_and_551_ssc_1 & (~
      and_dcpl_1246);
  assign act_regs_data_and_1528_cse = ActUnit_RunInst_switch_lp_and_553_ssc_1 & (~
      and_dcpl_1246);
  assign or_2273_cse = (z_out[4]) | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2])
      | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[1])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign and_2499_nl = nand_542_cse & nand_tmp_73;
  assign mux_938_nl = MUX_s_1_2_2((fsm_output[0]), nand_tmp_73, or_3395_cse);
  assign mux_939_cse = MUX_s_1_2_2(and_2499_nl, mux_938_nl, fsm_output[3]);
  assign nand_663_cse = ~((fsm_output[0]) & nand_tmp_73);
  assign nor_1578_cse = ~((fsm_output[3:1]!=3'b010) | nand_663_cse);
  assign mux_940_nl = MUX_s_1_2_2(mux_939_cse, nor_1578_cse, or_2273_cse);
  assign and_2031_cse = mux_940_nl & ActUnitRun_wen;
  assign or_2280_cse = (z_out[4]) | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]))
      | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2])
      | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[1])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_943_nl = MUX_s_1_2_2(mux_939_cse, nor_1578_cse, or_2280_cse);
  assign and_2033_cse = mux_943_nl & ActUnitRun_wen;
  assign or_2287_cse = (z_out[4]) | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2])
      | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[1])) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_946_nl = MUX_s_1_2_2(mux_939_cse, nor_1578_cse, or_2287_cse);
  assign and_2035_cse = mux_946_nl & ActUnitRun_wen;
  assign or_2294_cse = (z_out[4]) | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]))
      | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2])
      | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[1])) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_949_nl = MUX_s_1_2_2(mux_939_cse, nor_1578_cse, or_2294_cse);
  assign and_2037_cse = mux_949_nl & ActUnitRun_wen;
  assign or_2301_cse = (z_out[4]) | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]))
      | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[1])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_952_nl = MUX_s_1_2_2(mux_939_cse, nor_1578_cse, or_2301_cse);
  assign and_2039_cse = mux_952_nl & ActUnitRun_wen;
  assign or_2308_cse = (z_out[4]) | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]))
      | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]))
      | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[1])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_955_nl = MUX_s_1_2_2(mux_939_cse, nor_1578_cse, or_2308_cse);
  assign and_2041_cse = mux_955_nl & ActUnitRun_wen;
  assign or_2315_cse = (z_out[4]) | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]))
      | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[1])) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_958_nl = MUX_s_1_2_2(mux_939_cse, nor_1578_cse, or_2315_cse);
  assign and_2043_cse = mux_958_nl & ActUnitRun_wen;
  assign nand_685_cse = ~((~ (z_out[4])) & (nvhls_get_slc_2U_NVUINT8_return_3_sva[0])
      & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]) & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2])
      & (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]) & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1])
      & (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3])));
  assign mux_961_nl = MUX_s_1_2_2(mux_939_cse, nor_1578_cse, nand_685_cse);
  assign and_2045_cse = mux_961_nl & ActUnitRun_wen;
  assign or_2329_cse = (z_out[4]) | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2])
      | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[1])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]);
  assign mux_964_nl = MUX_s_1_2_2(or_tmp_1297, (~ mux_939_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_965_nl = MUX_s_1_2_2(mux_964_nl, or_tmp_1297, or_2329_cse);
  assign and_2047_cse = (~ mux_965_nl) & ActUnitRun_wen;
  assign or_2336_cse = (z_out[4]) | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]))
      | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2])
      | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[1])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]);
  assign mux_968_nl = MUX_s_1_2_2(or_tmp_1297, (~ mux_939_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_969_nl = MUX_s_1_2_2(mux_968_nl, or_tmp_1297, or_2336_cse);
  assign and_2049_cse = (~ mux_969_nl) & ActUnitRun_wen;
  assign or_2343_cse = (z_out[4]) | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign mux_972_nl = MUX_s_1_2_2(or_tmp_1297, (~ mux_939_cse), and_2484_cse);
  assign mux_973_nl = MUX_s_1_2_2(mux_972_nl, or_tmp_1297, or_2343_cse);
  assign and_2051_cse = (~ mux_973_nl) & ActUnitRun_wen;
  assign or_2350_cse = (z_out[4]) | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]))
      | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]);
  assign mux_976_nl = MUX_s_1_2_2(or_tmp_1297, (~ mux_939_cse), and_2484_cse);
  assign mux_977_nl = MUX_s_1_2_2(mux_976_nl, or_tmp_1297, or_2350_cse);
  assign and_2053_cse = (~ mux_977_nl) & ActUnitRun_wen;
  assign or_2357_cse = (z_out[4]) | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]))
      | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[1])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]);
  assign mux_980_nl = MUX_s_1_2_2(or_tmp_1297, (~ mux_939_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_981_nl = MUX_s_1_2_2(mux_980_nl, or_tmp_1297, or_2357_cse);
  assign and_2055_cse = (~ mux_981_nl) & ActUnitRun_wen;
  assign or_2364_cse = (z_out[4]) | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]))
      | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]))
      | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[1])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]);
  assign mux_984_nl = MUX_s_1_2_2(or_tmp_1297, (~ mux_939_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_985_nl = MUX_s_1_2_2(mux_984_nl, or_tmp_1297, or_2364_cse);
  assign and_2057_cse = (~ mux_985_nl) & ActUnitRun_wen;
  assign or_2371_cse = (z_out[4]) | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]))
      | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]);
  assign mux_988_nl = MUX_s_1_2_2(or_tmp_1297, (~ mux_939_cse), and_2494_cse);
  assign mux_989_nl = MUX_s_1_2_2(mux_988_nl, or_tmp_1297, or_2371_cse);
  assign and_2059_cse = (~ mux_989_nl) & ActUnitRun_wen;
  assign and_2533_cse = (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]) & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])
      & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2]) & (nvhls_get_slc_2U_NVUINT8_return_3_sva[1])
      & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]) & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_992_nl = MUX_s_1_2_2(or_tmp_1297, (~ mux_939_cse), and_2533_cse);
  assign mux_993_nl = MUX_s_1_2_2(mux_992_nl, or_tmp_1297, z_out[4]);
  assign and_2061_cse = (~ mux_993_nl) & ActUnitRun_wen;
  assign and_2535_nl = nand_542_cse & nand_tmp_104;
  assign mux_994_nl = MUX_s_1_2_2((fsm_output[0]), nand_tmp_104, or_3395_cse);
  assign mux_995_cse = MUX_s_1_2_2(and_2535_nl, mux_994_nl, fsm_output[3]);
  assign nand_704_cse = ~((fsm_output[0]) & nand_tmp_104);
  assign nor_1586_cse = ~((fsm_output[3:1]!=3'b010) | nand_704_cse);
  assign and_2571_nl = nand_542_cse & nand_tmp_120;
  assign mux_1051_nl = MUX_s_1_2_2((fsm_output[0]), nand_tmp_120, or_3395_cse);
  assign mux_1052_cse = MUX_s_1_2_2(and_2571_nl, mux_1051_nl, fsm_output[3]);
  assign nand_744_cse = ~((fsm_output[0]) & nand_tmp_120);
  assign nor_1594_cse = ~((fsm_output[3:1]!=3'b010) | nand_744_cse);
  assign and_2607_nl = nand_542_cse & nand_tmp_136;
  assign mux_1122_nl = MUX_s_1_2_2((fsm_output[0]), nand_tmp_136, or_3395_cse);
  assign mux_1123_cse = MUX_s_1_2_2(and_2607_nl, mux_1122_nl, fsm_output[3]);
  assign nand_784_cse = ~((fsm_output[0]) & nand_tmp_136);
  assign nor_1602_cse = ~((fsm_output[3:1]!=3'b010) | nand_784_cse);
  assign and_2643_nl = nand_542_cse & nand_tmp_152;
  assign mux_1179_nl = MUX_s_1_2_2((fsm_output[0]), nand_tmp_152, or_3395_cse);
  assign mux_1180_cse = MUX_s_1_2_2(and_2643_nl, mux_1179_nl, fsm_output[3]);
  assign nand_824_cse = ~((fsm_output[0]) & nand_tmp_152);
  assign nor_1610_cse = ~((fsm_output[3:1]!=3'b010) | nand_824_cse);
  assign and_1648_cse = (act_config_in_InstFetch_return_sva_7_2[5:3]==3'b111);
  assign nor_447_cse = ~((operator_6_false_acc_tmp[6:5]!=2'b00));
  assign ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_mx1
      = MUX_s_1_2_2(rva_in_PopNB_mioi_return_rsc_z_mxwt, ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva,
      is_start_sva);
  assign ActUnit_DecodeAxi_rva_in_reg_rw_sva_mx1 = MUX_s_1_2_2(rva_in_PopNB_mioi_data_rw_rsc_z_mxwt,
      ActUnit_DecodeAxi_rva_in_reg_rw_sva, is_start_sva);
  assign ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0 = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11:8]==4'b1001));
  assign ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_23_4_mx1_tmp_7_0
      = MUX_v_8_2_2((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7:0]), reg_ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_23_4_ftd_12,
      is_start_sva);
  assign act_mem_banks_read_read_data_lpi_1_dfm_1_31_0_mx1 = MUX_v_32_2_2(act_mem_banks_read_for_mux_15_itm,
      act_mem_banks_read_read_data_lpi_1_dfm_1_31_0, act_write_req_valid_lpi_1_dfm_5);
  assign act_mem_banks_read_read_data_lpi_1_dfm_1_63_32_mx1 = MUX_v_32_2_2(act_mem_banks_read_for_mux_14_itm,
      act_mem_banks_read_read_data_lpi_1_dfm_1_63_32, act_write_req_valid_lpi_1_dfm_5);
  assign act_mem_banks_read_read_data_lpi_1_dfm_1_95_64_mx1 = MUX_v_32_2_2(act_mem_banks_read_for_mux_13_itm,
      act_mem_banks_read_read_data_lpi_1_dfm_1_95_64, act_write_req_valid_lpi_1_dfm_5);
  assign act_mem_banks_read_read_data_lpi_1_dfm_1_127_96_mx1 = MUX_v_32_2_2(act_mem_banks_read_for_mux_12_itm,
      act_mem_banks_read_read_data_lpi_1_dfm_1_127_96, act_write_req_valid_lpi_1_dfm_5);
  assign act_mem_banks_read_read_data_lpi_1_dfm_1_159_128_mx1 = MUX_v_32_2_2(act_mem_banks_read_for_mux_11_itm,
      act_mem_banks_read_read_data_lpi_1_dfm_1_159_128, act_write_req_valid_lpi_1_dfm_5);
  assign act_mem_banks_read_read_data_lpi_1_dfm_1_191_160_mx1 = MUX_v_32_2_2(act_mem_banks_read_for_mux_10_itm,
      act_mem_banks_read_read_data_lpi_1_dfm_1_191_160, act_write_req_valid_lpi_1_dfm_5);
  assign act_mem_banks_read_read_data_lpi_1_dfm_1_223_192_mx1 = MUX_v_32_2_2(act_mem_banks_read_for_mux_9_itm,
      act_mem_banks_read_read_data_lpi_1_dfm_1_223_192, act_write_req_valid_lpi_1_dfm_5);
  assign act_mem_banks_read_read_data_lpi_1_dfm_1_255_224_mx1 = MUX_v_32_2_2(act_mem_banks_read_for_mux_8_itm,
      act_mem_banks_read_read_data_lpi_1_dfm_1_255_224, act_write_req_valid_lpi_1_dfm_5);
  assign act_mem_banks_read_read_data_lpi_1_dfm_1_287_256_mx1 = MUX_v_32_2_2(act_mem_banks_read_for_mux_7_itm,
      act_mem_banks_read_read_data_lpi_1_dfm_1_287_256, act_write_req_valid_lpi_1_dfm_5);
  assign act_mem_banks_read_read_data_lpi_1_dfm_1_319_288_mx1 = MUX_v_32_2_2(act_mem_banks_read_for_mux_6_itm,
      act_mem_banks_read_read_data_lpi_1_dfm_1_319_288, act_write_req_valid_lpi_1_dfm_5);
  assign act_mem_banks_read_read_data_lpi_1_dfm_1_351_320_mx1 = MUX_v_32_2_2(act_mem_banks_read_for_mux_5_itm,
      act_mem_banks_read_read_data_lpi_1_dfm_1_351_320, act_write_req_valid_lpi_1_dfm_5);
  assign act_mem_banks_read_read_data_lpi_1_dfm_1_383_352_mx1 = MUX_v_32_2_2(act_mem_banks_read_for_mux_4_itm,
      act_mem_banks_read_read_data_lpi_1_dfm_1_383_352, act_write_req_valid_lpi_1_dfm_5);
  assign act_mem_banks_read_read_data_lpi_1_dfm_1_415_384_mx1 = MUX_v_32_2_2(act_mem_banks_read_for_mux_3_itm,
      act_mem_banks_read_read_data_lpi_1_dfm_1_415_384, act_write_req_valid_lpi_1_dfm_5);
  assign act_mem_banks_read_read_data_lpi_1_dfm_1_447_416_mx1 = MUX_v_32_2_2(act_mem_banks_read_for_mux_2_itm,
      act_mem_banks_read_read_data_lpi_1_dfm_1_447_416, act_write_req_valid_lpi_1_dfm_5);
  assign act_mem_banks_read_read_data_lpi_1_dfm_1_479_448_mx1 = MUX_v_32_2_2(act_mem_banks_read_for_mux_1_itm,
      act_mem_banks_read_read_data_lpi_1_dfm_1_479_448, act_write_req_valid_lpi_1_dfm_5);
  assign act_mem_banks_read_read_data_lpi_1_dfm_1_511_480_mx1 = MUX_v_32_2_2(act_mem_banks_read_for_mux_itm,
      act_mem_banks_read_read_data_lpi_1_dfm_1_511_480, act_write_req_valid_lpi_1_dfm_5);
  assign nl_Gelu_for_1_else_if_acc_itm_mx1w0 = conv_u2s_3_4(Silu_for_1_else_if_Silu_for_else_if_mul_cmp_7_z[47:45])
      + 4'b1111;
  assign Gelu_for_1_else_if_acc_itm_mx1w0 = nl_Gelu_for_1_else_if_acc_itm_mx1w0[3:0];
  assign nl_Gelu_for_2_else_if_acc_itm_mx1w0 = conv_u2s_3_4(Silu_for_1_else_if_Silu_for_else_if_mul_cmp_z[47:45])
      + 4'b1111;
  assign Gelu_for_2_else_if_acc_itm_mx1w0 = nl_Gelu_for_2_else_if_acc_itm_mx1w0[3:0];
  assign nl_Gelu_for_3_else_if_acc_itm_mx1w0 = conv_u2s_3_4(Silu_for_1_else_if_Silu_for_else_if_mul_cmp_6_z[47:45])
      + 4'b1111;
  assign Gelu_for_3_else_if_acc_itm_mx1w0 = nl_Gelu_for_3_else_if_acc_itm_mx1w0[3:0];
  assign nl_Gelu_for_4_else_if_acc_itm_mx1w0 = conv_u2s_3_4(Silu_for_1_else_if_Silu_for_else_if_mul_cmp_5_z[47:45])
      + 4'b1111;
  assign Gelu_for_4_else_if_acc_itm_mx1w0 = nl_Gelu_for_4_else_if_acc_itm_mx1w0[3:0];
  assign nl_Gelu_for_5_else_if_acc_itm_mx1w0 = conv_u2s_3_4(Silu_for_1_else_if_Silu_for_else_if_mul_cmp_4_z[47:45])
      + 4'b1111;
  assign Gelu_for_5_else_if_acc_itm_mx1w0 = nl_Gelu_for_5_else_if_acc_itm_mx1w0[3:0];
  assign nl_Gelu_for_6_else_if_acc_itm_mx1w0 = conv_u2s_3_4(Silu_for_1_else_if_Silu_for_else_if_mul_cmp_3_z[47:45])
      + 4'b1111;
  assign Gelu_for_6_else_if_acc_itm_mx1w0 = nl_Gelu_for_6_else_if_acc_itm_mx1w0[3:0];
  assign nl_Gelu_for_7_else_if_acc_itm_mx1w0 = conv_u2s_3_4(Silu_for_1_else_if_Silu_for_else_if_mul_cmp_2_z[47:45])
      + 4'b1111;
  assign Gelu_for_7_else_if_acc_itm_mx1w0 = nl_Gelu_for_7_else_if_acc_itm_mx1w0[3:0];
  assign nl_Gelu_for_8_else_if_acc_itm_mx1w0 = conv_u2s_3_4(Silu_for_1_else_if_Silu_for_else_if_mul_cmp_1_z[47:45])
      + 4'b1111;
  assign Gelu_for_8_else_if_acc_itm_mx1w0 = nl_Gelu_for_8_else_if_acc_itm_mx1w0[3:0];
  assign operator_32_8_true_AC_TRN_AC_WRAP_1_less_15_tmp = $signed(26'b10000000000000000000000000)
      < $signed(({nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign Silu_for_else_and_1_tmp = Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign Silu_for_else_and_1_m1c_mx1 = MUX_s_1_2_2(Silu_for_else_and_1_m1c, Silu_for_else_and_1_tmp,
      Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
  assign operator_32_8_true_AC_TRN_AC_WRAP_1_less_14_tmp = $signed(26'b10000000000000000000000000)
      < $signed(({nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign Silu_for_else_and_3_tmp = Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign Silu_for_else_and_3_m1c_mx1 = MUX_s_1_2_2(Silu_for_else_and_3_m1c, Silu_for_else_and_3_tmp,
      Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
  assign operator_32_8_true_AC_TRN_AC_WRAP_1_less_13_tmp = $signed(26'b10000000000000000000000000)
      < $signed(({nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign Silu_for_else_and_5_tmp = Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign Silu_for_else_and_5_m1c_mx1 = MUX_s_1_2_2(Silu_for_else_and_5_m1c, Silu_for_else_and_5_tmp,
      Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
  assign operator_32_8_true_AC_TRN_AC_WRAP_1_less_12_tmp = $signed(26'b10000000000000000000000000)
      < $signed(({nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign Silu_for_else_and_7_tmp = Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign Silu_for_else_and_7_m1c_mx1 = MUX_s_1_2_2(Silu_for_else_and_7_m1c, Silu_for_else_and_7_tmp,
      Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
  assign operator_32_8_true_AC_TRN_AC_WRAP_1_less_11_tmp = $signed(26'b10000000000000000000000000)
      < $signed(({nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign Silu_for_else_and_9_tmp = Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign Silu_for_else_and_9_m1c_mx1 = MUX_s_1_2_2(Silu_for_else_and_9_m1c, Silu_for_else_and_9_tmp,
      Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
  assign operator_32_8_true_AC_TRN_AC_WRAP_1_less_10_tmp = $signed(26'b10000000000000000000000000)
      < $signed(({nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign Silu_for_else_and_11_tmp = Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign Silu_for_else_and_11_m1c_mx1 = MUX_s_1_2_2(Silu_for_else_and_11_m1c, Silu_for_else_and_11_tmp,
      Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
  assign operator_32_8_true_AC_TRN_AC_WRAP_1_less_9_tmp = $signed(26'b10000000000000000000000000)
      < $signed(({nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign Silu_for_else_and_13_tmp = Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign Silu_for_else_and_13_m1c_mx1 = MUX_s_1_2_2(Silu_for_else_and_13_m1c, Silu_for_else_and_13_tmp,
      Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
  assign operator_32_8_true_AC_TRN_AC_WRAP_1_less_8_tmp = $signed(26'b10000000000000000000000000)
      < $signed(({nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign Silu_for_else_and_15_tmp = Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign Silu_for_else_and_15_m1c_mx1 = MUX_s_1_2_2(Silu_for_else_and_15_m1c, Silu_for_else_and_15_tmp,
      Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
  assign Gelu_for_else_if_less_15_tmp = $signed(25'b1010000000000000000000000) <
      $signed(({nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign Gelu_for_else_if_less_14_tmp = $signed(25'b1010000000000000000000000) <
      $signed(({nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign Gelu_for_else_if_less_13_tmp = $signed(25'b1010000000000000000000000) <
      $signed(({nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign Gelu_for_else_if_less_12_tmp = $signed(25'b1010000000000000000000000) <
      $signed(({nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign Gelu_for_else_if_less_11_tmp = $signed(25'b1010000000000000000000000) <
      $signed(({nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign Gelu_for_else_if_less_10_tmp = $signed(25'b1010000000000000000000000) <
      $signed(({nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign Gelu_for_else_if_less_9_tmp = $signed(25'b1010000000000000000000000) < $signed(({nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign Gelu_for_else_if_less_8_tmp = $signed(25'b1010000000000000000000000) < $signed(({nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign Silu_for_else_and_17_m1c_mx0w1 = Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign Silu_for_else_and_17_m1c_mx1 = MUX_s_1_2_2(Silu_for_else_and_17_m1c, Silu_for_else_and_17_m1c_mx0w1,
      Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
  assign Silu_for_else_and_19_tmp = Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign Silu_for_else_and_19_m1c_mx1 = MUX_s_1_2_2(Silu_for_else_and_19_m1c, Silu_for_else_and_19_tmp,
      Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
  assign Silu_for_else_and_21_m1c_mx0w1 = Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign Silu_for_else_and_21_m1c_mx1 = MUX_s_1_2_2(Silu_for_else_and_21_m1c, Silu_for_else_and_21_m1c_mx0w1,
      Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
  assign Silu_for_else_and_23_m1c_mx0w1 = Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign Silu_for_else_and_23_m1c_mx1 = MUX_s_1_2_2(Silu_for_else_and_23_m1c, Silu_for_else_and_23_m1c_mx0w1,
      Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
  assign Silu_for_else_and_25_m1c_mx0w1 = Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign Silu_for_else_and_25_m1c_mx1 = MUX_s_1_2_2(Silu_for_else_and_25_m1c, Silu_for_else_and_25_m1c_mx0w1,
      Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
  assign Silu_for_else_and_27_m1c_mx0w1 = Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign Silu_for_else_and_27_m1c_mx1 = MUX_s_1_2_2(Silu_for_else_and_27_m1c, Silu_for_else_and_27_m1c_mx0w1,
      Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
  assign Silu_for_else_and_29_m1c_mx0w1 = Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign Silu_for_else_and_29_m1c_mx1 = MUX_s_1_2_2(Silu_for_else_and_29_m1c, Silu_for_else_and_29_m1c_mx0w1,
      Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
  assign Silu_for_else_and_31_m1c_mx0w1 = Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign Silu_for_else_and_31_m1c_mx1 = MUX_s_1_2_2(Silu_for_else_and_31_m1c, Silu_for_else_and_31_m1c_mx0w1,
      Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
  assign Gelu_for_else_and_1_tmp = Gelu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
      & Gelu_for_1_else_slc_32_svs;
  assign Gelu_for_else_and_1_m1c_mx1 = MUX_s_1_2_2(Gelu_for_else_and_1_m1c, Gelu_for_else_and_1_tmp,
      Gelu_for_1_slc_32_1_svs);
  assign Gelu_for_else_and_3_tmp = Gelu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
      & Gelu_for_2_else_slc_32_svs;
  assign Gelu_for_else_and_3_m1c_mx1 = MUX_s_1_2_2(Gelu_for_else_and_3_m1c, Gelu_for_else_and_3_tmp,
      Gelu_for_2_slc_32_1_svs);
  assign Gelu_for_else_and_5_tmp = Gelu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
      & Gelu_for_3_else_slc_32_svs;
  assign Gelu_for_else_and_5_m1c_mx1 = MUX_s_1_2_2(Gelu_for_else_and_5_m1c, Gelu_for_else_and_5_tmp,
      Gelu_for_3_slc_32_1_svs);
  assign Gelu_for_else_and_7_tmp = Gelu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
      & Gelu_for_4_else_slc_32_svs;
  assign Gelu_for_else_and_7_m1c_mx1 = MUX_s_1_2_2(Gelu_for_else_and_7_m1c, Gelu_for_else_and_7_tmp,
      Gelu_for_4_slc_32_1_svs);
  assign Gelu_for_else_and_9_tmp = Gelu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
      & Gelu_for_5_else_slc_32_svs;
  assign Gelu_for_else_and_9_m1c_mx1 = MUX_s_1_2_2(Gelu_for_else_and_9_m1c, Gelu_for_else_and_9_tmp,
      Gelu_for_5_slc_32_1_svs);
  assign Gelu_for_else_and_11_tmp = Gelu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
      & Gelu_for_6_else_slc_32_svs;
  assign Gelu_for_else_and_11_m1c_mx1 = MUX_s_1_2_2(Gelu_for_else_and_11_m1c, Gelu_for_else_and_11_tmp,
      Gelu_for_6_slc_32_1_svs);
  assign Gelu_for_else_and_13_tmp = Gelu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
      & Gelu_for_7_else_slc_32_svs;
  assign Gelu_for_else_and_13_m1c_mx1 = MUX_s_1_2_2(Gelu_for_else_and_13_m1c, Gelu_for_else_and_13_tmp,
      Gelu_for_7_slc_32_1_svs);
  assign Gelu_for_else_and_15_tmp = Gelu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
      & Gelu_for_8_else_slc_32_svs;
  assign Gelu_for_else_and_15_m1c_mx1 = MUX_s_1_2_2(Gelu_for_else_and_15_m1c, Gelu_for_else_and_15_tmp,
      Gelu_for_8_slc_32_1_svs);
  assign Gelu_for_else_and_17_tmp = Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & Gelu_for_9_else_slc_32_svs;
  assign Gelu_for_else_and_17_m1c_mx1 = MUX_s_1_2_2(Gelu_for_else_and_17_m1c, Gelu_for_else_and_17_tmp,
      Gelu_for_9_slc_32_1_svs);
  assign Gelu_for_else_and_19_tmp = Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & Gelu_for_10_else_slc_32_svs;
  assign Gelu_for_else_and_19_m1c_mx1 = MUX_s_1_2_2(Gelu_for_else_and_19_m1c, Gelu_for_else_and_19_tmp,
      Gelu_for_10_slc_32_1_svs);
  assign Gelu_for_else_and_21_tmp = Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & Gelu_for_11_else_slc_32_svs;
  assign Gelu_for_else_and_21_m1c_mx1 = MUX_s_1_2_2(Gelu_for_else_and_21_m1c, Gelu_for_else_and_21_tmp,
      Gelu_for_11_slc_32_1_svs);
  assign Gelu_for_else_and_23_tmp = Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & Gelu_for_12_else_slc_32_svs;
  assign Gelu_for_else_and_23_m1c_mx1 = MUX_s_1_2_2(Gelu_for_else_and_23_m1c, Gelu_for_else_and_23_tmp,
      Gelu_for_12_slc_32_1_svs);
  assign Gelu_for_else_and_25_tmp = Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & Gelu_for_13_else_slc_32_svs;
  assign Gelu_for_else_and_25_m1c_mx1 = MUX_s_1_2_2(Gelu_for_else_and_25_m1c, Gelu_for_else_and_25_tmp,
      Gelu_for_13_slc_32_1_svs);
  assign Gelu_for_else_and_27_tmp = Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & Gelu_for_14_else_slc_32_svs;
  assign Gelu_for_else_and_27_m1c_mx1 = MUX_s_1_2_2(Gelu_for_else_and_27_m1c, Gelu_for_else_and_27_tmp,
      Gelu_for_14_slc_32_1_svs);
  assign Gelu_for_else_and_29_tmp = Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & Gelu_for_15_else_slc_32_svs;
  assign Gelu_for_else_and_29_m1c_mx1 = MUX_s_1_2_2(Gelu_for_else_and_29_m1c, Gelu_for_else_and_29_tmp,
      Gelu_for_15_slc_32_1_svs);
  assign Gelu_for_else_and_31_tmp = Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & Gelu_for_16_else_slc_32_svs;
  assign Gelu_for_else_and_31_m1c_mx1 = MUX_s_1_2_2(Gelu_for_else_and_31_m1c, Gelu_for_else_and_31_tmp,
      Gelu_for_16_slc_32_1_svs);
  assign nl_act_read_addrs_sva_2_mx0w0 = ({(act_config_output_counter_sva_7_4[0])
      , act_config_output_counter_sva_3 , act_config_output_counter_sva_2_0}) + act_config_buffer_addr_base_sva;
  assign act_read_addrs_sva_2_mx0w0 = nl_act_read_addrs_sva_2_mx0w0[4:0];
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_2_mx0w2 = act_read_addrs_lpi_1_dfm_7
      & ({{4{ActUnit_DecodeAxiRead_unequal_tmp_1}}, ActUnit_DecodeAxiRead_unequal_tmp_1})
      & ({{4{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}}, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt})
      & ({{4{rva_in_PopNB_mioi_return_rsc_z_mxwt}}, rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign Tanh_for_and_1_cse_sva_mx0w0 = (act_config_in_InstFetch_return_sva_7_2[1:0]==2'b01);
  assign Tanh_for_and_2_cse_sva_mx0w0 = (act_config_in_InstFetch_return_sva_7_2[1:0]==2'b11);
  assign ActUnit_RunInst_switch_lp_equal_tmp_1_mx0w0 = (act_config_in_InstFetch_mux_tmp[7:4]==4'b0010);
  assign ActUnit_RunInst_switch_lp_equal_tmp_2_mx0w0 = (act_config_in_InstFetch_mux_tmp[7:4]==4'b0011);
  assign ActUnit_RunInst_switch_lp_equal_tmp_3_mx0w0 = (act_config_in_InstFetch_mux_tmp[7:4]==4'b0100);
  assign ActUnit_RunInst_switch_lp_equal_tmp_4_mx0w0 = (act_config_in_InstFetch_mux_tmp[7:4]==4'b0111);
  assign ActUnit_RunInst_switch_lp_equal_tmp_5_mx0w0 = (act_config_in_InstFetch_mux_tmp[7:4]==4'b1011);
  assign ActUnit_RunInst_switch_lp_equal_tmp_6_mx0w0 = (act_config_in_InstFetch_mux_tmp[7:4]==4'b1100);
  assign ActUnit_RunInst_switch_lp_equal_tmp_7_mx0w0 = (act_config_in_InstFetch_mux_tmp[7:4]==4'b1110);
  assign ActUnit_RunInst_switch_lp_equal_tmp_8_mx0w0 = (act_config_in_InstFetch_mux_tmp[7:4]==4'b1111);
  assign ActUnit_RunInst_switch_lp_nor_nl = ~(ActUnit_RunInst_switch_lp_equal_tmp_9
      | ActUnit_RunInst_switch_lp_equal_tmp_1_mx0w0 | ActUnit_RunInst_switch_lp_equal_tmp_2_mx0w0
      | ActUnit_RunInst_switch_lp_equal_tmp_3_mx0w0 | ActUnit_RunInst_switch_lp_equal_tmp_4_mx0w0
      | ActUnit_RunInst_switch_lp_equal_tmp_5_mx0w0 | ActUnit_RunInst_switch_lp_equal_tmp_6_mx0w0
      | ActUnit_RunInst_switch_lp_equal_tmp_7_mx0w0 | ActUnit_RunInst_switch_lp_equal_tmp_8_mx0w0);
  assign ActUnit_RunInst_switch_lp_nor_tmp_mx0 = MUX_s_1_2_2(ActUnit_RunInst_switch_lp_nor_nl,
      ActUnit_RunInst_switch_lp_nor_tmp, or_dcpl_823);
  assign nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      = MUX_s_1_4_2(reg_act_regs_data_0_0_ftd, act_regs_data_1_0_sva_31, act_regs_data_2_0_sva_31,
      act_regs_data_3_0_sva_31, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      = MUX_v_5_4_2(reg_act_regs_data_0_0_ftd_1, act_regs_data_1_0_sva_30_26, act_regs_data_2_0_sva_30_26,
      act_regs_data_3_0_sva_30_26, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm
      = MUX_v_22_4_2(reg_act_regs_data_0_0_ftd_3, act_regs_data_1_0_sva_21_0, act_regs_data_2_0_sva_21_0,
      act_regs_data_3_0_sva_21_0, act_config_in_InstFetch_mux_tmp[3:2]);
  assign Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs_mx0w0
      = $signed(1'b0) < $signed(({nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      = MUX_s_1_4_2(reg_act_regs_data_0_1_ftd, act_regs_data_1_1_sva_31, act_regs_data_2_1_sva_31,
      act_regs_data_3_1_sva_31, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      = MUX_v_5_4_2(reg_act_regs_data_0_1_ftd_1, act_regs_data_1_1_sva_30_26, act_regs_data_2_1_sva_30_26,
      act_regs_data_3_1_sva_30_26, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm
      = MUX_v_22_4_2(reg_act_regs_data_0_1_ftd_3, act_regs_data_1_1_sva_21_0, act_regs_data_2_1_sva_21_0,
      act_regs_data_3_1_sva_21_0, act_config_in_InstFetch_mux_tmp[3:2]);
  assign Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs_mx0w0
      = $signed(1'b0) < $signed(({nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      = MUX_s_1_4_2(act_regs_data_0_2_sva_31, act_regs_data_1_2_sva_31, act_regs_data_2_2_sva_31,
      act_regs_data_3_2_sva_31, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      = MUX_v_5_4_2(act_regs_data_0_2_sva_30_26, act_regs_data_1_2_sva_30_26, act_regs_data_2_2_sva_30_26,
      act_regs_data_3_2_sva_30_26, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm
      = MUX_v_22_4_2(act_regs_data_0_2_sva_21_0, act_regs_data_1_2_sva_21_0, act_regs_data_2_2_sva_21_0,
      act_regs_data_3_2_sva_21_0, act_config_in_InstFetch_mux_tmp[3:2]);
  assign Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs_mx0w0
      = $signed(1'b0) < $signed(({nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      = MUX_s_1_4_2(act_regs_data_0_3_sva_31, act_regs_data_1_3_sva_31, act_regs_data_2_3_sva_31,
      act_regs_data_3_3_sva_31, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      = MUX_v_5_4_2(act_regs_data_0_3_sva_30_26, act_regs_data_1_3_sva_30_26, act_regs_data_2_3_sva_30_26,
      act_regs_data_3_3_sva_30_26, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm
      = MUX_v_22_4_2(act_regs_data_0_3_sva_21_0, act_regs_data_1_3_sva_21_0, act_regs_data_2_3_sva_21_0,
      act_regs_data_3_3_sva_21_0, act_config_in_InstFetch_mux_tmp[3:2]);
  assign Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs_mx0w0
      = $signed(1'b0) < $signed(({nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      = MUX_s_1_4_2(act_regs_data_0_4_sva_31, act_regs_data_1_4_sva_31, act_regs_data_2_4_sva_31,
      act_regs_data_3_4_sva_31, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      = MUX_v_5_4_2(act_regs_data_0_4_sva_30_26, act_regs_data_1_4_sva_30_26, act_regs_data_2_4_sva_30_26,
      act_regs_data_3_4_sva_30_26, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm
      = MUX_v_22_4_2(act_regs_data_0_4_sva_21_0, act_regs_data_1_4_sva_21_0, act_regs_data_2_4_sva_21_0,
      act_regs_data_3_4_sva_21_0, act_config_in_InstFetch_mux_tmp[3:2]);
  assign Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs_mx0w0
      = $signed(1'b0) < $signed(({nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      = MUX_s_1_4_2(act_regs_data_0_5_sva_31, act_regs_data_1_5_sva_31, act_regs_data_2_5_sva_31,
      act_regs_data_3_5_sva_31, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      = MUX_v_5_4_2(act_regs_data_0_5_sva_30_26, act_regs_data_1_5_sva_30_26, act_regs_data_2_5_sva_30_26,
      act_regs_data_3_5_sva_30_26, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm
      = MUX_v_22_4_2(act_regs_data_0_5_sva_21_0, act_regs_data_1_5_sva_21_0, act_regs_data_2_5_sva_21_0,
      act_regs_data_3_5_sva_21_0, act_config_in_InstFetch_mux_tmp[3:2]);
  assign Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs_mx0w0
      = $signed(1'b0) < $signed(({nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      = MUX_s_1_4_2(act_regs_data_0_6_sva_31, act_regs_data_1_6_sva_31, act_regs_data_2_6_sva_31,
      act_regs_data_3_6_sva_31, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      = MUX_v_5_4_2(act_regs_data_0_6_sva_30_26, act_regs_data_1_6_sva_30_26, act_regs_data_2_6_sva_30_26,
      act_regs_data_3_6_sva_30_26, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm
      = MUX_v_22_4_2(act_regs_data_0_6_sva_21_0, act_regs_data_1_6_sva_21_0, act_regs_data_2_6_sva_21_0,
      act_regs_data_3_6_sva_21_0, act_config_in_InstFetch_mux_tmp[3:2]);
  assign Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs_mx0w0
      = $signed(1'b0) < $signed(({nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      = MUX_s_1_4_2(act_regs_data_0_7_sva_31, act_regs_data_1_7_sva_31, act_regs_data_2_7_sva_31,
      act_regs_data_3_7_sva_31, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      = MUX_v_5_4_2(act_regs_data_0_7_sva_30_26, act_regs_data_1_7_sva_30_26, act_regs_data_2_7_sva_30_26,
      act_regs_data_3_7_sva_30_26, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm
      = MUX_v_22_4_2(act_regs_data_0_7_sva_21_0, act_regs_data_1_7_sva_21_0, act_regs_data_2_7_sva_21_0,
      act_regs_data_3_7_sva_21_0, act_config_in_InstFetch_mux_tmp[3:2]);
  assign Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs_mx0w0
      = $signed(1'b0) < $signed(({nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      = MUX_s_1_4_2(act_regs_data_0_8_sva_31, act_regs_data_1_8_sva_31, act_regs_data_2_8_sva_31,
      act_regs_data_3_8_sva_31, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      = MUX_v_5_4_2(act_regs_data_0_8_sva_30_26, act_regs_data_1_8_sva_30_26, act_regs_data_2_8_sva_30_26,
      act_regs_data_3_8_sva_30_26, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm
      = MUX_v_22_4_2(act_regs_data_0_8_sva_21_0, act_regs_data_1_8_sva_21_0, act_regs_data_2_8_sva_21_0,
      act_regs_data_3_8_sva_21_0, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      = MUX_s_1_4_2(act_regs_data_0_9_sva_31, act_regs_data_1_9_sva_31, act_regs_data_2_9_sva_31,
      act_regs_data_3_9_sva_31, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      = MUX_v_5_4_2(act_regs_data_0_9_sva_30_26, act_regs_data_1_9_sva_30_26, act_regs_data_2_9_sva_30_26,
      act_regs_data_3_9_sva_30_26, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm
      = MUX_v_22_4_2(act_regs_data_0_9_sva_21_0, act_regs_data_1_9_sva_21_0, act_regs_data_2_9_sva_21_0,
      act_regs_data_3_9_sva_21_0, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      = MUX_s_1_4_2(reg_act_regs_data_0_10_ftd, act_regs_data_1_10_sva_31, act_regs_data_2_10_sva_31,
      act_regs_data_3_10_sva_31, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      = MUX_v_5_4_2(reg_act_regs_data_0_10_ftd_1, act_regs_data_1_10_sva_30_26, act_regs_data_2_10_sva_30_26,
      act_regs_data_3_10_sva_30_26, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm
      = MUX_v_22_4_2(reg_act_regs_data_0_10_ftd_3, act_regs_data_1_10_sva_21_0, act_regs_data_2_10_sva_21_0,
      act_regs_data_3_10_sva_21_0, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      = MUX_s_1_4_2(reg_act_regs_data_0_11_ftd, act_regs_data_1_11_sva_31, act_regs_data_2_11_sva_31,
      act_regs_data_3_11_sva_31, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      = MUX_v_5_4_2(reg_act_regs_data_0_11_ftd_1, act_regs_data_1_11_sva_30_26, act_regs_data_2_11_sva_30_26,
      act_regs_data_3_11_sva_30_26, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm
      = MUX_v_22_4_2(reg_act_regs_data_0_11_ftd_3, act_regs_data_1_11_sva_21_0, act_regs_data_2_11_sva_21_0,
      act_regs_data_3_11_sva_21_0, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      = MUX_s_1_4_2(reg_act_regs_data_0_12_ftd, act_regs_data_1_12_sva_31, act_regs_data_2_12_sva_31,
      act_regs_data_3_12_sva_31, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      = MUX_v_5_4_2(reg_act_regs_data_0_12_ftd_1, act_regs_data_1_12_sva_30_26, act_regs_data_2_12_sva_30_26,
      act_regs_data_3_12_sva_30_26, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm
      = MUX_v_22_4_2(reg_act_regs_data_0_12_ftd_3, act_regs_data_1_12_sva_21_0, act_regs_data_2_12_sva_21_0,
      act_regs_data_3_12_sva_21_0, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      = MUX_s_1_4_2(reg_act_regs_data_0_13_ftd, act_regs_data_1_13_sva_31, act_regs_data_2_13_sva_31,
      act_regs_data_3_13_sva_31, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      = MUX_v_5_4_2(reg_act_regs_data_0_13_ftd_1, act_regs_data_1_13_sva_30_26, act_regs_data_2_13_sva_30_26,
      act_regs_data_3_13_sva_30_26, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm
      = MUX_v_22_4_2(reg_act_regs_data_0_13_ftd_3, act_regs_data_1_13_sva_21_0, act_regs_data_2_13_sva_21_0,
      act_regs_data_3_13_sva_21_0, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      = MUX_s_1_4_2(act_regs_data_0_14_sva_31, act_regs_data_1_14_sva_31, act_regs_data_2_14_sva_31,
      act_regs_data_3_14_sva_31, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      = MUX_v_5_4_2(act_regs_data_0_14_sva_30_26, act_regs_data_1_14_sva_30_26, act_regs_data_2_14_sva_30_26,
      act_regs_data_3_14_sva_30_26, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm
      = MUX_v_22_4_2(act_regs_data_0_14_sva_21_0, act_regs_data_1_14_sva_21_0, act_regs_data_2_14_sva_21_0,
      act_regs_data_3_14_sva_21_0, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      = MUX_s_1_4_2(act_regs_data_0_15_sva_31, act_regs_data_1_15_sva_31, act_regs_data_2_15_sva_31,
      act_regs_data_3_15_sva_31, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      = MUX_v_5_4_2(act_regs_data_0_15_sva_30_26, act_regs_data_1_15_sva_30_26, act_regs_data_2_15_sva_30_26,
      act_regs_data_3_15_sva_30_26, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm
      = MUX_v_22_4_2(act_regs_data_0_15_sva_21_0, act_regs_data_1_15_sva_21_0, act_regs_data_2_15_sva_21_0,
      act_regs_data_3_15_sva_21_0, act_config_in_InstFetch_mux_tmp[3:2]);
  assign act_config_in_InstFetch_mux_tmp = MUX_v_8_32_2(act_config_inst_regs_0_sva_dfm_5,
      act_config_inst_regs_1_sva_dfm_5, act_config_inst_regs_2_sva_dfm_5, act_config_inst_regs_3_sva_dfm_5,
      act_config_inst_regs_4_sva_dfm_5, act_config_inst_regs_5_sva_dfm_5, act_config_inst_regs_6_sva_dfm_5,
      act_config_inst_regs_7_sva_dfm_5, act_config_inst_regs_8_sva_dfm_5, act_config_inst_regs_9_sva_dfm_5,
      act_config_inst_regs_10_sva_dfm_5, act_config_inst_regs_11_sva_dfm_5, act_config_inst_regs_12_sva_dfm_5,
      act_config_inst_regs_13_sva_dfm_5, act_config_inst_regs_14_sva_dfm_5, act_config_inst_regs_15_sva_dfm_5,
      act_config_inst_regs_16_sva_dfm_6, act_config_inst_regs_17_sva_dfm_6, act_config_inst_regs_18_sva_dfm_6,
      act_config_inst_regs_19_sva_dfm_6, act_config_inst_regs_20_sva_dfm_6, act_config_inst_regs_21_sva_dfm_6,
      act_config_inst_regs_22_sva_dfm_6, act_config_inst_regs_23_sva_dfm_6, act_config_inst_regs_24_sva_dfm_6,
      act_config_inst_regs_25_sva_dfm_6, act_config_inst_regs_26_sva_dfm_6, act_config_inst_regs_27_sva_dfm_6,
      act_config_inst_regs_28_sva_dfm_6, act_config_inst_regs_29_sva_dfm_6, act_config_inst_regs_30_sva_dfm_6,
      act_config_inst_regs_31_sva_dfm_6, act_config_inst_counter_sva);
  assign operator_32_8_true_AC_TRN_AC_WRAP_less_tmp = $signed(27'b100000000000000000000000000)
      < $signed(({nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign operator_32_8_true_AC_TRN_AC_WRAP_less_1_tmp = $signed(27'b100000000000000000000000000)
      < $signed(({nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign operator_32_8_true_AC_TRN_AC_WRAP_less_2_tmp = $signed(27'b100000000000000000000000000)
      < $signed(({nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign operator_32_8_true_AC_TRN_AC_WRAP_less_3_tmp = $signed(27'b100000000000000000000000000)
      < $signed(({nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign operator_32_8_true_AC_TRN_AC_WRAP_less_4_tmp = $signed(27'b100000000000000000000000000)
      < $signed(({nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign operator_32_8_true_AC_TRN_AC_WRAP_less_5_tmp = $signed(27'b100000000000000000000000000)
      < $signed(({nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign operator_32_8_true_AC_TRN_AC_WRAP_less_6_tmp = $signed(27'b100000000000000000000000000)
      < $signed(({nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign operator_32_8_true_AC_TRN_AC_WRAP_less_7_tmp = $signed(27'b100000000000000000000000000)
      < $signed(({nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign operator_32_8_true_AC_TRN_AC_WRAP_less_8_tmp = $signed(27'b100000000000000000000000000)
      < $signed(({nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign operator_32_8_true_AC_TRN_AC_WRAP_less_9_tmp = $signed(27'b100000000000000000000000000)
      < $signed(({nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign operator_32_8_true_AC_TRN_AC_WRAP_less_10_tmp = $signed(27'b100000000000000000000000000)
      < $signed(({nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign operator_32_8_true_AC_TRN_AC_WRAP_less_11_tmp = $signed(27'b100000000000000000000000000)
      < $signed(({nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign operator_32_8_true_AC_TRN_AC_WRAP_less_12_tmp = $signed(27'b100000000000000000000000000)
      < $signed(({nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign operator_32_8_true_AC_TRN_AC_WRAP_less_13_tmp = $signed(27'b100000000000000000000000000)
      < $signed(({nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign operator_32_8_true_AC_TRN_AC_WRAP_less_14_tmp = $signed(27'b100000000000000000000000000)
      < $signed(({nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign operator_32_8_true_AC_TRN_AC_WRAP_less_15_tmp = $signed(27'b100000000000000000000000000)
      < $signed(({nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign Gelu_for_if_less_tmp = $signed(27'b101100000000000000000000000) < $signed(({nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign Gelu_for_if_less_1_tmp = $signed(27'b101100000000000000000000000) < $signed(({nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign Gelu_for_if_less_2_tmp = $signed(27'b101100000000000000000000000) < $signed(({nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign Gelu_for_if_less_3_tmp = $signed(27'b101100000000000000000000000) < $signed(({nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign Gelu_for_if_less_4_tmp = $signed(27'b101100000000000000000000000) < $signed(({nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign Gelu_for_if_less_5_tmp = $signed(27'b101100000000000000000000000) < $signed(({nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign Gelu_for_if_less_6_tmp = $signed(27'b101100000000000000000000000) < $signed(({nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign Gelu_for_if_less_7_tmp = $signed(27'b101100000000000000000000000) < $signed(({nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign Gelu_for_if_less_8_tmp = $signed(27'b101100000000000000000000000) < $signed(({nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign Gelu_for_if_less_9_tmp = $signed(27'b101100000000000000000000000) < $signed(({nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign Gelu_for_if_less_10_tmp = $signed(27'b101100000000000000000000000) < $signed(({nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign Gelu_for_if_less_11_tmp = $signed(27'b101100000000000000000000000) < $signed(({nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign Gelu_for_if_less_12_tmp = $signed(27'b101100000000000000000000000) < $signed(({nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign Gelu_for_if_less_13_tmp = $signed(27'b101100000000000000000000000) < $signed(({nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign Gelu_for_if_less_14_tmp = $signed(27'b101100000000000000000000000) < $signed(({nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign Gelu_for_if_less_15_tmp = $signed(27'b101100000000000000000000000) < $signed(({nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      , nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
  assign ActUnit_RunInst_switch_lp_equal_tmp_9 = (act_config_in_InstFetch_mux_tmp[7:4]==4'b0001);
  assign Tanh_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1
      = $signed(({nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , (nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0[2])}))
      < $signed(1'b1);
  assign Tanh_for_15_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1
      = $signed(({nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , (nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0[2])}))
      < $signed(1'b1);
  assign Tanh_for_14_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1
      = $signed(({nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , (nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0[2])}))
      < $signed(1'b1);
  assign Tanh_for_13_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1
      = $signed(({nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , (nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0[2])}))
      < $signed(1'b1);
  assign Tanh_for_12_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1
      = $signed(({nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , (nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0[2])}))
      < $signed(1'b1);
  assign Tanh_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1
      = $signed(({nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , (nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0[2])}))
      < $signed(1'b1);
  assign Tanh_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1
      = $signed(({nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , (nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0[2])}))
      < $signed(1'b1);
  assign Tanh_for_9_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1
      = $signed(({nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , (nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0[2])}))
      < $signed(1'b1);
  assign Tanh_for_8_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1
      = $signed(({nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , (nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0[2])}))
      < $signed(1'b1);
  assign Tanh_for_7_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1
      = $signed(({nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , (nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0[2])}))
      < $signed(1'b1);
  assign Tanh_for_6_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1
      = $signed(({nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , (nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0[2])}))
      < $signed(1'b1);
  assign Tanh_for_5_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1
      = $signed(({nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , (nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0[2])}))
      < $signed(1'b1);
  assign Tanh_for_4_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1
      = $signed(({nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , (nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0[2])}))
      < $signed(1'b1);
  assign Tanh_for_3_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1
      = $signed(({nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , (nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0[2])}))
      < $signed(1'b1);
  assign Tanh_for_2_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1
      = $signed(({nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , (nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0[2])}))
      < $signed(1'b1);
  assign Tanh_for_1_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1
      = $signed(({nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
      , nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
      , nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      , (nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0[2])}))
      < $signed(1'b1);
  assign ActUnit_RunInst_switch_lp_and_32_tmp_mx0w1 = (act_config_in_InstFetch_return_sva_7_2[1:0]==2'b10)
      & act_port_PopNB_mioi_return_rsc_z_mxwt;
  assign ActUnit_RunInst_switch_lp_and_16_tmp_mx0w1 = (act_config_in_InstFetch_return_sva_7_2[1:0]==2'b01)
      & act_port_PopNB_mioi_return_rsc_z_mxwt;
  assign act_config_InstIncr_if_equal_1_tmp = act_config_inst_counter_sva_dfm_3 ==
      (operator_6_false_acc_tmp[4:0]);
  assign act_config_InstIncr_act_config_InstIncr_if_and_svs_1 = act_config_InstIncr_if_equal_1_tmp
      & nor_447_cse;
  assign ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_30_26_2 =
      MUX_v_5_64_2(act_regs_data_0_0_sva_dfm_2_30_26, act_regs_data_0_1_sva_dfm_2_30_26,
      act_regs_data_0_2_sva_dfm_2_30_26, act_regs_data_0_3_sva_dfm_2_30_26, act_regs_data_0_4_sva_dfm_2_30_26,
      act_regs_data_0_5_sva_dfm_2_30_26, act_regs_data_0_6_sva_dfm_2_30_26, act_regs_data_0_7_sva_dfm_2_30_26,
      act_regs_data_0_8_sva_dfm_2_30_26, act_regs_data_0_9_sva_dfm_2_30_26, act_regs_data_0_10_sva_dfm_2_30_26,
      act_regs_data_0_11_sva_dfm_2_30_26, act_regs_data_0_12_sva_dfm_2_30_26, act_regs_data_0_13_sva_dfm_2_30_26,
      act_regs_data_0_14_sva_dfm_2_30_26, act_regs_data_0_15_sva_dfm_2_30_26, act_regs_data_1_0_sva_dfm_2_30_26,
      act_regs_data_1_1_sva_dfm_2_30_26, act_regs_data_1_2_sva_dfm_2_30_26, act_regs_data_1_3_sva_dfm_2_30_26,
      act_regs_data_1_4_sva_dfm_2_30_26, act_regs_data_1_5_sva_dfm_2_30_26, act_regs_data_1_6_sva_dfm_2_30_26,
      act_regs_data_1_7_sva_dfm_2_30_26, act_regs_data_1_8_sva_dfm_2_30_26, act_regs_data_1_9_sva_dfm_2_30_26,
      act_regs_data_1_10_sva_dfm_2_30_26, act_regs_data_1_11_sva_dfm_2_30_26, act_regs_data_1_12_sva_dfm_2_30_26,
      act_regs_data_1_13_sva_dfm_2_30_26, act_regs_data_1_14_sva_dfm_2_30_26, act_regs_data_1_15_sva_dfm_2_30_26,
      act_regs_data_2_0_sva_dfm_2_30_26, act_regs_data_2_1_sva_dfm_2_30_26, act_regs_data_2_2_sva_dfm_2_30_26,
      act_regs_data_2_3_sva_dfm_2_30_26, act_regs_data_2_4_sva_dfm_2_30_26, act_regs_data_2_5_sva_dfm_2_30_26,
      act_regs_data_2_6_sva_dfm_2_30_26, act_regs_data_2_7_sva_dfm_2_30_26, act_regs_data_2_8_sva_dfm_2_30_26,
      act_regs_data_2_9_sva_dfm_2_30_26, act_regs_data_2_10_sva_dfm_2_30_26, act_regs_data_2_11_sva_dfm_2_30_26,
      act_regs_data_2_12_sva_dfm_2_30_26, act_regs_data_2_13_sva_dfm_2_30_26, act_regs_data_2_14_sva_dfm_2_30_26,
      act_regs_data_2_15_sva_dfm_2_30_26, act_regs_data_3_0_sva_dfm_2_30_26, act_regs_data_3_1_sva_dfm_2_30_26,
      act_regs_data_3_2_sva_dfm_2_30_26, act_regs_data_3_3_sva_dfm_2_30_26, act_regs_data_3_4_sva_dfm_2_30_26,
      act_regs_data_3_5_sva_dfm_2_30_26, act_regs_data_3_6_sva_dfm_2_30_26, act_regs_data_3_7_sva_dfm_2_30_26,
      act_regs_data_3_8_sva_dfm_2_30_26, act_regs_data_3_9_sva_dfm_2_30_26, act_regs_data_3_10_sva_dfm_2_30_26,
      act_regs_data_3_11_sva_dfm_2_30_26, act_regs_data_3_12_sva_dfm_2_30_26, act_regs_data_3_13_sva_dfm_2_30_26,
      act_regs_data_3_14_sva_dfm_2_30_26, act_regs_data_3_15_sva_dfm_2_30_26, {nvhls_get_slc_2U_NVUINT8_return_2_sva
      , ActUnit_PushOutput_if_for_i_4_0_sva_3_0});
  assign ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_31 = MUX_s_1_64_2(reg_act_regs_data_0_0_ftd,
      reg_act_regs_data_0_1_ftd, act_regs_data_0_2_sva_31, act_regs_data_0_3_sva_31,
      act_regs_data_0_4_sva_31, act_regs_data_0_5_sva_31, act_regs_data_0_6_sva_31,
      act_regs_data_0_7_sva_31, act_regs_data_0_8_sva_31, act_regs_data_0_9_sva_31,
      reg_act_regs_data_0_10_ftd, reg_act_regs_data_0_11_ftd, reg_act_regs_data_0_12_ftd,
      reg_act_regs_data_0_13_ftd, act_regs_data_0_14_sva_31, act_regs_data_0_15_sva_31,
      act_regs_data_1_0_sva_31, act_regs_data_1_1_sva_31, act_regs_data_1_2_sva_31,
      act_regs_data_1_3_sva_31, act_regs_data_1_4_sva_31, act_regs_data_1_5_sva_31,
      act_regs_data_1_6_sva_31, act_regs_data_1_7_sva_31, act_regs_data_1_8_sva_31,
      act_regs_data_1_9_sva_31, act_regs_data_1_10_sva_31, act_regs_data_1_11_sva_31,
      act_regs_data_1_12_sva_31, act_regs_data_1_13_sva_31, act_regs_data_1_14_sva_31,
      act_regs_data_1_15_sva_31, act_regs_data_2_0_sva_31, act_regs_data_2_1_sva_31,
      act_regs_data_2_2_sva_31, act_regs_data_2_3_sva_31, act_regs_data_2_4_sva_31,
      act_regs_data_2_5_sva_31, act_regs_data_2_6_sva_31, act_regs_data_2_7_sva_31,
      act_regs_data_2_8_sva_31, act_regs_data_2_9_sva_31, act_regs_data_2_10_sva_31,
      act_regs_data_2_11_sva_31, act_regs_data_2_12_sva_31, act_regs_data_2_13_sva_31,
      act_regs_data_2_14_sva_31, act_regs_data_2_15_sva_31, act_regs_data_3_0_sva_31,
      act_regs_data_3_1_sva_31, act_regs_data_3_2_sva_31, act_regs_data_3_3_sva_31,
      act_regs_data_3_4_sva_31, act_regs_data_3_5_sva_31, act_regs_data_3_6_sva_31,
      act_regs_data_3_7_sva_31, act_regs_data_3_8_sva_31, act_regs_data_3_9_sva_31,
      act_regs_data_3_10_sva_31, act_regs_data_3_11_sva_31, act_regs_data_3_12_sva_31,
      act_regs_data_3_13_sva_31, act_regs_data_3_14_sva_31, act_regs_data_3_15_sva_31,
      {(act_config_in_InstFetch_return_sva_7_2[1:0]) , ActUnit_PushOutput_if_for_i_4_0_sva_3_0});
  assign ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_30_26
      = MUX_v_5_64_2(reg_act_regs_data_0_0_ftd_1, reg_act_regs_data_0_1_ftd_1, act_regs_data_0_2_sva_30_26,
      act_regs_data_0_3_sva_30_26, act_regs_data_0_4_sva_30_26, act_regs_data_0_5_sva_30_26,
      act_regs_data_0_6_sva_30_26, act_regs_data_0_7_sva_30_26, act_regs_data_0_8_sva_30_26,
      act_regs_data_0_9_sva_30_26, reg_act_regs_data_0_10_ftd_1, reg_act_regs_data_0_11_ftd_1,
      reg_act_regs_data_0_12_ftd_1, reg_act_regs_data_0_13_ftd_1, act_regs_data_0_14_sva_30_26,
      act_regs_data_0_15_sva_30_26, act_regs_data_1_0_sva_30_26, act_regs_data_1_1_sva_30_26,
      act_regs_data_1_2_sva_30_26, act_regs_data_1_3_sva_30_26, act_regs_data_1_4_sva_30_26,
      act_regs_data_1_5_sva_30_26, act_regs_data_1_6_sva_30_26, act_regs_data_1_7_sva_30_26,
      act_regs_data_1_8_sva_30_26, act_regs_data_1_9_sva_30_26, act_regs_data_1_10_sva_30_26,
      act_regs_data_1_11_sva_30_26, act_regs_data_1_12_sva_30_26, act_regs_data_1_13_sva_30_26,
      act_regs_data_1_14_sva_30_26, act_regs_data_1_15_sva_30_26, act_regs_data_2_0_sva_30_26,
      act_regs_data_2_1_sva_30_26, act_regs_data_2_2_sva_30_26, act_regs_data_2_3_sva_30_26,
      act_regs_data_2_4_sva_30_26, act_regs_data_2_5_sva_30_26, act_regs_data_2_6_sva_30_26,
      act_regs_data_2_7_sva_30_26, act_regs_data_2_8_sva_30_26, act_regs_data_2_9_sva_30_26,
      act_regs_data_2_10_sva_30_26, act_regs_data_2_11_sva_30_26, act_regs_data_2_12_sva_30_26,
      act_regs_data_2_13_sva_30_26, act_regs_data_2_14_sva_30_26, act_regs_data_2_15_sva_30_26,
      act_regs_data_3_0_sva_30_26, act_regs_data_3_1_sva_30_26, act_regs_data_3_2_sva_30_26,
      act_regs_data_3_3_sva_30_26, act_regs_data_3_4_sva_30_26, act_regs_data_3_5_sva_30_26,
      act_regs_data_3_6_sva_30_26, act_regs_data_3_7_sva_30_26, act_regs_data_3_8_sva_30_26,
      act_regs_data_3_9_sva_30_26, act_regs_data_3_10_sva_30_26, act_regs_data_3_11_sva_30_26,
      act_regs_data_3_12_sva_30_26, act_regs_data_3_13_sva_30_26, act_regs_data_3_14_sva_30_26,
      act_regs_data_3_15_sva_30_26, {(act_config_in_InstFetch_return_sva_7_2[1:0])
      , ActUnit_PushOutput_if_for_i_4_0_sva_3_0});
  assign ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_21_0 =
      MUX_v_22_64_2(reg_act_regs_data_0_0_ftd_3, reg_act_regs_data_0_1_ftd_3, act_regs_data_0_2_sva_21_0,
      act_regs_data_0_3_sva_21_0, act_regs_data_0_4_sva_21_0, act_regs_data_0_5_sva_21_0,
      act_regs_data_0_6_sva_21_0, act_regs_data_0_7_sva_21_0, act_regs_data_0_8_sva_21_0,
      act_regs_data_0_9_sva_21_0, reg_act_regs_data_0_10_ftd_3, reg_act_regs_data_0_11_ftd_3,
      reg_act_regs_data_0_12_ftd_3, reg_act_regs_data_0_13_ftd_3, act_regs_data_0_14_sva_21_0,
      act_regs_data_0_15_sva_21_0, act_regs_data_1_0_sva_21_0, act_regs_data_1_1_sva_21_0,
      act_regs_data_1_2_sva_21_0, act_regs_data_1_3_sva_21_0, act_regs_data_1_4_sva_21_0,
      act_regs_data_1_5_sva_21_0, act_regs_data_1_6_sva_21_0, act_regs_data_1_7_sva_21_0,
      act_regs_data_1_8_sva_21_0, act_regs_data_1_9_sva_21_0, act_regs_data_1_10_sva_21_0,
      act_regs_data_1_11_sva_21_0, act_regs_data_1_12_sva_21_0, act_regs_data_1_13_sva_21_0,
      act_regs_data_1_14_sva_21_0, act_regs_data_1_15_sva_21_0, act_regs_data_2_0_sva_21_0,
      act_regs_data_2_1_sva_21_0, act_regs_data_2_2_sva_21_0, act_regs_data_2_3_sva_21_0,
      act_regs_data_2_4_sva_21_0, act_regs_data_2_5_sva_21_0, act_regs_data_2_6_sva_21_0,
      act_regs_data_2_7_sva_21_0, act_regs_data_2_8_sva_21_0, act_regs_data_2_9_sva_21_0,
      act_regs_data_2_10_sva_21_0, act_regs_data_2_11_sva_21_0, act_regs_data_2_12_sva_21_0,
      act_regs_data_2_13_sva_21_0, act_regs_data_2_14_sva_21_0, act_regs_data_2_15_sva_21_0,
      act_regs_data_3_0_sva_21_0, act_regs_data_3_1_sva_21_0, act_regs_data_3_2_sva_21_0,
      act_regs_data_3_3_sva_21_0, act_regs_data_3_4_sva_21_0, act_regs_data_3_5_sva_21_0,
      act_regs_data_3_6_sva_21_0, act_regs_data_3_7_sva_21_0, act_regs_data_3_8_sva_21_0,
      act_regs_data_3_9_sva_21_0, act_regs_data_3_10_sva_21_0, act_regs_data_3_11_sva_21_0,
      act_regs_data_3_12_sva_21_0, act_regs_data_3_13_sva_21_0, act_regs_data_3_14_sva_21_0,
      act_regs_data_3_15_sva_21_0, {(act_config_in_InstFetch_return_sva_7_2[1:0])
      , ActUnit_PushOutput_if_for_i_4_0_sva_3_0});
  assign act_config_ActConfigRead_else_unequal_tmp_1 = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7:0]==8'b00000010));
  assign act_config_ActConfigRead_unequal_tmp_1 = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7:0]==8'b00000001));
  assign ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_2_tmp
      = ~(act_config_is_zero_first_sva | ActUnit_RunInst_switch_lp_and_32_tmp | ActUnit_RunInst_switch_lp_equal_tmp_2
      | ActUnit_RunInst_switch_lp_equal_tmp_3 | ActUnit_RunInst_switch_lp_equal_tmp_4
      | ActUnit_RunInst_switch_lp_equal_tmp_5 | ActUnit_RunInst_switch_lp_equal_tmp_6
      | ActUnit_RunInst_switch_lp_equal_tmp_7 | ActUnit_RunInst_switch_lp_equal_tmp_8
      | ActUnit_RunInst_switch_lp_nor_tmp);
  assign ActUnit_DecodeAxiRead_unequal_tmp_1 = ~((rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11:8]==4'b1000));
  assign ActUnit_DecodeAxi_if_or_7_tmp_1 = ActUnit_DecodeAxiRead_unequal_tmp_1 |
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_6_nl = act_read_addrs_lpi_1_dfm_7
      & ({{4{ActUnit_DecodeAxiRead_unequal_tmp_1}}, ActUnit_DecodeAxiRead_unequal_tmp_1})
      & (signext_5_1(~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)) & ({{4{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_nl = ~(ActUnit_RunInst_switch_lp_and_32_tmp
      | ActUnit_RunInst_switch_lp_equal_tmp_2 | ActUnit_RunInst_switch_lp_equal_tmp_3
      | ActUnit_RunInst_switch_lp_equal_tmp_4 | ActUnit_RunInst_switch_lp_equal_tmp_5
      | ActUnit_RunInst_switch_lp_equal_tmp_6 | ActUnit_RunInst_switch_lp_equal_tmp_7
      | ActUnit_RunInst_switch_lp_equal_tmp_8 | ActUnit_RunInst_switch_lp_nor_tmp);
  assign ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_and_18_nl = ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_30_26
      & (signext_5_1(~ act_config_is_zero_first_sva)) & (signext_5_1(ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_nl));
  assign while_mux_53_ssc_mx0 = MUX_v_5_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_6_nl,
      ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_and_18_nl, is_start_sva);
  assign while_and_88_tmp_1 = ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_mx1
      & (~ is_start_sva);
  assign ActUnit_DecodeAxiWrite_else_not_17_nl = ~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0;
  assign act_read_addrs_lpi_1_dfm_7 = MUX_v_5_2_2(5'b00000, (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4:0]),
      ActUnit_DecodeAxiWrite_else_not_17_nl);
  assign Tanh_for_nor_cse_sva_mx0w0 = ~((act_config_in_InstFetch_return_sva_7_2[1:0]!=2'b00));
  assign Tanh_for_and_cse_sva_mx0w0 = (act_config_in_InstFetch_return_sva_7_2[1:0]==2'b10);
  assign operator_32_8_true_AC_TRN_AC_WRAP_7_less_15_tmp = 26'b11000000000000000000000000
      < ({ActUnit_RunInst_case_15_nv_scvector_cctor_data_0_sva_30_26 , reg_ActUnit_RunInst_case_15_nv_scvector_cctor_data_0_ftd_rsp_0
      , reg_ActUnit_RunInst_case_15_nv_scvector_cctor_data_0_ftd_rsp_1 , reg_ActUnit_RunInst_case_15_nv_scvector_cctor_data_0_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_6_less_15_tmp = 25'b1000000000000000000000000
      < ({ActUnit_RunInst_case_15_nv_scvector_cctor_data_0_sva_30_26 , reg_ActUnit_RunInst_case_15_nv_scvector_cctor_data_0_ftd_rsp_0
      , reg_ActUnit_RunInst_case_15_nv_scvector_cctor_data_0_ftd_rsp_1 , reg_ActUnit_RunInst_case_15_nv_scvector_cctor_data_0_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_3_less_15_tmp = 26'b10000000000000000000000000
      < ({reg_ActUnit_RunInst_case_14_nv_scvector_cctor_data_0_ftd_1_30_26 , reg_ActUnit_RunInst_case_14_nv_scvector_cctor_data_0_1_ftd_rsp_0
      , reg_ActUnit_RunInst_case_14_nv_scvector_cctor_data_0_1_ftd_rsp_1 , reg_ActUnit_RunInst_case_14_nv_scvector_cctor_data_0_1_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_7_less_14_tmp = 26'b11000000000000000000000000
      < ({nv_scvector_cctor_nv_scvector_6_for_2_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
      , reg_nv_scvector_cctor_nv_scvector_6_for_2_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_6_for_2_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_2_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_6_less_14_tmp = 25'b1000000000000000000000000
      < ({nv_scvector_cctor_nv_scvector_6_for_2_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
      , reg_nv_scvector_cctor_nv_scvector_6_for_2_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_6_for_2_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_2_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_3_less_14_tmp = 26'b10000000000000000000000000
      < ({reg_nv_scvector_cctor_nv_scvector_5_for_2_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
      , reg_nv_scvector_cctor_nv_scvector_5_for_2_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_2_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_5_for_2_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_7_less_13_tmp = 26'b11000000000000000000000000
      < ({nv_scvector_cctor_nv_scvector_6_for_3_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
      , reg_nv_scvector_cctor_nv_scvector_6_for_3_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_6_for_3_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_3_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_6_less_13_tmp = 25'b1000000000000000000000000
      < ({nv_scvector_cctor_nv_scvector_6_for_3_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
      , reg_nv_scvector_cctor_nv_scvector_6_for_3_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_6_for_3_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_3_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_3_less_13_tmp = 26'b10000000000000000000000000
      < ({reg_nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
      , reg_nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_7_less_12_tmp = 26'b11000000000000000000000000
      < ({nv_scvector_cctor_nv_scvector_6_for_4_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
      , reg_nv_scvector_cctor_nv_scvector_6_for_4_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_6_for_4_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_4_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_6_less_12_tmp = 25'b1000000000000000000000000
      < ({nv_scvector_cctor_nv_scvector_6_for_4_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
      , reg_nv_scvector_cctor_nv_scvector_6_for_4_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_6_for_4_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_4_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_3_less_12_tmp = 26'b10000000000000000000000000
      < ({reg_nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
      , reg_nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_7_less_11_tmp = 26'b11000000000000000000000000
      < ({nv_scvector_cctor_nv_scvector_6_for_5_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
      , reg_nv_scvector_cctor_nv_scvector_6_for_5_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_6_for_5_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_5_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_6_less_11_tmp = 25'b1000000000000000000000000
      < ({nv_scvector_cctor_nv_scvector_6_for_5_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
      , reg_nv_scvector_cctor_nv_scvector_6_for_5_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_6_for_5_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_5_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_3_less_11_tmp = 26'b10000000000000000000000000
      < ({reg_nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
      , reg_nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_7_less_10_tmp = 26'b11000000000000000000000000
      < ({nv_scvector_cctor_nv_scvector_6_for_6_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
      , reg_nv_scvector_cctor_nv_scvector_6_for_6_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_6_for_6_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_6_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_6_less_10_tmp = 25'b1000000000000000000000000
      < ({nv_scvector_cctor_nv_scvector_6_for_6_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
      , reg_nv_scvector_cctor_nv_scvector_6_for_6_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_6_for_6_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_6_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_3_less_10_tmp = 26'b10000000000000000000000000
      < ({reg_nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
      , reg_nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_7_less_9_tmp = 26'b11000000000000000000000000
      < ({nv_scvector_cctor_nv_scvector_6_for_7_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
      , reg_nv_scvector_cctor_nv_scvector_6_for_7_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_6_for_7_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_7_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_6_less_9_tmp = 25'b1000000000000000000000000
      < ({nv_scvector_cctor_nv_scvector_6_for_7_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
      , reg_nv_scvector_cctor_nv_scvector_6_for_7_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_6_for_7_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_7_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_3_less_9_tmp = 26'b10000000000000000000000000
      < ({reg_nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
      , reg_nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_7_less_8_tmp = 26'b11000000000000000000000000
      < ({nv_scvector_cctor_nv_scvector_6_for_8_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
      , reg_nv_scvector_cctor_nv_scvector_6_for_8_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_6_for_8_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_8_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_6_less_8_tmp = 25'b1000000000000000000000000
      < ({nv_scvector_cctor_nv_scvector_6_for_8_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
      , reg_nv_scvector_cctor_nv_scvector_6_for_8_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_6_for_8_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_8_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_3_less_8_tmp = 26'b10000000000000000000000000
      < ({reg_nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
      , reg_nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_7_less_7_tmp = 26'b11000000000000000000000000
      < ({nv_scvector_cctor_nv_scvector_6_for_9_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
      , reg_nv_scvector_cctor_nv_scvector_6_for_9_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_6_for_9_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_9_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_6_less_7_tmp = 25'b1000000000000000000000000
      < ({nv_scvector_cctor_nv_scvector_6_for_9_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
      , reg_nv_scvector_cctor_nv_scvector_6_for_9_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_6_for_9_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_9_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_3_less_7_tmp = 26'b10000000000000000000000000
      < ({reg_nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
      , reg_nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_7_less_6_tmp = 26'b11000000000000000000000000
      < ({nv_scvector_cctor_nv_scvector_6_for_10_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
      , reg_nv_scvector_cctor_nv_scvector_6_for_10_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_6_for_10_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_10_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_6_less_6_tmp = 25'b1000000000000000000000000
      < ({nv_scvector_cctor_nv_scvector_6_for_10_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
      , reg_nv_scvector_cctor_nv_scvector_6_for_10_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_6_for_10_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_10_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_3_less_6_tmp = 26'b10000000000000000000000000
      < ({reg_nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
      , reg_nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_7_less_5_tmp = 26'b11000000000000000000000000
      < ({nv_scvector_cctor_nv_scvector_6_for_11_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
      , reg_nv_scvector_cctor_nv_scvector_6_for_11_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_6_for_11_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_11_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_6_less_5_tmp = 25'b1000000000000000000000000
      < ({nv_scvector_cctor_nv_scvector_6_for_11_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
      , reg_nv_scvector_cctor_nv_scvector_6_for_11_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_6_for_11_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_11_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_3_less_5_tmp = 26'b10000000000000000000000000
      < ({reg_nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
      , reg_nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_7_less_4_tmp = 26'b11000000000000000000000000
      < ({nv_scvector_cctor_nv_scvector_6_for_12_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
      , reg_nv_scvector_cctor_nv_scvector_6_for_12_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_6_for_12_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_12_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_6_less_4_tmp = 25'b1000000000000000000000000
      < ({nv_scvector_cctor_nv_scvector_6_for_12_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
      , reg_nv_scvector_cctor_nv_scvector_6_for_12_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_6_for_12_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_12_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_3_less_4_tmp = 26'b10000000000000000000000000
      < ({reg_nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
      , reg_nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_7_less_3_tmp = 26'b11000000000000000000000000
      < ({nv_scvector_cctor_nv_scvector_6_for_13_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
      , reg_nv_scvector_cctor_nv_scvector_6_for_13_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_6_for_13_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_13_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_6_less_3_tmp = 25'b1000000000000000000000000
      < ({nv_scvector_cctor_nv_scvector_6_for_13_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
      , reg_nv_scvector_cctor_nv_scvector_6_for_13_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_6_for_13_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_13_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_3_less_3_tmp = 26'b10000000000000000000000000
      < ({reg_nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
      , reg_nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_7_less_2_tmp = 26'b11000000000000000000000000
      < ({nv_scvector_cctor_nv_scvector_6_for_14_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
      , reg_nv_scvector_cctor_nv_scvector_6_for_14_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_6_for_14_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_14_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_6_less_2_tmp = 25'b1000000000000000000000000
      < ({nv_scvector_cctor_nv_scvector_6_for_14_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
      , reg_nv_scvector_cctor_nv_scvector_6_for_14_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_6_for_14_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_14_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_3_less_2_tmp = 26'b10000000000000000000000000
      < ({reg_nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
      , reg_nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_7_less_1_tmp = 26'b11000000000000000000000000
      < ({nv_scvector_cctor_nv_scvector_6_for_15_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
      , reg_nv_scvector_cctor_nv_scvector_6_for_15_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_6_for_15_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_15_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_6_less_1_tmp = 25'b1000000000000000000000000
      < ({nv_scvector_cctor_nv_scvector_6_for_15_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
      , reg_nv_scvector_cctor_nv_scvector_6_for_15_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_6_for_15_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_15_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_3_less_1_tmp = 26'b10000000000000000000000000
      < ({reg_nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
      , reg_nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_7_less_tmp = 26'b11000000000000000000000000
      < ({nv_scvector_cctor_nv_scvector_6_for_16_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
      , reg_nv_scvector_cctor_nv_scvector_6_for_16_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_6_for_16_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_16_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_6_less_tmp = 25'b1000000000000000000000000
      < ({nv_scvector_cctor_nv_scvector_6_for_16_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
      , reg_nv_scvector_cctor_nv_scvector_6_for_16_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_6_for_16_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_6_for_16_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1});
  assign operator_32_8_true_AC_TRN_AC_WRAP_3_less_tmp = 26'b10000000000000000000000000
      < ({reg_nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
      , reg_nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1});
  assign ActUnit_RunInst_switch_lp_and_48_tmp_1 = (act_config_in_InstFetch_return_sva_7_2[1:0]==2'b11)
      & act_port_PopNB_mioi_return_rsc_z_mxwt;
  assign ActUnit_RunInst_switch_lp_and_tmp_mx0w0 = Tanh_for_nor_cse_sva_mx0w0 & act_port_PopNB_mioi_return_rsc_z_mxwt;
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_8_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[31:0])
      & (signext_32_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{31{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{31{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{31{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_0_lpi_1_dfm_7 = MUX_v_32_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_8_nl,
      ({act_write_data_data_0_0_sva_31 , act_write_data_data_0_0_sva_30_26 , reg_act_write_data_data_0_0_2_ftd
      , reg_act_write_data_data_0_0_2_ftd_1 , act_write_data_data_0_0_sva_21_0}),
      while_and_1_tmp);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_9_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[63:32])
      & (signext_32_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{31{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{31{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{31{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_1_lpi_1_dfm_7 = MUX_v_32_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_9_nl,
      ({act_write_data_data_0_1_sva_31 , act_write_data_data_0_1_sva_30_26 , act_write_data_data_0_1_sva_25
      , act_write_data_data_0_1_sva_24_22 , act_write_data_data_0_1_sva_21_0}), while_and_1_tmp);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_10_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[95:64])
      & (signext_32_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{31{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{31{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{31{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_2_lpi_1_dfm_7 = MUX_v_32_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_10_nl,
      ({act_write_data_data_0_2_sva_31 , act_write_data_data_0_2_sva_30_26 , act_write_data_data_0_2_sva_25
      , act_write_data_data_0_2_sva_24_22 , act_write_data_data_0_2_sva_21_0}), while_and_1_tmp);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_11_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[127:96])
      & (signext_32_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{31{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{31{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{31{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_3_lpi_1_dfm_7 = MUX_v_32_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_11_nl,
      ({act_write_data_data_0_3_sva_31 , act_write_data_data_0_3_sva_30_26 , act_write_data_data_0_3_sva_25
      , act_write_data_data_0_3_sva_24_22 , act_write_data_data_0_3_sva_21_0}), while_and_1_tmp);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_12_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[159:128])
      & (signext_32_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{31{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{31{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{31{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_4_lpi_1_dfm_7 = MUX_v_32_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_12_nl,
      ({act_write_data_data_0_4_sva_31 , act_write_data_data_0_4_sva_30_26 , act_write_data_data_0_4_sva_25
      , act_write_data_data_0_4_sva_24_22 , act_write_data_data_0_4_sva_21_0}), while_and_1_tmp);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_13_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[191:160])
      & (signext_32_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{31{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{31{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{31{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_5_lpi_1_dfm_7 = MUX_v_32_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_13_nl,
      ({act_write_data_data_0_5_sva_31 , act_write_data_data_0_5_sva_30_26 , act_write_data_data_0_5_sva_25
      , act_write_data_data_0_5_sva_24_22 , act_write_data_data_0_5_sva_21_0}), while_and_1_tmp);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_14_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[223:192])
      & (signext_32_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{31{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{31{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{31{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_6_lpi_1_dfm_7 = MUX_v_32_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_14_nl,
      ({act_write_data_data_0_6_sva_31 , act_write_data_data_0_6_sva_30_26 , act_write_data_data_0_6_sva_25
      , act_write_data_data_0_6_sva_24_22 , act_write_data_data_0_6_sva_21_0}), while_and_1_tmp);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_15_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[255:224])
      & (signext_32_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{31{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{31{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{31{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_7_lpi_1_dfm_7 = MUX_v_32_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_15_nl,
      ({act_write_data_data_0_7_sva_31 , act_write_data_data_0_7_sva_30_26 , act_write_data_data_0_7_sva_25
      , act_write_data_data_0_7_sva_24_22 , act_write_data_data_0_7_sva_21_0}), while_and_1_tmp);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_16_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[287:256])
      & (signext_32_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{31{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{31{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{31{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_8_lpi_1_dfm_7 = MUX_v_32_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_16_nl,
      ({act_write_data_data_0_8_sva_31 , act_write_data_data_0_8_sva_30_26 , act_write_data_data_0_8_sva_25
      , act_write_data_data_0_8_sva_24_22 , act_write_data_data_0_8_sva_21_0}), while_and_1_tmp);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_17_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[319:288])
      & (signext_32_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{31{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{31{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{31{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_9_lpi_1_dfm_7 = MUX_v_32_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_17_nl,
      ({act_write_data_data_0_9_sva_31 , act_write_data_data_0_9_sva_30_26 , act_write_data_data_0_9_sva_25
      , act_write_data_data_0_9_sva_24_22 , act_write_data_data_0_9_sva_21_0}), while_and_1_tmp);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_18_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[351:320])
      & (signext_32_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{31{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{31{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{31{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_10_lpi_1_dfm_7 = MUX_v_32_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_18_nl,
      ({act_write_data_data_0_10_sva_31 , act_write_data_data_0_10_sva_30_26 , act_write_data_data_0_10_sva_25
      , act_write_data_data_0_10_sva_24_22 , act_write_data_data_0_10_sva_21_0}),
      while_and_1_tmp);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_19_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[383:352])
      & (signext_32_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{31{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{31{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{31{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_11_lpi_1_dfm_7 = MUX_v_32_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_19_nl,
      ({act_write_data_data_0_11_sva_31 , act_write_data_data_0_11_sva_30_26 , act_write_data_data_0_11_sva_25
      , act_write_data_data_0_11_sva_24_22 , act_write_data_data_0_11_sva_21_0}),
      while_and_1_tmp);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_20_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[415:384])
      & (signext_32_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{31{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{31{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{31{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_12_lpi_1_dfm_7 = MUX_v_32_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_20_nl,
      ({act_write_data_data_0_12_sva_31 , act_write_data_data_0_12_sva_30_26 , act_write_data_data_0_12_sva_25
      , act_write_data_data_0_12_sva_24_22 , act_write_data_data_0_12_sva_21_0}),
      while_and_1_tmp);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_21_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[447:416])
      & (signext_32_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{31{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{31{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{31{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_13_lpi_1_dfm_7 = MUX_v_32_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_21_nl,
      ({act_write_data_data_0_13_sva_31 , act_write_data_data_0_13_sva_30_26 , act_write_data_data_0_13_sva_25
      , act_write_data_data_0_13_sva_24_22 , act_write_data_data_0_13_sva_21_0}),
      while_and_1_tmp);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_22_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[479:448])
      & (signext_32_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{31{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{31{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{31{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign act_write_data_data_0_14_lpi_1_dfm_7 = MUX_v_32_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_22_nl,
      ({act_write_data_data_0_14_sva_31 , act_write_data_data_0_14_sva_30_26 , act_write_data_data_0_14_sva_25
      , act_write_data_data_0_14_sva_24_22 , act_write_data_data_0_14_sva_21_0}),
      while_and_1_tmp);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_23_itm = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[511:480])
      & (signext_32_1(~ ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0)) & ({{31{ActUnit_DecodeAxiRead_unequal_tmp_1}},
      ActUnit_DecodeAxiRead_unequal_tmp_1}) & ({{31{rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}},
      rva_in_PopNB_mioi_data_rw_rsc_z_mxwt}) & ({{31{rva_in_PopNB_mioi_return_rsc_z_mxwt}},
      rva_in_PopNB_mioi_return_rsc_z_mxwt});
  assign while_mux_32_nl = MUX_s_1_2_2((ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_23_itm[31]),
      act_write_data_data_0_15_sva_2_31, while_and_1_tmp);
  assign while_mux_427_nl = MUX_v_5_2_2((ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_23_itm[30:26]),
      act_write_data_data_0_15_sva_2_30_26, while_and_1_tmp);
  assign while_mux_428_nl = MUX_s_1_2_2((ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_23_itm[25]),
      reg_act_write_data_data_0_15_2_ftd, while_and_1_tmp);
  assign while_mux_430_nl = MUX_v_3_2_2((ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_23_itm[24:22]),
      reg_act_write_data_data_0_15_2_ftd_1, while_and_1_tmp);
  assign while_mux_429_nl = MUX_v_22_2_2((ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_23_itm[21:0]),
      act_write_data_data_0_15_sva_2_21_0, while_and_1_tmp);
  assign while_while_nand_nl = ~((~ ActUnit_RunInst_switch_lp_and_32_tmp) & is_start_sva);
  assign act_write_data_data_0_15_lpi_1_dfm_7 = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      ({while_mux_32_nl , while_mux_427_nl , while_mux_428_nl , while_mux_430_nl
      , while_mux_429_nl}), while_while_nand_nl);
  assign while_and_1_tmp = ActUnit_RunInst_switch_lp_and_32_tmp & is_start_sva;
  assign act_config_ActConfigRead_else_else_not_21 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7:0]==8'b00000011);
  assign while_asn_2035 = (~ while_and_88_tmp_1) | ActUnit_DecodeAxi_if_or_7_tmp_1;
  assign while_asn_2037 = (~(act_config_ActConfigRead_unequal_tmp_1 | ActUnit_DecodeAxi_if_or_7_tmp_1))
      & while_and_88_tmp_1;
  assign while_asn_2039 = act_config_ActConfigRead_unequal_tmp_1 & (~ ActUnit_DecodeAxi_if_or_7_tmp_1)
      & while_and_88_tmp_1;
  assign nl_Silu_for_y_1_sva_1_22_0_1 = ({1'b1 , (Silu_for_1_else_if_Silu_for_else_if_mul_cmp_z[43:22])})
      + 23'b00110011001100110011001;
  assign Silu_for_y_1_sva_1_22_0_1 = nl_Silu_for_y_1_sva_1_22_0_1[22:0];
  assign Silu_for_else_and_ssc_1 = (~ Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign Silu_for_else_else_else_and_1_ssc_1 = Gelu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
      & Gelu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Silu_for_else_and_1_m1c_mx1;
  assign nl_Silu_for_y_2_sva_1_22_0_1 = ({1'b1 , (Silu_for_1_else_if_Silu_for_else_if_mul_cmp_7_z[43:22])})
      + 23'b00110011001100110011001;
  assign Silu_for_y_2_sva_1_22_0_1 = nl_Silu_for_y_2_sva_1_22_0_1[22:0];
  assign Silu_for_else_and_2_ssc_1 = (~ Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign Silu_for_else_else_else_and_3_ssc_1 = Gelu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
      & Gelu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Silu_for_else_and_3_m1c_mx1;
  assign nl_Silu_for_y_3_sva_1_22_0_1 = ({1'b1 , (Silu_for_1_else_if_Silu_for_else_if_mul_cmp_6_z[43:22])})
      + 23'b00110011001100110011001;
  assign Silu_for_y_3_sva_1_22_0_1 = nl_Silu_for_y_3_sva_1_22_0_1[22:0];
  assign Silu_for_else_and_4_ssc_1 = (~ Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign Silu_for_else_else_else_and_5_ssc_1 = Gelu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
      & Gelu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Silu_for_else_and_5_m1c_mx1;
  assign nl_Silu_for_y_4_sva_1_22_0_1 = ({1'b1 , (Silu_for_1_else_if_Silu_for_else_if_mul_cmp_5_z[43:22])})
      + 23'b00110011001100110011001;
  assign Silu_for_y_4_sva_1_22_0_1 = nl_Silu_for_y_4_sva_1_22_0_1[22:0];
  assign Silu_for_else_and_6_ssc_1 = (~ Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign Silu_for_else_else_else_and_7_ssc_1 = Gelu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
      & Gelu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Silu_for_else_and_7_m1c_mx1;
  assign nl_Silu_for_y_5_sva_1_22_0_1 = ({1'b1 , (Silu_for_1_else_if_Silu_for_else_if_mul_cmp_4_z[43:22])})
      + 23'b00110011001100110011001;
  assign Silu_for_y_5_sva_1_22_0_1 = nl_Silu_for_y_5_sva_1_22_0_1[22:0];
  assign Silu_for_else_and_8_ssc_1 = (~ Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign Silu_for_else_else_else_and_9_ssc_1 = Gelu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
      & Gelu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Silu_for_else_and_9_m1c_mx1;
  assign nl_Silu_for_y_6_sva_1_22_0_1 = ({1'b1 , (Silu_for_1_else_if_Silu_for_else_if_mul_cmp_3_z[43:22])})
      + 23'b00110011001100110011001;
  assign Silu_for_y_6_sva_1_22_0_1 = nl_Silu_for_y_6_sva_1_22_0_1[22:0];
  assign Silu_for_else_and_10_ssc_1 = (~ Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign Silu_for_else_else_else_and_11_ssc_1 = Gelu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
      & Gelu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Silu_for_else_and_11_m1c_mx1;
  assign nl_Silu_for_y_7_sva_1_22_0_1 = ({1'b1 , (Silu_for_1_else_if_Silu_for_else_if_mul_cmp_2_z[43:22])})
      + 23'b00110011001100110011001;
  assign Silu_for_y_7_sva_1_22_0_1 = nl_Silu_for_y_7_sva_1_22_0_1[22:0];
  assign Silu_for_else_and_12_ssc_1 = (~ Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign Silu_for_else_else_else_and_13_ssc_1 = Gelu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
      & Gelu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Silu_for_else_and_13_m1c_mx1;
  assign nl_Silu_for_y_8_sva_1_22_0_1 = ({1'b1 , (Silu_for_1_else_if_Silu_for_else_if_mul_cmp_1_z[43:22])})
      + 23'b00110011001100110011001;
  assign Silu_for_y_8_sva_1_22_0_1 = nl_Silu_for_y_8_sva_1_22_0_1[22:0];
  assign Silu_for_else_and_14_ssc_1 = (~ Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign Silu_for_else_else_else_and_15_ssc_1 = Gelu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
      & Gelu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Silu_for_else_and_15_m1c_mx1;
  assign Silu_for_else_and_39_ssc_1 = (~ Gelu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs)
      & Silu_for_else_and_15_m1c_mx1;
  assign Silu_for_else_else_else_and_14_ssc_1 = (~ Gelu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      & Gelu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Silu_for_else_and_15_m1c_mx1;
  assign Silu_for_else_and_38_ssc_1 = (~ Gelu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs)
      & Silu_for_else_and_13_m1c_mx1;
  assign Silu_for_else_else_else_and_12_ssc_1 = (~ Gelu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      & Gelu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Silu_for_else_and_13_m1c_mx1;
  assign Silu_for_else_and_37_ssc_1 = (~ Gelu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs)
      & Silu_for_else_and_11_m1c_mx1;
  assign Silu_for_else_else_else_and_10_ssc_1 = (~ Gelu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      & Gelu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Silu_for_else_and_11_m1c_mx1;
  assign Silu_for_else_and_36_ssc_1 = (~ Gelu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs)
      & Silu_for_else_and_9_m1c_mx1;
  assign Silu_for_else_else_else_and_8_ssc_1 = (~ Gelu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      & Gelu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Silu_for_else_and_9_m1c_mx1;
  assign Silu_for_else_and_35_ssc_1 = (~ Gelu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs)
      & Silu_for_else_and_7_m1c_mx1;
  assign Silu_for_else_else_else_and_6_ssc_1 = (~ Gelu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      & Gelu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Silu_for_else_and_7_m1c_mx1;
  assign Silu_for_else_and_34_ssc_1 = (~ Gelu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs)
      & Silu_for_else_and_5_m1c_mx1;
  assign Silu_for_else_else_else_and_4_ssc_1 = (~ Gelu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      & Gelu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Silu_for_else_and_5_m1c_mx1;
  assign Silu_for_else_and_33_ssc_1 = (~ Gelu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs)
      & Silu_for_else_and_3_m1c_mx1;
  assign Silu_for_else_else_else_and_2_ssc_1 = (~ Gelu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      & Gelu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Silu_for_else_and_3_m1c_mx1;
  assign Silu_for_else_and_32_ssc_1 = (~ Gelu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs)
      & Silu_for_else_and_1_m1c_mx1;
  assign Silu_for_else_else_else_and_ssc_1 = (~ Gelu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      & Gelu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Silu_for_else_and_1_m1c_mx1;
  assign ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_21_0_mx0w1
      = MUX_v_22_64_2(act_regs_data_0_0_sva_dfm_2_21_0, act_regs_data_0_1_sva_dfm_2_21_0,
      act_regs_data_0_2_sva_dfm_2_21_0, act_regs_data_0_3_sva_dfm_2_21_0, act_regs_data_0_4_sva_dfm_2_21_0,
      act_regs_data_0_5_sva_dfm_2_21_0, act_regs_data_0_6_sva_dfm_2_21_0, act_regs_data_0_7_sva_dfm_2_21_0,
      act_regs_data_0_8_sva_dfm_2_21_0, act_regs_data_0_9_sva_dfm_2_21_0, act_regs_data_0_10_sva_dfm_2_21_0,
      act_regs_data_0_11_sva_dfm_2_21_0, act_regs_data_0_12_sva_dfm_2_21_0, act_regs_data_0_13_sva_dfm_2_21_0,
      act_regs_data_0_14_sva_dfm_2_21_0, act_regs_data_0_15_sva_dfm_2_21_0, act_regs_data_1_0_sva_dfm_2_21_0,
      act_regs_data_1_1_sva_dfm_2_21_0, act_regs_data_1_2_sva_dfm_2_21_0, act_regs_data_1_3_sva_dfm_2_21_0,
      act_regs_data_1_4_sva_dfm_2_21_0, act_regs_data_1_5_sva_dfm_2_21_0, act_regs_data_1_6_sva_dfm_2_21_0,
      act_regs_data_1_7_sva_dfm_2_21_0, act_regs_data_1_8_sva_dfm_2_21_0, act_regs_data_1_9_sva_dfm_2_21_0,
      act_regs_data_1_10_sva_dfm_2_21_0, act_regs_data_1_11_sva_dfm_2_21_0, act_regs_data_1_12_sva_dfm_2_21_0,
      act_regs_data_1_13_sva_dfm_2_21_0, act_regs_data_1_14_sva_dfm_2_21_0, act_regs_data_1_15_sva_dfm_2_21_0,
      act_regs_data_2_0_sva_dfm_2_21_0, act_regs_data_2_1_sva_dfm_2_21_0, act_regs_data_2_2_sva_dfm_2_21_0,
      act_regs_data_2_3_sva_dfm_2_21_0, act_regs_data_2_4_sva_dfm_2_21_0, act_regs_data_2_5_sva_dfm_2_21_0,
      act_regs_data_2_6_sva_dfm_2_21_0, act_regs_data_2_7_sva_dfm_2_21_0, act_regs_data_2_8_sva_dfm_2_21_0,
      act_regs_data_2_9_sva_dfm_2_21_0, act_regs_data_2_10_sva_dfm_2_21_0, act_regs_data_2_11_sva_dfm_2_21_0,
      act_regs_data_2_12_sva_dfm_2_21_0, act_regs_data_2_13_sva_dfm_2_21_0, act_regs_data_2_14_sva_dfm_2_21_0,
      act_regs_data_2_15_sva_dfm_2_21_0, act_regs_data_3_0_sva_dfm_2_21_0, act_regs_data_3_1_sva_dfm_2_21_0,
      act_regs_data_3_2_sva_dfm_2_21_0, act_regs_data_3_3_sva_dfm_2_21_0, act_regs_data_3_4_sva_dfm_2_21_0,
      act_regs_data_3_5_sva_dfm_2_21_0, act_regs_data_3_6_sva_dfm_2_21_0, act_regs_data_3_7_sva_dfm_2_21_0,
      act_regs_data_3_8_sva_dfm_2_21_0, act_regs_data_3_9_sva_dfm_2_21_0, act_regs_data_3_10_sva_dfm_2_21_0,
      act_regs_data_3_11_sva_dfm_2_21_0, act_regs_data_3_12_sva_dfm_2_21_0, act_regs_data_3_13_sva_dfm_2_21_0,
      act_regs_data_3_14_sva_dfm_2_21_0, act_regs_data_3_15_sva_dfm_2_21_0, {nvhls_get_slc_2U_NVUINT8_return_2_sva
      , ActUnit_PushOutput_if_for_i_4_0_sva_3_0});
  assign Silu_for_else_mux_40_nl = MUX_s_1_2_2((Silu_for_y_1_sva_1_22_0_1[22]), (Silu_for_16_else_else_if_acc_itm[1]),
      Silu_for_else_and_30_ssc_1);
  assign Silu_for_y_lpi_1_dfm_4_31_1 = Silu_for_else_mux_40_nl & (~(Silu_for_else_and_47_ssc_1
      | Silu_for_else_else_else_and_30_ssc_1 | Silu_for_else_else_else_and_31_ssc_1))
      & Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  assign Silu_for_else_or_15_itm = Silu_for_else_else_else_and_30_ssc_1 | Silu_for_else_else_else_and_31_ssc_1;
  assign Silu_for_else_Silu_for_else_mux1h_47_nl = MUX1HOT_v_2_4_2((Silu_for_y_1_sva_1_22_0_1[21:20]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1[1:0]),
      (reg_Silu_for_16_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1[21:20]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:20]),
      {(~ Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_30_ssc_1 , Silu_for_else_and_47_ssc_1 , Silu_for_else_or_15_itm});
  assign Silu_for_else_Silu_for_else_mux1h_64_nl = MUX1HOT_v_20_4_2((Silu_for_y_1_sva_1_22_0_1[19:0]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:2]),
      (reg_Silu_for_16_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1[19:0]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[19:0]),
      {(~ Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_30_ssc_1 , Silu_for_else_and_47_ssc_1 , Silu_for_else_or_15_itm});
  assign Silu_for_y_lpi_1_dfm_4_21_0_1 = MUX_v_22_2_2(22'b0000000000000000000000,
      ({Silu_for_else_Silu_for_else_mux1h_47_nl , Silu_for_else_Silu_for_else_mux1h_64_nl}),
      Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
  assign Silu_for_else_Silu_for_else_mux1h_15_nl = MUX1HOT_v_5_3_2((signext_5_1(Silu_for_y_1_sva_1_22_0_1[22])),
      (signext_5_1(Silu_for_16_else_else_if_acc_itm[1])), reg_nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26,
      {(~ Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_30_ssc_1 , Silu_for_else_else_else_and_31_ssc_1});
  assign Silu_for_else_nor_31_nl = ~(Silu_for_else_and_47_ssc_1 | Silu_for_else_else_else_and_30_ssc_1);
  assign Silu_for_y_lpi_1_dfm_4_30_26_1 = Silu_for_else_Silu_for_else_mux1h_15_nl
      & (signext_5_1(Silu_for_else_nor_31_nl)) & ({{4{Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs}},
      Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs});
  assign Silu_for_else_mux_41_nl = MUX_s_1_2_2((Silu_for_y_8_sva_1_22_0_1[22]), (Silu_for_15_else_else_if_acc_itm[1]),
      Silu_for_else_and_28_ssc_1);
  assign Silu_for_y_15_lpi_1_dfm_4_31_1 = Silu_for_else_mux_41_nl & (~(Silu_for_else_and_46_ssc_1
      | Silu_for_else_else_else_and_28_ssc_1 | Silu_for_else_else_else_and_29_ssc_1))
      & Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  assign Silu_for_else_or_14_itm = Silu_for_else_else_else_and_28_ssc_1 | Silu_for_else_else_else_and_29_ssc_1;
  assign Silu_for_else_Silu_for_else_mux1h_46_nl = MUX1HOT_v_2_4_2((Silu_for_y_8_sva_1_22_0_1[21:20]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1[1:0]),
      (reg_Silu_for_15_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1[21:20]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:20]),
      {(~ Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_28_ssc_1 , Silu_for_else_and_46_ssc_1 , Silu_for_else_or_14_itm});
  assign Silu_for_else_Silu_for_else_mux1h_66_nl = MUX1HOT_v_20_4_2((Silu_for_y_8_sva_1_22_0_1[19:0]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:2]),
      (reg_Silu_for_15_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1[19:0]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[19:0]),
      {(~ Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_28_ssc_1 , Silu_for_else_and_46_ssc_1 , Silu_for_else_or_14_itm});
  assign Silu_for_y_15_lpi_1_dfm_4_21_0_1 = MUX_v_22_2_2(22'b0000000000000000000000,
      ({Silu_for_else_Silu_for_else_mux1h_46_nl , Silu_for_else_Silu_for_else_mux1h_66_nl}),
      Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
  assign Silu_for_else_Silu_for_else_mux1h_14_nl = MUX1HOT_v_5_3_2((signext_5_1(Silu_for_y_8_sva_1_22_0_1[22])),
      (signext_5_1(Silu_for_15_else_else_if_acc_itm[1])), reg_nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26,
      {(~ Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_28_ssc_1 , Silu_for_else_else_else_and_29_ssc_1});
  assign Silu_for_else_nor_29_nl = ~(Silu_for_else_and_46_ssc_1 | Silu_for_else_else_else_and_28_ssc_1);
  assign Silu_for_y_15_lpi_1_dfm_4_30_26_1 = Silu_for_else_Silu_for_else_mux1h_14_nl
      & (signext_5_1(Silu_for_else_nor_29_nl)) & ({{4{Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs}},
      Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs});
  assign Silu_for_else_mux_42_nl = MUX_s_1_2_2((Silu_for_y_7_sva_1_22_0_1[22]), (Silu_for_14_else_else_if_acc_itm[1]),
      Silu_for_else_and_26_ssc_1);
  assign Silu_for_y_14_lpi_1_dfm_4_31_1 = Silu_for_else_mux_42_nl & (~(Silu_for_else_and_45_ssc_1
      | Silu_for_else_else_else_and_26_ssc_1 | Silu_for_else_else_else_and_27_ssc_1))
      & Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  assign Silu_for_else_or_13_itm = Silu_for_else_else_else_and_26_ssc_1 | Silu_for_else_else_else_and_27_ssc_1;
  assign Silu_for_else_Silu_for_else_mux1h_45_nl = MUX1HOT_v_2_4_2((Silu_for_y_7_sva_1_22_0_1[21:20]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1[1:0]),
      (reg_Silu_for_14_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1[21:20]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:20]),
      {(~ Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_26_ssc_1 , Silu_for_else_and_45_ssc_1 , Silu_for_else_or_13_itm});
  assign Silu_for_else_Silu_for_else_mux1h_68_nl = MUX1HOT_v_20_4_2((Silu_for_y_7_sva_1_22_0_1[19:0]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:2]),
      (reg_Silu_for_14_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1[19:0]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[19:0]),
      {(~ Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_26_ssc_1 , Silu_for_else_and_45_ssc_1 , Silu_for_else_or_13_itm});
  assign Silu_for_y_14_lpi_1_dfm_4_21_0_1 = MUX_v_22_2_2(22'b0000000000000000000000,
      ({Silu_for_else_Silu_for_else_mux1h_45_nl , Silu_for_else_Silu_for_else_mux1h_68_nl}),
      Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
  assign Silu_for_else_Silu_for_else_mux1h_13_nl = MUX1HOT_v_5_3_2((signext_5_1(Silu_for_y_7_sva_1_22_0_1[22])),
      (signext_5_1(Silu_for_14_else_else_if_acc_itm[1])), reg_nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26,
      {(~ Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_26_ssc_1 , Silu_for_else_else_else_and_27_ssc_1});
  assign Silu_for_else_nor_27_nl = ~(Silu_for_else_and_45_ssc_1 | Silu_for_else_else_else_and_26_ssc_1);
  assign Silu_for_y_14_lpi_1_dfm_4_30_26_1 = Silu_for_else_Silu_for_else_mux1h_13_nl
      & (signext_5_1(Silu_for_else_nor_27_nl)) & ({{4{Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs}},
      Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs});
  assign Silu_for_else_mux_43_nl = MUX_s_1_2_2((Silu_for_y_6_sva_1_22_0_1[22]), (Silu_for_13_else_else_if_acc_itm[1]),
      Silu_for_else_and_24_ssc_1);
  assign Silu_for_y_13_lpi_1_dfm_4_31_1 = Silu_for_else_mux_43_nl & (~(Silu_for_else_and_44_ssc_1
      | Silu_for_else_else_else_and_24_ssc_1 | Silu_for_else_else_else_and_25_ssc_1))
      & Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  assign Silu_for_else_or_12_itm = Silu_for_else_else_else_and_24_ssc_1 | Silu_for_else_else_else_and_25_ssc_1;
  assign Silu_for_else_Silu_for_else_mux1h_44_nl = MUX1HOT_v_2_4_2((Silu_for_y_6_sva_1_22_0_1[21:20]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1[1:0]),
      (reg_Silu_for_13_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1[21:20]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:20]),
      {(~ Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_24_ssc_1 , Silu_for_else_and_44_ssc_1 , Silu_for_else_or_12_itm});
  assign Silu_for_else_Silu_for_else_mux1h_70_nl = MUX1HOT_v_20_4_2((Silu_for_y_6_sva_1_22_0_1[19:0]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:2]),
      (reg_Silu_for_13_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1[19:0]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[19:0]),
      {(~ Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_24_ssc_1 , Silu_for_else_and_44_ssc_1 , Silu_for_else_or_12_itm});
  assign Silu_for_y_13_lpi_1_dfm_4_21_0_1 = MUX_v_22_2_2(22'b0000000000000000000000,
      ({Silu_for_else_Silu_for_else_mux1h_44_nl , Silu_for_else_Silu_for_else_mux1h_70_nl}),
      Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
  assign Silu_for_else_Silu_for_else_mux1h_12_nl = MUX1HOT_v_5_3_2((signext_5_1(Silu_for_y_6_sva_1_22_0_1[22])),
      (signext_5_1(Silu_for_13_else_else_if_acc_itm[1])), reg_nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26,
      {(~ Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_24_ssc_1 , Silu_for_else_else_else_and_25_ssc_1});
  assign Silu_for_else_nor_25_nl = ~(Silu_for_else_and_44_ssc_1 | Silu_for_else_else_else_and_24_ssc_1);
  assign Silu_for_y_13_lpi_1_dfm_4_30_26_1 = Silu_for_else_Silu_for_else_mux1h_12_nl
      & (signext_5_1(Silu_for_else_nor_25_nl)) & ({{4{Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs}},
      Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs});
  assign Silu_for_else_mux_44_nl = MUX_s_1_2_2((Silu_for_y_5_sva_1_22_0_1[22]), (Silu_for_12_else_else_if_acc_itm[1]),
      Silu_for_else_and_22_ssc_1);
  assign Silu_for_y_12_lpi_1_dfm_4_31_1 = Silu_for_else_mux_44_nl & (~(Silu_for_else_and_43_ssc_1
      | Silu_for_else_else_else_and_22_ssc_1 | Silu_for_else_else_else_and_23_ssc_1))
      & Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  assign Silu_for_else_or_11_itm = Silu_for_else_else_else_and_22_ssc_1 | Silu_for_else_else_else_and_23_ssc_1;
  assign Silu_for_else_Silu_for_else_mux1h_43_nl = MUX1HOT_v_2_4_2((Silu_for_y_5_sva_1_22_0_1[21:20]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1[1:0]),
      (reg_Silu_for_12_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1[21:20]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:20]),
      {(~ Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_22_ssc_1 , Silu_for_else_and_43_ssc_1 , Silu_for_else_or_11_itm});
  assign Silu_for_else_Silu_for_else_mux1h_72_nl = MUX1HOT_v_20_4_2((Silu_for_y_5_sva_1_22_0_1[19:0]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:2]),
      (reg_Silu_for_12_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1[19:0]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[19:0]),
      {(~ Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_22_ssc_1 , Silu_for_else_and_43_ssc_1 , Silu_for_else_or_11_itm});
  assign Silu_for_y_12_lpi_1_dfm_4_21_0_1 = MUX_v_22_2_2(22'b0000000000000000000000,
      ({Silu_for_else_Silu_for_else_mux1h_43_nl , Silu_for_else_Silu_for_else_mux1h_72_nl}),
      Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
  assign Silu_for_else_Silu_for_else_mux1h_11_nl = MUX1HOT_v_5_3_2((signext_5_1(Silu_for_y_5_sva_1_22_0_1[22])),
      (signext_5_1(Silu_for_12_else_else_if_acc_itm[1])), reg_nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26,
      {(~ Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_22_ssc_1 , Silu_for_else_else_else_and_23_ssc_1});
  assign Silu_for_else_nor_23_nl = ~(Silu_for_else_and_43_ssc_1 | Silu_for_else_else_else_and_22_ssc_1);
  assign Silu_for_y_12_lpi_1_dfm_4_30_26_1 = Silu_for_else_Silu_for_else_mux1h_11_nl
      & (signext_5_1(Silu_for_else_nor_23_nl)) & ({{4{Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs}},
      Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs});
  assign Silu_for_else_mux_45_nl = MUX_s_1_2_2((Silu_for_y_4_sva_1_22_0_1[22]), (Silu_for_11_else_else_if_acc_itm[1]),
      Silu_for_else_and_20_ssc_1);
  assign Silu_for_y_11_lpi_1_dfm_4_31_1 = Silu_for_else_mux_45_nl & (~(Silu_for_else_and_42_ssc_1
      | Silu_for_else_else_else_and_20_ssc_1 | Silu_for_else_else_else_and_21_ssc_1))
      & Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  assign Silu_for_else_or_10_itm = Silu_for_else_else_else_and_20_ssc_1 | Silu_for_else_else_else_and_21_ssc_1;
  assign Silu_for_else_Silu_for_else_mux1h_42_nl = MUX1HOT_v_2_4_2((Silu_for_y_4_sva_1_22_0_1[21:20]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1[1:0]),
      (reg_Silu_for_11_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1[21:20]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:20]),
      {(~ Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_20_ssc_1 , Silu_for_else_and_42_ssc_1 , Silu_for_else_or_10_itm});
  assign Silu_for_else_Silu_for_else_mux1h_74_nl = MUX1HOT_v_20_4_2((Silu_for_y_4_sva_1_22_0_1[19:0]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:2]),
      (reg_Silu_for_11_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1[19:0]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[19:0]),
      {(~ Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_20_ssc_1 , Silu_for_else_and_42_ssc_1 , Silu_for_else_or_10_itm});
  assign Silu_for_y_11_lpi_1_dfm_4_21_0_1 = MUX_v_22_2_2(22'b0000000000000000000000,
      ({Silu_for_else_Silu_for_else_mux1h_42_nl , Silu_for_else_Silu_for_else_mux1h_74_nl}),
      Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
  assign Silu_for_else_Silu_for_else_mux1h_10_nl = MUX1HOT_v_5_3_2((signext_5_1(Silu_for_y_4_sva_1_22_0_1[22])),
      (signext_5_1(Silu_for_11_else_else_if_acc_itm[1])), reg_nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26,
      {(~ Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_20_ssc_1 , Silu_for_else_else_else_and_21_ssc_1});
  assign Silu_for_else_nor_21_nl = ~(Silu_for_else_and_42_ssc_1 | Silu_for_else_else_else_and_20_ssc_1);
  assign Silu_for_y_11_lpi_1_dfm_4_30_26_1 = Silu_for_else_Silu_for_else_mux1h_10_nl
      & (signext_5_1(Silu_for_else_nor_21_nl)) & ({{4{Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs}},
      Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs});
  assign Silu_for_else_mux_46_nl = MUX_s_1_2_2((Silu_for_y_3_sva_1_22_0_1[22]), (Silu_for_10_else_else_if_acc_itm[1]),
      Silu_for_else_and_18_ssc_1);
  assign Silu_for_y_10_lpi_1_dfm_4_31_1 = Silu_for_else_mux_46_nl & (~(Silu_for_else_and_41_ssc_1
      | Silu_for_else_else_else_and_18_ssc_1 | Silu_for_else_else_else_and_19_ssc_1))
      & Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  assign Silu_for_else_or_9_itm = Silu_for_else_else_else_and_18_ssc_1 | Silu_for_else_else_else_and_19_ssc_1;
  assign Silu_for_else_Silu_for_else_mux1h_41_nl = MUX1HOT_v_2_4_2((Silu_for_y_3_sva_1_22_0_1[21:20]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1[1:0]),
      (reg_Silu_for_10_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1[21:20]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:20]),
      {(~ Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_18_ssc_1 , Silu_for_else_and_41_ssc_1 , Silu_for_else_or_9_itm});
  assign Silu_for_else_Silu_for_else_mux1h_76_nl = MUX1HOT_v_20_4_2((Silu_for_y_3_sva_1_22_0_1[19:0]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:2]),
      (reg_Silu_for_10_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1[19:0]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[19:0]),
      {(~ Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_18_ssc_1 , Silu_for_else_and_41_ssc_1 , Silu_for_else_or_9_itm});
  assign Silu_for_y_10_lpi_1_dfm_4_21_0_1 = MUX_v_22_2_2(22'b0000000000000000000000,
      ({Silu_for_else_Silu_for_else_mux1h_41_nl , Silu_for_else_Silu_for_else_mux1h_76_nl}),
      Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
  assign Silu_for_else_Silu_for_else_mux1h_9_nl = MUX1HOT_v_5_3_2((signext_5_1(Silu_for_y_3_sva_1_22_0_1[22])),
      (signext_5_1(Silu_for_10_else_else_if_acc_itm[1])), reg_nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26,
      {(~ Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_18_ssc_1 , Silu_for_else_else_else_and_19_ssc_1});
  assign Silu_for_else_nor_19_nl = ~(Silu_for_else_and_41_ssc_1 | Silu_for_else_else_else_and_18_ssc_1);
  assign Silu_for_y_10_lpi_1_dfm_4_30_26_1 = Silu_for_else_Silu_for_else_mux1h_9_nl
      & (signext_5_1(Silu_for_else_nor_19_nl)) & ({{4{Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs}},
      Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs});
  assign Silu_for_else_mux_47_nl = MUX_s_1_2_2((Silu_for_y_2_sva_1_22_0_1[22]), (Silu_for_9_else_else_if_acc_itm[1]),
      Silu_for_else_and_16_ssc_1);
  assign Silu_for_y_9_lpi_1_dfm_4_31_1 = Silu_for_else_mux_47_nl & (~(Silu_for_else_and_40_ssc_1
      | Silu_for_else_else_else_and_16_ssc_1 | Silu_for_else_else_else_and_17_ssc_1))
      & Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  assign Silu_for_else_or_8_itm = Silu_for_else_else_else_and_16_ssc_1 | Silu_for_else_else_else_and_17_ssc_1;
  assign Silu_for_else_Silu_for_else_mux1h_40_nl = MUX1HOT_v_2_4_2((Silu_for_y_2_sva_1_22_0_1[21:20]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1[1:0]),
      (Silu_for_9_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0[21:20]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:20]),
      {(~ Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_16_ssc_1 , Silu_for_else_and_40_ssc_1 , Silu_for_else_or_8_itm});
  assign Silu_for_else_Silu_for_else_mux1h_78_nl = MUX1HOT_v_20_4_2((Silu_for_y_2_sva_1_22_0_1[19:0]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:2]),
      (Silu_for_9_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0[19:0]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[19:0]),
      {(~ Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_16_ssc_1 , Silu_for_else_and_40_ssc_1 , Silu_for_else_or_8_itm});
  assign Silu_for_y_9_lpi_1_dfm_4_21_0_1 = MUX_v_22_2_2(22'b0000000000000000000000,
      ({Silu_for_else_Silu_for_else_mux1h_40_nl , Silu_for_else_Silu_for_else_mux1h_78_nl}),
      Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
  assign Silu_for_else_Silu_for_else_mux1h_8_nl = MUX1HOT_v_5_3_2((signext_5_1(Silu_for_y_2_sva_1_22_0_1[22])),
      (signext_5_1(Silu_for_9_else_else_if_acc_itm[1])), reg_nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26,
      {(~ Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_16_ssc_1 , Silu_for_else_else_else_and_17_ssc_1});
  assign Silu_for_else_nor_17_nl = ~(Silu_for_else_and_40_ssc_1 | Silu_for_else_else_else_and_16_ssc_1);
  assign Silu_for_y_9_lpi_1_dfm_4_30_26_1 = Silu_for_else_Silu_for_else_mux1h_8_nl
      & (signext_5_1(Silu_for_else_nor_17_nl)) & ({{4{Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs}},
      Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs});
  assign Gelu_for_else_Gelu_for_else_mux1h_15_nl = MUX1HOT_s_1_3_2((Gelu_for_2_else_if_acc_itm_mx1w0[3]),
      (Gelu_for_1_else_else_if_mul_cmp_1_z[46]), (Gelu_for_y_sva_4_27_22_1[5]), {(~
      Gelu_for_16_else_slc_32_svs) , Gelu_for_else_and_30_ssc_1 , Gelu_for_else_else_else_and_30_ssc_1});
  assign Gelu_for_y_lpi_1_dfm_4_31_1 = Gelu_for_else_Gelu_for_else_mux1h_15_nl &
      (~(Gelu_for_else_and_47_ssc_1 | Gelu_for_else_else_else_and_31_ssc_1)) & Gelu_for_16_slc_32_1_svs;
  assign Gelu_for_else_or_nl = Gelu_for_else_and_47_ssc_1 | Gelu_for_else_else_else_and_30_ssc_1;
  assign Gelu_for_else_Gelu_for_else_mux1h_47_nl = MUX1HOT_v_22_4_2((Silu_for_1_else_if_Silu_for_else_if_mul_cmp_z[44:23]),
      (Gelu_for_1_else_else_if_mul_cmp_1_z[45:24]), (Gelu_for_1_else_else_else_if_mul_cmp_1_z[45:24]),
      act_write_data_data_0_15_sva_2_21_0, {(~ Gelu_for_16_else_slc_32_svs) , Gelu_for_else_and_30_ssc_1
      , Gelu_for_else_or_nl , Gelu_for_else_else_else_and_31_ssc_1});
  assign Gelu_for_y_lpi_1_dfm_4_21_0_1 = MUX_v_22_2_2(22'b0000000000000000000000,
      Gelu_for_else_Gelu_for_else_mux1h_47_nl, Gelu_for_16_slc_32_1_svs);
  assign Gelu_for_else_Gelu_for_else_mux1h_31_nl = MUX1HOT_v_5_4_2((signext_5_1(Gelu_for_2_else_if_acc_itm_mx1w0[3])),
      (signext_5_1(Gelu_for_1_else_else_if_mul_cmp_1_z[46])), (signext_5_2(Gelu_for_y_sva_4_27_22_1[5:4])),
      act_write_data_data_0_15_sva_2_30_26, {(~ Gelu_for_16_else_slc_32_svs) , Gelu_for_else_and_30_ssc_1
      , Gelu_for_else_else_else_and_30_ssc_1 , Gelu_for_else_else_else_and_31_ssc_1});
  assign Gelu_for_y_lpi_1_dfm_4_30_26 = Gelu_for_else_Gelu_for_else_mux1h_31_nl &
      (signext_5_1(~ Gelu_for_else_and_47_ssc_1)) & ({{4{Gelu_for_16_slc_32_1_svs}},
      Gelu_for_16_slc_32_1_svs});
  assign Gelu_for_else_Gelu_for_else_mux1h_63_nl = MUX1HOT_s_1_4_2((Gelu_for_2_else_if_acc_itm_mx1w0[3]),
      (Gelu_for_1_else_else_if_mul_cmp_1_z[46]), (Gelu_for_y_sva_4_27_22_1[3]), reg_act_write_data_data_0_15_2_ftd,
      {(~ Gelu_for_16_else_slc_32_svs) , Gelu_for_else_and_30_ssc_1 , Gelu_for_else_else_else_and_30_ssc_1
      , Gelu_for_else_else_else_and_31_ssc_1});
  assign Gelu_for_y_lpi_1_dfm_4_25 = Gelu_for_else_Gelu_for_else_mux1h_63_nl & (~
      Gelu_for_else_and_47_ssc_1) & Gelu_for_16_slc_32_1_svs;
  assign Gelu_for_else_Gelu_for_else_mux1h_79_nl = MUX1HOT_v_3_5_2((Gelu_for_2_else_if_acc_itm_mx1w0[2:0]),
      (signext_3_1(Gelu_for_1_else_else_if_mul_cmp_1_z[46])), (Gelu_for_1_else_else_else_if_mul_cmp_1_z[48:46]),
      (Gelu_for_y_sva_4_27_22_1[2:0]), reg_act_write_data_data_0_15_2_ftd_1, {(~
      Gelu_for_16_else_slc_32_svs) , Gelu_for_else_and_30_ssc_1 , Gelu_for_else_and_47_ssc_1
      , Gelu_for_else_else_else_and_30_ssc_1 , Gelu_for_else_else_else_and_31_ssc_1});
  assign Gelu_for_y_lpi_1_dfm_4_24_22 = MUX_v_3_2_2(3'b000, Gelu_for_else_Gelu_for_else_mux1h_79_nl,
      Gelu_for_16_slc_32_1_svs);
  assign Gelu_for_else_Gelu_for_else_mux1h_14_nl = MUX1HOT_s_1_3_2((Gelu_for_8_else_if_acc_itm_mx1w0[3]),
      (Gelu_for_1_else_else_if_mul_cmp_2_z[46]), (Gelu_for_y_15_sva_4_27_22_1[5]),
      {(~ Gelu_for_15_else_slc_32_svs) , Gelu_for_else_and_28_ssc_1 , Gelu_for_else_else_else_and_28_ssc_1});
  assign Gelu_for_y_15_lpi_1_dfm_4_31_1 = Gelu_for_else_Gelu_for_else_mux1h_14_nl
      & (~(Gelu_for_else_and_46_ssc_1 | Gelu_for_else_else_else_and_29_ssc_1)) &
      Gelu_for_15_slc_32_1_svs;
  assign Gelu_for_else_or_1_nl = Gelu_for_else_and_46_ssc_1 | Gelu_for_else_else_else_and_28_ssc_1;
  assign Gelu_for_else_Gelu_for_else_mux1h_46_nl = MUX1HOT_v_22_4_2((Silu_for_1_else_if_Silu_for_else_if_mul_cmp_1_z[44:23]),
      (Gelu_for_1_else_else_if_mul_cmp_2_z[45:24]), (Gelu_for_1_else_else_else_if_mul_cmp_2_z[45:24]),
      act_write_data_data_0_14_sva_21_0, {(~ Gelu_for_15_else_slc_32_svs) , Gelu_for_else_and_28_ssc_1
      , Gelu_for_else_or_1_nl , Gelu_for_else_else_else_and_29_ssc_1});
  assign Gelu_for_y_15_lpi_1_dfm_4_21_0_1 = MUX_v_22_2_2(22'b0000000000000000000000,
      Gelu_for_else_Gelu_for_else_mux1h_46_nl, Gelu_for_15_slc_32_1_svs);
  assign Gelu_for_else_Gelu_for_else_mux1h_30_nl = MUX1HOT_v_5_4_2((signext_5_1(Gelu_for_8_else_if_acc_itm_mx1w0[3])),
      (signext_5_1(Gelu_for_1_else_else_if_mul_cmp_2_z[46])), (signext_5_2(Gelu_for_y_15_sva_4_27_22_1[5:4])),
      act_write_data_data_0_14_sva_30_26, {(~ Gelu_for_15_else_slc_32_svs) , Gelu_for_else_and_28_ssc_1
      , Gelu_for_else_else_else_and_28_ssc_1 , Gelu_for_else_else_else_and_29_ssc_1});
  assign Gelu_for_y_15_lpi_1_dfm_4_30_26 = Gelu_for_else_Gelu_for_else_mux1h_30_nl
      & (signext_5_1(~ Gelu_for_else_and_46_ssc_1)) & ({{4{Gelu_for_15_slc_32_1_svs}},
      Gelu_for_15_slc_32_1_svs});
  assign Gelu_for_else_Gelu_for_else_mux1h_62_nl = MUX1HOT_s_1_4_2((Gelu_for_8_else_if_acc_itm_mx1w0[3]),
      (Gelu_for_1_else_else_if_mul_cmp_2_z[46]), (Gelu_for_y_15_sva_4_27_22_1[3]),
      act_write_data_data_0_14_sva_25, {(~ Gelu_for_15_else_slc_32_svs) , Gelu_for_else_and_28_ssc_1
      , Gelu_for_else_else_else_and_28_ssc_1 , Gelu_for_else_else_else_and_29_ssc_1});
  assign Gelu_for_y_15_lpi_1_dfm_4_25 = Gelu_for_else_Gelu_for_else_mux1h_62_nl &
      (~ Gelu_for_else_and_46_ssc_1) & Gelu_for_15_slc_32_1_svs;
  assign Gelu_for_else_Gelu_for_else_mux1h_78_nl = MUX1HOT_v_3_5_2((Gelu_for_8_else_if_acc_itm_mx1w0[2:0]),
      (signext_3_1(Gelu_for_1_else_else_if_mul_cmp_2_z[46])), (Gelu_for_1_else_else_else_if_mul_cmp_2_z[48:46]),
      (Gelu_for_y_15_sva_4_27_22_1[2:0]), act_write_data_data_0_14_sva_24_22, {(~
      Gelu_for_15_else_slc_32_svs) , Gelu_for_else_and_28_ssc_1 , Gelu_for_else_and_46_ssc_1
      , Gelu_for_else_else_else_and_28_ssc_1 , Gelu_for_else_else_else_and_29_ssc_1});
  assign Gelu_for_y_15_lpi_1_dfm_4_24_22 = MUX_v_3_2_2(3'b000, Gelu_for_else_Gelu_for_else_mux1h_78_nl,
      Gelu_for_15_slc_32_1_svs);
  assign Gelu_for_else_Gelu_for_else_mux1h_13_nl = MUX1HOT_s_1_3_2((Gelu_for_7_else_if_acc_itm_mx1w0[3]),
      (Gelu_for_1_else_else_if_mul_cmp_3_z[46]), (Gelu_for_y_14_sva_4_27_22_1[5]),
      {(~ Gelu_for_14_else_slc_32_svs) , Gelu_for_else_and_26_ssc_1 , Gelu_for_else_else_else_and_26_ssc_1});
  assign Gelu_for_y_14_lpi_1_dfm_4_31_1 = Gelu_for_else_Gelu_for_else_mux1h_13_nl
      & (~(Gelu_for_else_and_45_ssc_1 | Gelu_for_else_else_else_and_27_ssc_1)) &
      Gelu_for_14_slc_32_1_svs;
  assign Gelu_for_else_or_2_nl = Gelu_for_else_and_45_ssc_1 | Gelu_for_else_else_else_and_26_ssc_1;
  assign Gelu_for_else_Gelu_for_else_mux1h_45_nl = MUX1HOT_v_22_4_2((Silu_for_1_else_if_Silu_for_else_if_mul_cmp_2_z[44:23]),
      (Gelu_for_1_else_else_if_mul_cmp_3_z[45:24]), (Gelu_for_1_else_else_else_if_mul_cmp_3_z[45:24]),
      act_write_data_data_0_13_sva_21_0, {(~ Gelu_for_14_else_slc_32_svs) , Gelu_for_else_and_26_ssc_1
      , Gelu_for_else_or_2_nl , Gelu_for_else_else_else_and_27_ssc_1});
  assign Gelu_for_y_14_lpi_1_dfm_4_21_0_1 = MUX_v_22_2_2(22'b0000000000000000000000,
      Gelu_for_else_Gelu_for_else_mux1h_45_nl, Gelu_for_14_slc_32_1_svs);
  assign Gelu_for_else_Gelu_for_else_mux1h_29_nl = MUX1HOT_v_5_4_2((signext_5_1(Gelu_for_7_else_if_acc_itm_mx1w0[3])),
      (signext_5_1(Gelu_for_1_else_else_if_mul_cmp_3_z[46])), (signext_5_2(Gelu_for_y_14_sva_4_27_22_1[5:4])),
      act_write_data_data_0_13_sva_30_26, {(~ Gelu_for_14_else_slc_32_svs) , Gelu_for_else_and_26_ssc_1
      , Gelu_for_else_else_else_and_26_ssc_1 , Gelu_for_else_else_else_and_27_ssc_1});
  assign Gelu_for_y_14_lpi_1_dfm_4_30_26 = Gelu_for_else_Gelu_for_else_mux1h_29_nl
      & (signext_5_1(~ Gelu_for_else_and_45_ssc_1)) & ({{4{Gelu_for_14_slc_32_1_svs}},
      Gelu_for_14_slc_32_1_svs});
  assign Gelu_for_else_Gelu_for_else_mux1h_61_nl = MUX1HOT_s_1_4_2((Gelu_for_7_else_if_acc_itm_mx1w0[3]),
      (Gelu_for_1_else_else_if_mul_cmp_3_z[46]), (Gelu_for_y_14_sva_4_27_22_1[3]),
      act_write_data_data_0_13_sva_25, {(~ Gelu_for_14_else_slc_32_svs) , Gelu_for_else_and_26_ssc_1
      , Gelu_for_else_else_else_and_26_ssc_1 , Gelu_for_else_else_else_and_27_ssc_1});
  assign Gelu_for_y_14_lpi_1_dfm_4_25 = Gelu_for_else_Gelu_for_else_mux1h_61_nl &
      (~ Gelu_for_else_and_45_ssc_1) & Gelu_for_14_slc_32_1_svs;
  assign Gelu_for_else_Gelu_for_else_mux1h_77_nl = MUX1HOT_v_3_5_2((Gelu_for_7_else_if_acc_itm_mx1w0[2:0]),
      (signext_3_1(Gelu_for_1_else_else_if_mul_cmp_3_z[46])), (Gelu_for_1_else_else_else_if_mul_cmp_3_z[48:46]),
      (Gelu_for_y_14_sva_4_27_22_1[2:0]), act_write_data_data_0_13_sva_24_22, {(~
      Gelu_for_14_else_slc_32_svs) , Gelu_for_else_and_26_ssc_1 , Gelu_for_else_and_45_ssc_1
      , Gelu_for_else_else_else_and_26_ssc_1 , Gelu_for_else_else_else_and_27_ssc_1});
  assign Gelu_for_y_14_lpi_1_dfm_4_24_22 = MUX_v_3_2_2(3'b000, Gelu_for_else_Gelu_for_else_mux1h_77_nl,
      Gelu_for_14_slc_32_1_svs);
  assign Gelu_for_else_Gelu_for_else_mux1h_12_nl = MUX1HOT_s_1_3_2((Gelu_for_6_else_if_acc_itm_mx1w0[3]),
      (Gelu_for_1_else_else_if_mul_cmp_4_z[46]), (Gelu_for_y_13_sva_4_27_22_1[5]),
      {(~ Gelu_for_13_else_slc_32_svs) , Gelu_for_else_and_24_ssc_1 , Gelu_for_else_else_else_and_24_ssc_1});
  assign Gelu_for_y_13_lpi_1_dfm_4_31_1 = Gelu_for_else_Gelu_for_else_mux1h_12_nl
      & (~(Gelu_for_else_and_44_ssc_1 | Gelu_for_else_else_else_and_25_ssc_1)) &
      Gelu_for_13_slc_32_1_svs;
  assign Gelu_for_else_or_3_nl = Gelu_for_else_and_44_ssc_1 | Gelu_for_else_else_else_and_24_ssc_1;
  assign Gelu_for_else_Gelu_for_else_mux1h_44_nl = MUX1HOT_v_22_4_2((Silu_for_1_else_if_Silu_for_else_if_mul_cmp_3_z[44:23]),
      (Gelu_for_1_else_else_if_mul_cmp_4_z[45:24]), (Gelu_for_1_else_else_else_if_mul_cmp_4_z[45:24]),
      act_write_data_data_0_12_sva_21_0, {(~ Gelu_for_13_else_slc_32_svs) , Gelu_for_else_and_24_ssc_1
      , Gelu_for_else_or_3_nl , Gelu_for_else_else_else_and_25_ssc_1});
  assign Gelu_for_y_13_lpi_1_dfm_4_21_0_1 = MUX_v_22_2_2(22'b0000000000000000000000,
      Gelu_for_else_Gelu_for_else_mux1h_44_nl, Gelu_for_13_slc_32_1_svs);
  assign Gelu_for_else_Gelu_for_else_mux1h_28_nl = MUX1HOT_v_5_4_2((signext_5_1(Gelu_for_6_else_if_acc_itm_mx1w0[3])),
      (signext_5_1(Gelu_for_1_else_else_if_mul_cmp_4_z[46])), (signext_5_2(Gelu_for_y_13_sva_4_27_22_1[5:4])),
      act_write_data_data_0_12_sva_30_26, {(~ Gelu_for_13_else_slc_32_svs) , Gelu_for_else_and_24_ssc_1
      , Gelu_for_else_else_else_and_24_ssc_1 , Gelu_for_else_else_else_and_25_ssc_1});
  assign Gelu_for_y_13_lpi_1_dfm_4_30_26 = Gelu_for_else_Gelu_for_else_mux1h_28_nl
      & (signext_5_1(~ Gelu_for_else_and_44_ssc_1)) & ({{4{Gelu_for_13_slc_32_1_svs}},
      Gelu_for_13_slc_32_1_svs});
  assign Gelu_for_else_Gelu_for_else_mux1h_60_nl = MUX1HOT_s_1_4_2((Gelu_for_6_else_if_acc_itm_mx1w0[3]),
      (Gelu_for_1_else_else_if_mul_cmp_4_z[46]), (Gelu_for_y_13_sva_4_27_22_1[3]),
      act_write_data_data_0_12_sva_25, {(~ Gelu_for_13_else_slc_32_svs) , Gelu_for_else_and_24_ssc_1
      , Gelu_for_else_else_else_and_24_ssc_1 , Gelu_for_else_else_else_and_25_ssc_1});
  assign Gelu_for_y_13_lpi_1_dfm_4_25 = Gelu_for_else_Gelu_for_else_mux1h_60_nl &
      (~ Gelu_for_else_and_44_ssc_1) & Gelu_for_13_slc_32_1_svs;
  assign Gelu_for_else_Gelu_for_else_mux1h_76_nl = MUX1HOT_v_3_5_2((Gelu_for_6_else_if_acc_itm_mx1w0[2:0]),
      (signext_3_1(Gelu_for_1_else_else_if_mul_cmp_4_z[46])), (Gelu_for_1_else_else_else_if_mul_cmp_4_z[48:46]),
      (Gelu_for_y_13_sva_4_27_22_1[2:0]), act_write_data_data_0_12_sva_24_22, {(~
      Gelu_for_13_else_slc_32_svs) , Gelu_for_else_and_24_ssc_1 , Gelu_for_else_and_44_ssc_1
      , Gelu_for_else_else_else_and_24_ssc_1 , Gelu_for_else_else_else_and_25_ssc_1});
  assign Gelu_for_y_13_lpi_1_dfm_4_24_22 = MUX_v_3_2_2(3'b000, Gelu_for_else_Gelu_for_else_mux1h_76_nl,
      Gelu_for_13_slc_32_1_svs);
  assign Gelu_for_else_Gelu_for_else_mux1h_11_nl = MUX1HOT_s_1_3_2((Gelu_for_5_else_if_acc_itm_mx1w0[3]),
      (Gelu_for_1_else_else_if_mul_cmp_5_z[46]), (Gelu_for_y_12_sva_4_27_22_1[5]),
      {(~ Gelu_for_12_else_slc_32_svs) , Gelu_for_else_and_22_ssc_1 , Gelu_for_else_else_else_and_22_ssc_1});
  assign Gelu_for_y_12_lpi_1_dfm_4_31_1 = Gelu_for_else_Gelu_for_else_mux1h_11_nl
      & (~(Gelu_for_else_and_43_ssc_1 | Gelu_for_else_else_else_and_23_ssc_1)) &
      Gelu_for_12_slc_32_1_svs;
  assign Gelu_for_else_or_4_nl = Gelu_for_else_and_43_ssc_1 | Gelu_for_else_else_else_and_22_ssc_1;
  assign Gelu_for_else_Gelu_for_else_mux1h_43_nl = MUX1HOT_v_22_4_2((Silu_for_1_else_if_Silu_for_else_if_mul_cmp_4_z[44:23]),
      (Gelu_for_1_else_else_if_mul_cmp_5_z[45:24]), (Gelu_for_1_else_else_else_if_mul_cmp_5_z[45:24]),
      act_write_data_data_0_11_sva_21_0, {(~ Gelu_for_12_else_slc_32_svs) , Gelu_for_else_and_22_ssc_1
      , Gelu_for_else_or_4_nl , Gelu_for_else_else_else_and_23_ssc_1});
  assign Gelu_for_y_12_lpi_1_dfm_4_21_0_1 = MUX_v_22_2_2(22'b0000000000000000000000,
      Gelu_for_else_Gelu_for_else_mux1h_43_nl, Gelu_for_12_slc_32_1_svs);
  assign Gelu_for_else_Gelu_for_else_mux1h_27_nl = MUX1HOT_v_5_4_2((signext_5_1(Gelu_for_5_else_if_acc_itm_mx1w0[3])),
      (signext_5_1(Gelu_for_1_else_else_if_mul_cmp_5_z[46])), (signext_5_2(Gelu_for_y_12_sva_4_27_22_1[5:4])),
      act_write_data_data_0_11_sva_30_26, {(~ Gelu_for_12_else_slc_32_svs) , Gelu_for_else_and_22_ssc_1
      , Gelu_for_else_else_else_and_22_ssc_1 , Gelu_for_else_else_else_and_23_ssc_1});
  assign Gelu_for_y_12_lpi_1_dfm_4_30_26 = Gelu_for_else_Gelu_for_else_mux1h_27_nl
      & (signext_5_1(~ Gelu_for_else_and_43_ssc_1)) & ({{4{Gelu_for_12_slc_32_1_svs}},
      Gelu_for_12_slc_32_1_svs});
  assign Gelu_for_else_Gelu_for_else_mux1h_59_nl = MUX1HOT_s_1_4_2((Gelu_for_5_else_if_acc_itm_mx1w0[3]),
      (Gelu_for_1_else_else_if_mul_cmp_5_z[46]), (Gelu_for_y_12_sva_4_27_22_1[3]),
      act_write_data_data_0_11_sva_25, {(~ Gelu_for_12_else_slc_32_svs) , Gelu_for_else_and_22_ssc_1
      , Gelu_for_else_else_else_and_22_ssc_1 , Gelu_for_else_else_else_and_23_ssc_1});
  assign Gelu_for_y_12_lpi_1_dfm_4_25 = Gelu_for_else_Gelu_for_else_mux1h_59_nl &
      (~ Gelu_for_else_and_43_ssc_1) & Gelu_for_12_slc_32_1_svs;
  assign Gelu_for_else_Gelu_for_else_mux1h_75_nl = MUX1HOT_v_3_5_2((Gelu_for_5_else_if_acc_itm_mx1w0[2:0]),
      (signext_3_1(Gelu_for_1_else_else_if_mul_cmp_5_z[46])), (Gelu_for_1_else_else_else_if_mul_cmp_5_z[48:46]),
      (Gelu_for_y_12_sva_4_27_22_1[2:0]), act_write_data_data_0_11_sva_24_22, {(~
      Gelu_for_12_else_slc_32_svs) , Gelu_for_else_and_22_ssc_1 , Gelu_for_else_and_43_ssc_1
      , Gelu_for_else_else_else_and_22_ssc_1 , Gelu_for_else_else_else_and_23_ssc_1});
  assign Gelu_for_y_12_lpi_1_dfm_4_24_22 = MUX_v_3_2_2(3'b000, Gelu_for_else_Gelu_for_else_mux1h_75_nl,
      Gelu_for_12_slc_32_1_svs);
  assign Gelu_for_else_Gelu_for_else_mux1h_10_nl = MUX1HOT_s_1_3_2((Gelu_for_4_else_if_acc_itm_mx1w0[3]),
      (Gelu_for_1_else_else_if_mul_cmp_6_z[46]), (Gelu_for_y_11_sva_4_27_22_1[5]),
      {(~ Gelu_for_11_else_slc_32_svs) , Gelu_for_else_and_20_ssc_1 , Gelu_for_else_else_else_and_20_ssc_1});
  assign Gelu_for_y_11_lpi_1_dfm_4_31_1 = Gelu_for_else_Gelu_for_else_mux1h_10_nl
      & (~(Gelu_for_else_and_42_ssc_1 | Gelu_for_else_else_else_and_21_ssc_1)) &
      Gelu_for_11_slc_32_1_svs;
  assign Gelu_for_else_or_5_nl = Gelu_for_else_and_42_ssc_1 | Gelu_for_else_else_else_and_20_ssc_1;
  assign Gelu_for_else_Gelu_for_else_mux1h_42_nl = MUX1HOT_v_22_4_2((Silu_for_1_else_if_Silu_for_else_if_mul_cmp_5_z[44:23]),
      (Gelu_for_1_else_else_if_mul_cmp_6_z[45:24]), (Gelu_for_1_else_else_else_if_mul_cmp_6_z[45:24]),
      act_write_data_data_0_10_sva_21_0, {(~ Gelu_for_11_else_slc_32_svs) , Gelu_for_else_and_20_ssc_1
      , Gelu_for_else_or_5_nl , Gelu_for_else_else_else_and_21_ssc_1});
  assign Gelu_for_y_11_lpi_1_dfm_4_21_0_1 = MUX_v_22_2_2(22'b0000000000000000000000,
      Gelu_for_else_Gelu_for_else_mux1h_42_nl, Gelu_for_11_slc_32_1_svs);
  assign Gelu_for_else_Gelu_for_else_mux1h_26_nl = MUX1HOT_v_5_4_2((signext_5_1(Gelu_for_4_else_if_acc_itm_mx1w0[3])),
      (signext_5_1(Gelu_for_1_else_else_if_mul_cmp_6_z[46])), (signext_5_2(Gelu_for_y_11_sva_4_27_22_1[5:4])),
      act_write_data_data_0_10_sva_30_26, {(~ Gelu_for_11_else_slc_32_svs) , Gelu_for_else_and_20_ssc_1
      , Gelu_for_else_else_else_and_20_ssc_1 , Gelu_for_else_else_else_and_21_ssc_1});
  assign Gelu_for_y_11_lpi_1_dfm_4_30_26 = Gelu_for_else_Gelu_for_else_mux1h_26_nl
      & (signext_5_1(~ Gelu_for_else_and_42_ssc_1)) & ({{4{Gelu_for_11_slc_32_1_svs}},
      Gelu_for_11_slc_32_1_svs});
  assign Gelu_for_else_Gelu_for_else_mux1h_58_nl = MUX1HOT_s_1_4_2((Gelu_for_4_else_if_acc_itm_mx1w0[3]),
      (Gelu_for_1_else_else_if_mul_cmp_6_z[46]), (Gelu_for_y_11_sva_4_27_22_1[3]),
      act_write_data_data_0_10_sva_25, {(~ Gelu_for_11_else_slc_32_svs) , Gelu_for_else_and_20_ssc_1
      , Gelu_for_else_else_else_and_20_ssc_1 , Gelu_for_else_else_else_and_21_ssc_1});
  assign Gelu_for_y_11_lpi_1_dfm_4_25 = Gelu_for_else_Gelu_for_else_mux1h_58_nl &
      (~ Gelu_for_else_and_42_ssc_1) & Gelu_for_11_slc_32_1_svs;
  assign Gelu_for_else_Gelu_for_else_mux1h_74_nl = MUX1HOT_v_3_5_2((Gelu_for_4_else_if_acc_itm_mx1w0[2:0]),
      (signext_3_1(Gelu_for_1_else_else_if_mul_cmp_6_z[46])), (Gelu_for_1_else_else_else_if_mul_cmp_6_z[48:46]),
      (Gelu_for_y_11_sva_4_27_22_1[2:0]), act_write_data_data_0_10_sva_24_22, {(~
      Gelu_for_11_else_slc_32_svs) , Gelu_for_else_and_20_ssc_1 , Gelu_for_else_and_42_ssc_1
      , Gelu_for_else_else_else_and_20_ssc_1 , Gelu_for_else_else_else_and_21_ssc_1});
  assign Gelu_for_y_11_lpi_1_dfm_4_24_22 = MUX_v_3_2_2(3'b000, Gelu_for_else_Gelu_for_else_mux1h_74_nl,
      Gelu_for_11_slc_32_1_svs);
  assign Gelu_for_else_Gelu_for_else_mux1h_9_nl = MUX1HOT_s_1_3_2((Gelu_for_3_else_if_acc_itm_mx1w0[3]),
      (Gelu_for_1_else_else_if_mul_cmp_7_z[46]), (Gelu_for_y_10_sva_4_27_22_1[5]),
      {(~ Gelu_for_10_else_slc_32_svs) , Gelu_for_else_and_18_ssc_1 , Gelu_for_else_else_else_and_18_ssc_1});
  assign Gelu_for_y_10_lpi_1_dfm_4_31_1 = Gelu_for_else_Gelu_for_else_mux1h_9_nl
      & (~(Gelu_for_else_and_41_ssc_1 | Gelu_for_else_else_else_and_19_ssc_1)) &
      Gelu_for_10_slc_32_1_svs;
  assign Gelu_for_else_or_6_nl = Gelu_for_else_and_41_ssc_1 | Gelu_for_else_else_else_and_18_ssc_1;
  assign Gelu_for_else_Gelu_for_else_mux1h_41_nl = MUX1HOT_v_22_4_2((Silu_for_1_else_if_Silu_for_else_if_mul_cmp_6_z[44:23]),
      (Gelu_for_1_else_else_if_mul_cmp_7_z[45:24]), (Gelu_for_1_else_else_else_if_mul_cmp_7_z[45:24]),
      act_write_data_data_0_1_sva_21_0, {(~ Gelu_for_10_else_slc_32_svs) , Gelu_for_else_and_18_ssc_1
      , Gelu_for_else_or_6_nl , Gelu_for_else_else_else_and_19_ssc_1});
  assign Gelu_for_y_10_lpi_1_dfm_4_21_0_1 = MUX_v_22_2_2(22'b0000000000000000000000,
      Gelu_for_else_Gelu_for_else_mux1h_41_nl, Gelu_for_10_slc_32_1_svs);
  assign Gelu_for_else_Gelu_for_else_mux1h_25_nl = MUX1HOT_v_5_4_2((signext_5_1(Gelu_for_3_else_if_acc_itm_mx1w0[3])),
      (signext_5_1(Gelu_for_1_else_else_if_mul_cmp_7_z[46])), (signext_5_2(Gelu_for_y_10_sva_4_27_22_1[5:4])),
      act_write_data_data_0_1_sva_30_26, {(~ Gelu_for_10_else_slc_32_svs) , Gelu_for_else_and_18_ssc_1
      , Gelu_for_else_else_else_and_18_ssc_1 , Gelu_for_else_else_else_and_19_ssc_1});
  assign Gelu_for_y_10_lpi_1_dfm_4_30_26 = Gelu_for_else_Gelu_for_else_mux1h_25_nl
      & (signext_5_1(~ Gelu_for_else_and_41_ssc_1)) & ({{4{Gelu_for_10_slc_32_1_svs}},
      Gelu_for_10_slc_32_1_svs});
  assign Gelu_for_else_Gelu_for_else_mux1h_57_nl = MUX1HOT_s_1_4_2((Gelu_for_3_else_if_acc_itm_mx1w0[3]),
      (Gelu_for_1_else_else_if_mul_cmp_7_z[46]), (Gelu_for_y_10_sva_4_27_22_1[3]),
      act_write_data_data_0_1_sva_25, {(~ Gelu_for_10_else_slc_32_svs) , Gelu_for_else_and_18_ssc_1
      , Gelu_for_else_else_else_and_18_ssc_1 , Gelu_for_else_else_else_and_19_ssc_1});
  assign Gelu_for_y_10_lpi_1_dfm_4_25 = Gelu_for_else_Gelu_for_else_mux1h_57_nl &
      (~ Gelu_for_else_and_41_ssc_1) & Gelu_for_10_slc_32_1_svs;
  assign Gelu_for_else_Gelu_for_else_mux1h_73_nl = MUX1HOT_v_3_5_2((Gelu_for_3_else_if_acc_itm_mx1w0[2:0]),
      (signext_3_1(Gelu_for_1_else_else_if_mul_cmp_7_z[46])), (Gelu_for_1_else_else_else_if_mul_cmp_7_z[48:46]),
      (Gelu_for_y_10_sva_4_27_22_1[2:0]), act_write_data_data_0_1_sva_24_22, {(~
      Gelu_for_10_else_slc_32_svs) , Gelu_for_else_and_18_ssc_1 , Gelu_for_else_and_41_ssc_1
      , Gelu_for_else_else_else_and_18_ssc_1 , Gelu_for_else_else_else_and_19_ssc_1});
  assign Gelu_for_y_10_lpi_1_dfm_4_24_22 = MUX_v_3_2_2(3'b000, Gelu_for_else_Gelu_for_else_mux1h_73_nl,
      Gelu_for_10_slc_32_1_svs);
  assign Gelu_for_else_Gelu_for_else_mux1h_8_nl = MUX1HOT_s_1_3_2((Gelu_for_1_else_if_acc_itm_mx1w0[3]),
      (Gelu_for_1_else_else_if_mul_cmp_8_z[46]), (Gelu_for_y_9_sva_4_27_22_1[5]),
      {(~ Gelu_for_9_else_slc_32_svs) , Gelu_for_else_and_16_ssc_1 , Gelu_for_else_else_else_and_16_ssc_1});
  assign Gelu_for_y_9_lpi_1_dfm_4_31_1 = Gelu_for_else_Gelu_for_else_mux1h_8_nl &
      (~(Gelu_for_else_and_40_ssc_1 | Gelu_for_else_else_else_and_17_ssc_1)) & Gelu_for_9_slc_32_1_svs;
  assign Gelu_for_else_or_7_nl = Gelu_for_else_and_40_ssc_1 | Gelu_for_else_else_else_and_16_ssc_1;
  assign Gelu_for_else_Gelu_for_else_mux1h_40_nl = MUX1HOT_v_22_4_2((Silu_for_1_else_if_Silu_for_else_if_mul_cmp_7_z[44:23]),
      (Gelu_for_1_else_else_if_mul_cmp_8_z[45:24]), (Gelu_for_1_else_else_else_if_mul_cmp_8_z[45:24]),
      act_write_data_data_0_9_sva_21_0, {(~ Gelu_for_9_else_slc_32_svs) , Gelu_for_else_and_16_ssc_1
      , Gelu_for_else_or_7_nl , Gelu_for_else_else_else_and_17_ssc_1});
  assign Gelu_for_y_9_lpi_1_dfm_4_21_0_1 = MUX_v_22_2_2(22'b0000000000000000000000,
      Gelu_for_else_Gelu_for_else_mux1h_40_nl, Gelu_for_9_slc_32_1_svs);
  assign Gelu_for_else_Gelu_for_else_mux1h_24_nl = MUX1HOT_v_5_4_2((signext_5_1(Gelu_for_1_else_if_acc_itm_mx1w0[3])),
      (signext_5_1(Gelu_for_1_else_else_if_mul_cmp_8_z[46])), (signext_5_2(Gelu_for_y_9_sva_4_27_22_1[5:4])),
      act_write_data_data_0_9_sva_30_26, {(~ Gelu_for_9_else_slc_32_svs) , Gelu_for_else_and_16_ssc_1
      , Gelu_for_else_else_else_and_16_ssc_1 , Gelu_for_else_else_else_and_17_ssc_1});
  assign Gelu_for_y_9_lpi_1_dfm_4_30_26 = Gelu_for_else_Gelu_for_else_mux1h_24_nl
      & (signext_5_1(~ Gelu_for_else_and_40_ssc_1)) & ({{4{Gelu_for_9_slc_32_1_svs}},
      Gelu_for_9_slc_32_1_svs});
  assign Gelu_for_else_Gelu_for_else_mux1h_56_nl = MUX1HOT_s_1_4_2((Gelu_for_1_else_if_acc_itm_mx1w0[3]),
      (Gelu_for_1_else_else_if_mul_cmp_8_z[46]), (Gelu_for_y_9_sva_4_27_22_1[3]),
      act_write_data_data_0_9_sva_25, {(~ Gelu_for_9_else_slc_32_svs) , Gelu_for_else_and_16_ssc_1
      , Gelu_for_else_else_else_and_16_ssc_1 , Gelu_for_else_else_else_and_17_ssc_1});
  assign Gelu_for_y_9_lpi_1_dfm_4_25 = Gelu_for_else_Gelu_for_else_mux1h_56_nl &
      (~ Gelu_for_else_and_40_ssc_1) & Gelu_for_9_slc_32_1_svs;
  assign Gelu_for_else_Gelu_for_else_mux1h_72_nl = MUX1HOT_v_3_5_2((Gelu_for_1_else_if_acc_itm_mx1w0[2:0]),
      (signext_3_1(Gelu_for_1_else_else_if_mul_cmp_8_z[46])), (Gelu_for_1_else_else_else_if_mul_cmp_8_z[48:46]),
      (Gelu_for_y_9_sva_4_27_22_1[2:0]), act_write_data_data_0_9_sva_24_22, {(~ Gelu_for_9_else_slc_32_svs)
      , Gelu_for_else_and_16_ssc_1 , Gelu_for_else_and_40_ssc_1 , Gelu_for_else_else_else_and_16_ssc_1
      , Gelu_for_else_else_else_and_17_ssc_1});
  assign Gelu_for_y_9_lpi_1_dfm_4_24_22 = MUX_v_3_2_2(3'b000, Gelu_for_else_Gelu_for_else_mux1h_72_nl,
      Gelu_for_9_slc_32_1_svs);
  assign Gelu_for_else_Gelu_for_else_mux1h_7_nl = MUX1HOT_s_1_3_2((Gelu_for_8_else_if_acc_itm[3]),
      (Gelu_for_1_else_else_if_mul_cmp_9_z[46]), (Gelu_for_y_8_sva_4_27_22_1[5]),
      {(~ Gelu_for_8_else_slc_32_svs) , Gelu_for_else_and_14_ssc_1 , Gelu_for_else_else_else_and_14_ssc_1});
  assign Gelu_for_y_8_lpi_1_dfm_4_31_1 = Gelu_for_else_Gelu_for_else_mux1h_7_nl &
      (~(Gelu_for_else_and_39_ssc_1 | Gelu_for_else_else_else_and_15_ssc_1)) & Gelu_for_8_slc_32_1_svs;
  assign Gelu_for_else_or_8_nl = Gelu_for_else_and_39_ssc_1 | Gelu_for_else_else_else_and_14_ssc_1;
  assign Gelu_for_else_Gelu_for_else_mux1h_39_nl = MUX1HOT_v_22_4_2(Silu_for_2_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0,
      (Gelu_for_1_else_else_if_mul_cmp_9_z[45:24]), (Gelu_for_1_else_else_else_if_mul_cmp_9_z[45:24]),
      act_write_data_data_0_8_sva_21_0, {(~ Gelu_for_8_else_slc_32_svs) , Gelu_for_else_and_14_ssc_1
      , Gelu_for_else_or_8_nl , Gelu_for_else_else_else_and_15_ssc_1});
  assign Gelu_for_y_8_lpi_1_dfm_4_21_0_1 = MUX_v_22_2_2(22'b0000000000000000000000,
      Gelu_for_else_Gelu_for_else_mux1h_39_nl, Gelu_for_8_slc_32_1_svs);
  assign Gelu_for_else_Gelu_for_else_mux1h_23_nl = MUX1HOT_v_5_4_2((signext_5_1(Gelu_for_8_else_if_acc_itm[3])),
      (signext_5_1(Gelu_for_1_else_else_if_mul_cmp_9_z[46])), (signext_5_2(Gelu_for_y_8_sva_4_27_22_1[5:4])),
      act_write_data_data_0_8_sva_30_26, {(~ Gelu_for_8_else_slc_32_svs) , Gelu_for_else_and_14_ssc_1
      , Gelu_for_else_else_else_and_14_ssc_1 , Gelu_for_else_else_else_and_15_ssc_1});
  assign Gelu_for_y_8_lpi_1_dfm_4_30_26 = Gelu_for_else_Gelu_for_else_mux1h_23_nl
      & (signext_5_1(~ Gelu_for_else_and_39_ssc_1)) & ({{4{Gelu_for_8_slc_32_1_svs}},
      Gelu_for_8_slc_32_1_svs});
  assign Gelu_for_else_Gelu_for_else_mux1h_55_nl = MUX1HOT_s_1_4_2((Gelu_for_8_else_if_acc_itm[3]),
      (Gelu_for_1_else_else_if_mul_cmp_9_z[46]), (Gelu_for_y_8_sva_4_27_22_1[3]),
      act_write_data_data_0_8_sva_25, {(~ Gelu_for_8_else_slc_32_svs) , Gelu_for_else_and_14_ssc_1
      , Gelu_for_else_else_else_and_14_ssc_1 , Gelu_for_else_else_else_and_15_ssc_1});
  assign Gelu_for_y_8_lpi_1_dfm_4_25 = Gelu_for_else_Gelu_for_else_mux1h_55_nl &
      (~ Gelu_for_else_and_39_ssc_1) & Gelu_for_8_slc_32_1_svs;
  assign Gelu_for_else_Gelu_for_else_mux1h_71_nl = MUX1HOT_v_3_5_2((Gelu_for_8_else_if_acc_itm[2:0]),
      (signext_3_1(Gelu_for_1_else_else_if_mul_cmp_9_z[46])), (Gelu_for_1_else_else_else_if_mul_cmp_9_z[48:46]),
      (Gelu_for_y_8_sva_4_27_22_1[2:0]), act_write_data_data_0_8_sva_24_22, {(~ Gelu_for_8_else_slc_32_svs)
      , Gelu_for_else_and_14_ssc_1 , Gelu_for_else_and_39_ssc_1 , Gelu_for_else_else_else_and_14_ssc_1
      , Gelu_for_else_else_else_and_15_ssc_1});
  assign Gelu_for_y_8_lpi_1_dfm_4_24_22 = MUX_v_3_2_2(3'b000, Gelu_for_else_Gelu_for_else_mux1h_71_nl,
      Gelu_for_8_slc_32_1_svs);
  assign Gelu_for_else_Gelu_for_else_mux1h_6_nl = MUX1HOT_s_1_3_2((Gelu_for_7_else_if_acc_itm[3]),
      (Gelu_for_1_else_else_if_mul_cmp_10_z[46]), (Gelu_for_y_7_sva_4_27_22_1[5]),
      {(~ Gelu_for_7_else_slc_32_svs) , Gelu_for_else_and_12_ssc_1 , Gelu_for_else_else_else_and_12_ssc_1});
  assign Gelu_for_y_7_lpi_1_dfm_4_31_1 = Gelu_for_else_Gelu_for_else_mux1h_6_nl &
      (~(Gelu_for_else_and_38_ssc_1 | Gelu_for_else_else_else_and_13_ssc_1)) & Gelu_for_7_slc_32_1_svs;
  assign Gelu_for_else_or_9_nl = Gelu_for_else_and_38_ssc_1 | Gelu_for_else_else_else_and_12_ssc_1;
  assign Gelu_for_else_Gelu_for_else_mux1h_38_nl = MUX1HOT_v_22_4_2(reg_Silu_for_16_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1,
      (Gelu_for_1_else_else_if_mul_cmp_10_z[45:24]), (Gelu_for_1_else_else_else_if_mul_cmp_10_z[45:24]),
      act_write_data_data_0_7_sva_21_0, {(~ Gelu_for_7_else_slc_32_svs) , Gelu_for_else_and_12_ssc_1
      , Gelu_for_else_or_9_nl , Gelu_for_else_else_else_and_13_ssc_1});
  assign Gelu_for_y_7_lpi_1_dfm_4_21_0_1 = MUX_v_22_2_2(22'b0000000000000000000000,
      Gelu_for_else_Gelu_for_else_mux1h_38_nl, Gelu_for_7_slc_32_1_svs);
  assign Gelu_for_else_Gelu_for_else_mux1h_22_nl = MUX1HOT_v_5_4_2((signext_5_1(Gelu_for_7_else_if_acc_itm[3])),
      (signext_5_1(Gelu_for_1_else_else_if_mul_cmp_10_z[46])), (signext_5_2(Gelu_for_y_7_sva_4_27_22_1[5:4])),
      act_write_data_data_0_7_sva_30_26, {(~ Gelu_for_7_else_slc_32_svs) , Gelu_for_else_and_12_ssc_1
      , Gelu_for_else_else_else_and_12_ssc_1 , Gelu_for_else_else_else_and_13_ssc_1});
  assign Gelu_for_y_7_lpi_1_dfm_4_30_26 = Gelu_for_else_Gelu_for_else_mux1h_22_nl
      & (signext_5_1(~ Gelu_for_else_and_38_ssc_1)) & ({{4{Gelu_for_7_slc_32_1_svs}},
      Gelu_for_7_slc_32_1_svs});
  assign Gelu_for_else_Gelu_for_else_mux1h_54_nl = MUX1HOT_s_1_4_2((Gelu_for_7_else_if_acc_itm[3]),
      (Gelu_for_1_else_else_if_mul_cmp_10_z[46]), (Gelu_for_y_7_sva_4_27_22_1[3]),
      act_write_data_data_0_7_sva_25, {(~ Gelu_for_7_else_slc_32_svs) , Gelu_for_else_and_12_ssc_1
      , Gelu_for_else_else_else_and_12_ssc_1 , Gelu_for_else_else_else_and_13_ssc_1});
  assign Gelu_for_y_7_lpi_1_dfm_4_25 = Gelu_for_else_Gelu_for_else_mux1h_54_nl &
      (~ Gelu_for_else_and_38_ssc_1) & Gelu_for_7_slc_32_1_svs;
  assign Gelu_for_else_Gelu_for_else_mux1h_70_nl = MUX1HOT_v_3_5_2((Gelu_for_7_else_if_acc_itm[2:0]),
      (signext_3_1(Gelu_for_1_else_else_if_mul_cmp_10_z[46])), (Gelu_for_1_else_else_else_if_mul_cmp_10_z[48:46]),
      (Gelu_for_y_7_sva_4_27_22_1[2:0]), act_write_data_data_0_7_sva_24_22, {(~ Gelu_for_7_else_slc_32_svs)
      , Gelu_for_else_and_12_ssc_1 , Gelu_for_else_and_38_ssc_1 , Gelu_for_else_else_else_and_12_ssc_1
      , Gelu_for_else_else_else_and_13_ssc_1});
  assign Gelu_for_y_7_lpi_1_dfm_4_24_22 = MUX_v_3_2_2(3'b000, Gelu_for_else_Gelu_for_else_mux1h_70_nl,
      Gelu_for_7_slc_32_1_svs);
  assign Gelu_for_else_Gelu_for_else_mux1h_5_nl = MUX1HOT_s_1_3_2((Gelu_for_6_else_if_acc_itm[3]),
      (Gelu_for_1_else_else_if_mul_cmp_11_z[46]), (Gelu_for_y_6_sva_4_27_22_1[5]),
      {(~ Gelu_for_6_else_slc_32_svs) , Gelu_for_else_and_10_ssc_1 , Gelu_for_else_else_else_and_10_ssc_1});
  assign Gelu_for_y_6_lpi_1_dfm_4_31_1 = Gelu_for_else_Gelu_for_else_mux1h_5_nl &
      (~(Gelu_for_else_and_37_ssc_1 | Gelu_for_else_else_else_and_11_ssc_1)) & Gelu_for_6_slc_32_1_svs;
  assign Gelu_for_else_or_10_nl = Gelu_for_else_and_37_ssc_1 | Gelu_for_else_else_else_and_10_ssc_1;
  assign Gelu_for_else_Gelu_for_else_mux1h_37_nl = MUX1HOT_v_22_4_2(reg_Silu_for_15_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1,
      (Gelu_for_1_else_else_if_mul_cmp_11_z[45:24]), (Gelu_for_1_else_else_else_if_mul_cmp_11_z[45:24]),
      act_write_data_data_0_6_sva_21_0, {(~ Gelu_for_6_else_slc_32_svs) , Gelu_for_else_and_10_ssc_1
      , Gelu_for_else_or_10_nl , Gelu_for_else_else_else_and_11_ssc_1});
  assign Gelu_for_y_6_lpi_1_dfm_4_21_0_1 = MUX_v_22_2_2(22'b0000000000000000000000,
      Gelu_for_else_Gelu_for_else_mux1h_37_nl, Gelu_for_6_slc_32_1_svs);
  assign Gelu_for_else_Gelu_for_else_mux1h_21_nl = MUX1HOT_v_5_4_2((signext_5_1(Gelu_for_6_else_if_acc_itm[3])),
      (signext_5_1(Gelu_for_1_else_else_if_mul_cmp_11_z[46])), (signext_5_2(Gelu_for_y_6_sva_4_27_22_1[5:4])),
      act_write_data_data_0_6_sva_30_26, {(~ Gelu_for_6_else_slc_32_svs) , Gelu_for_else_and_10_ssc_1
      , Gelu_for_else_else_else_and_10_ssc_1 , Gelu_for_else_else_else_and_11_ssc_1});
  assign Gelu_for_y_6_lpi_1_dfm_4_30_26 = Gelu_for_else_Gelu_for_else_mux1h_21_nl
      & (signext_5_1(~ Gelu_for_else_and_37_ssc_1)) & ({{4{Gelu_for_6_slc_32_1_svs}},
      Gelu_for_6_slc_32_1_svs});
  assign Gelu_for_else_Gelu_for_else_mux1h_53_nl = MUX1HOT_s_1_4_2((Gelu_for_6_else_if_acc_itm[3]),
      (Gelu_for_1_else_else_if_mul_cmp_11_z[46]), (Gelu_for_y_6_sva_4_27_22_1[3]),
      act_write_data_data_0_6_sva_25, {(~ Gelu_for_6_else_slc_32_svs) , Gelu_for_else_and_10_ssc_1
      , Gelu_for_else_else_else_and_10_ssc_1 , Gelu_for_else_else_else_and_11_ssc_1});
  assign Gelu_for_y_6_lpi_1_dfm_4_25 = Gelu_for_else_Gelu_for_else_mux1h_53_nl &
      (~ Gelu_for_else_and_37_ssc_1) & Gelu_for_6_slc_32_1_svs;
  assign Gelu_for_else_Gelu_for_else_mux1h_69_nl = MUX1HOT_v_3_5_2((Gelu_for_6_else_if_acc_itm[2:0]),
      (signext_3_1(Gelu_for_1_else_else_if_mul_cmp_11_z[46])), (Gelu_for_1_else_else_else_if_mul_cmp_11_z[48:46]),
      (Gelu_for_y_6_sva_4_27_22_1[2:0]), act_write_data_data_0_6_sva_24_22, {(~ Gelu_for_6_else_slc_32_svs)
      , Gelu_for_else_and_10_ssc_1 , Gelu_for_else_and_37_ssc_1 , Gelu_for_else_else_else_and_10_ssc_1
      , Gelu_for_else_else_else_and_11_ssc_1});
  assign Gelu_for_y_6_lpi_1_dfm_4_24_22 = MUX_v_3_2_2(3'b000, Gelu_for_else_Gelu_for_else_mux1h_69_nl,
      Gelu_for_6_slc_32_1_svs);
  assign Gelu_for_else_Gelu_for_else_mux1h_4_nl = MUX1HOT_s_1_3_2((Gelu_for_5_else_if_acc_itm[3]),
      (Gelu_for_1_else_else_if_mul_cmp_12_z[46]), (Gelu_for_y_5_sva_4_27_22_1[5]),
      {(~ Gelu_for_5_else_slc_32_svs) , Gelu_for_else_and_8_ssc_1 , Gelu_for_else_else_else_and_8_ssc_1});
  assign Gelu_for_y_5_lpi_1_dfm_4_31_1 = Gelu_for_else_Gelu_for_else_mux1h_4_nl &
      (~(Gelu_for_else_and_36_ssc_1 | Gelu_for_else_else_else_and_9_ssc_1)) & Gelu_for_5_slc_32_1_svs;
  assign Gelu_for_else_or_11_nl = Gelu_for_else_and_36_ssc_1 | Gelu_for_else_else_else_and_8_ssc_1;
  assign Gelu_for_else_Gelu_for_else_mux1h_36_nl = MUX1HOT_v_22_4_2(reg_Silu_for_14_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1,
      (Gelu_for_1_else_else_if_mul_cmp_12_z[45:24]), (Gelu_for_1_else_else_else_if_mul_cmp_12_z[45:24]),
      act_write_data_data_0_5_sva_21_0, {(~ Gelu_for_5_else_slc_32_svs) , Gelu_for_else_and_8_ssc_1
      , Gelu_for_else_or_11_nl , Gelu_for_else_else_else_and_9_ssc_1});
  assign Gelu_for_y_5_lpi_1_dfm_4_21_0_1 = MUX_v_22_2_2(22'b0000000000000000000000,
      Gelu_for_else_Gelu_for_else_mux1h_36_nl, Gelu_for_5_slc_32_1_svs);
  assign Gelu_for_else_Gelu_for_else_mux1h_20_nl = MUX1HOT_v_5_4_2((signext_5_1(Gelu_for_5_else_if_acc_itm[3])),
      (signext_5_1(Gelu_for_1_else_else_if_mul_cmp_12_z[46])), (signext_5_2(Gelu_for_y_5_sva_4_27_22_1[5:4])),
      act_write_data_data_0_5_sva_30_26, {(~ Gelu_for_5_else_slc_32_svs) , Gelu_for_else_and_8_ssc_1
      , Gelu_for_else_else_else_and_8_ssc_1 , Gelu_for_else_else_else_and_9_ssc_1});
  assign Gelu_for_y_5_lpi_1_dfm_4_30_26 = Gelu_for_else_Gelu_for_else_mux1h_20_nl
      & (signext_5_1(~ Gelu_for_else_and_36_ssc_1)) & ({{4{Gelu_for_5_slc_32_1_svs}},
      Gelu_for_5_slc_32_1_svs});
  assign Gelu_for_else_Gelu_for_else_mux1h_52_nl = MUX1HOT_s_1_4_2((Gelu_for_5_else_if_acc_itm[3]),
      (Gelu_for_1_else_else_if_mul_cmp_12_z[46]), (Gelu_for_y_5_sva_4_27_22_1[3]),
      act_write_data_data_0_5_sva_25, {(~ Gelu_for_5_else_slc_32_svs) , Gelu_for_else_and_8_ssc_1
      , Gelu_for_else_else_else_and_8_ssc_1 , Gelu_for_else_else_else_and_9_ssc_1});
  assign Gelu_for_y_5_lpi_1_dfm_4_25 = Gelu_for_else_Gelu_for_else_mux1h_52_nl &
      (~ Gelu_for_else_and_36_ssc_1) & Gelu_for_5_slc_32_1_svs;
  assign Gelu_for_else_Gelu_for_else_mux1h_68_nl = MUX1HOT_v_3_5_2((Gelu_for_5_else_if_acc_itm[2:0]),
      (signext_3_1(Gelu_for_1_else_else_if_mul_cmp_12_z[46])), (Gelu_for_1_else_else_else_if_mul_cmp_12_z[48:46]),
      (Gelu_for_y_5_sva_4_27_22_1[2:0]), act_write_data_data_0_5_sva_24_22, {(~ Gelu_for_5_else_slc_32_svs)
      , Gelu_for_else_and_8_ssc_1 , Gelu_for_else_and_36_ssc_1 , Gelu_for_else_else_else_and_8_ssc_1
      , Gelu_for_else_else_else_and_9_ssc_1});
  assign Gelu_for_y_5_lpi_1_dfm_4_24_22 = MUX_v_3_2_2(3'b000, Gelu_for_else_Gelu_for_else_mux1h_68_nl,
      Gelu_for_5_slc_32_1_svs);
  assign Gelu_for_else_Gelu_for_else_mux1h_3_nl = MUX1HOT_s_1_3_2((Gelu_for_4_else_if_acc_itm[3]),
      (Gelu_for_1_else_else_if_mul_cmp_13_z[46]), (Gelu_for_y_4_sva_4_27_22_1[5]),
      {(~ Gelu_for_4_else_slc_32_svs) , Gelu_for_else_and_6_ssc_1 , Gelu_for_else_else_else_and_6_ssc_1});
  assign Gelu_for_y_4_lpi_1_dfm_4_31_1 = Gelu_for_else_Gelu_for_else_mux1h_3_nl &
      (~(Gelu_for_else_and_35_ssc_1 | Gelu_for_else_else_else_and_7_ssc_1)) & Gelu_for_4_slc_32_1_svs;
  assign Gelu_for_else_or_12_nl = Gelu_for_else_and_35_ssc_1 | Gelu_for_else_else_else_and_6_ssc_1;
  assign Gelu_for_else_Gelu_for_else_mux1h_35_nl = MUX1HOT_v_22_4_2(reg_Silu_for_13_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1,
      (Gelu_for_1_else_else_if_mul_cmp_13_z[45:24]), (Gelu_for_1_else_else_else_if_mul_cmp_13_z[45:24]),
      act_write_data_data_0_4_sva_21_0, {(~ Gelu_for_4_else_slc_32_svs) , Gelu_for_else_and_6_ssc_1
      , Gelu_for_else_or_12_nl , Gelu_for_else_else_else_and_7_ssc_1});
  assign Gelu_for_y_4_lpi_1_dfm_4_21_0_1 = MUX_v_22_2_2(22'b0000000000000000000000,
      Gelu_for_else_Gelu_for_else_mux1h_35_nl, Gelu_for_4_slc_32_1_svs);
  assign Gelu_for_else_Gelu_for_else_mux1h_19_nl = MUX1HOT_v_5_4_2((signext_5_1(Gelu_for_4_else_if_acc_itm[3])),
      (signext_5_1(Gelu_for_1_else_else_if_mul_cmp_13_z[46])), (signext_5_2(Gelu_for_y_4_sva_4_27_22_1[5:4])),
      act_write_data_data_0_4_sva_30_26, {(~ Gelu_for_4_else_slc_32_svs) , Gelu_for_else_and_6_ssc_1
      , Gelu_for_else_else_else_and_6_ssc_1 , Gelu_for_else_else_else_and_7_ssc_1});
  assign Gelu_for_y_4_lpi_1_dfm_4_30_26 = Gelu_for_else_Gelu_for_else_mux1h_19_nl
      & (signext_5_1(~ Gelu_for_else_and_35_ssc_1)) & ({{4{Gelu_for_4_slc_32_1_svs}},
      Gelu_for_4_slc_32_1_svs});
  assign Gelu_for_else_Gelu_for_else_mux1h_51_nl = MUX1HOT_s_1_4_2((Gelu_for_4_else_if_acc_itm[3]),
      (Gelu_for_1_else_else_if_mul_cmp_13_z[46]), (Gelu_for_y_4_sva_4_27_22_1[3]),
      act_write_data_data_0_4_sva_25, {(~ Gelu_for_4_else_slc_32_svs) , Gelu_for_else_and_6_ssc_1
      , Gelu_for_else_else_else_and_6_ssc_1 , Gelu_for_else_else_else_and_7_ssc_1});
  assign Gelu_for_y_4_lpi_1_dfm_4_25 = Gelu_for_else_Gelu_for_else_mux1h_51_nl &
      (~ Gelu_for_else_and_35_ssc_1) & Gelu_for_4_slc_32_1_svs;
  assign Gelu_for_else_Gelu_for_else_mux1h_67_nl = MUX1HOT_v_3_5_2((Gelu_for_4_else_if_acc_itm[2:0]),
      (signext_3_1(Gelu_for_1_else_else_if_mul_cmp_13_z[46])), (Gelu_for_1_else_else_else_if_mul_cmp_13_z[48:46]),
      (Gelu_for_y_4_sva_4_27_22_1[2:0]), act_write_data_data_0_4_sva_24_22, {(~ Gelu_for_4_else_slc_32_svs)
      , Gelu_for_else_and_6_ssc_1 , Gelu_for_else_and_35_ssc_1 , Gelu_for_else_else_else_and_6_ssc_1
      , Gelu_for_else_else_else_and_7_ssc_1});
  assign Gelu_for_y_4_lpi_1_dfm_4_24_22 = MUX_v_3_2_2(3'b000, Gelu_for_else_Gelu_for_else_mux1h_67_nl,
      Gelu_for_4_slc_32_1_svs);
  assign Gelu_for_else_Gelu_for_else_mux1h_2_nl = MUX1HOT_s_1_3_2((Gelu_for_3_else_if_acc_itm[3]),
      (Gelu_for_1_else_else_if_mul_cmp_14_z[46]), (Gelu_for_y_3_sva_4_27_22_1[5]),
      {(~ Gelu_for_3_else_slc_32_svs) , Gelu_for_else_and_4_ssc_1 , Gelu_for_else_else_else_and_4_ssc_1});
  assign Gelu_for_y_3_lpi_1_dfm_4_31_1 = Gelu_for_else_Gelu_for_else_mux1h_2_nl &
      (~(Gelu_for_else_and_34_ssc_1 | Gelu_for_else_else_else_and_5_ssc_1)) & Gelu_for_3_slc_32_1_svs;
  assign Gelu_for_else_or_13_nl = Gelu_for_else_and_34_ssc_1 | Gelu_for_else_else_else_and_4_ssc_1;
  assign Gelu_for_else_Gelu_for_else_mux1h_34_nl = MUX1HOT_v_22_4_2(reg_Silu_for_12_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1,
      (Gelu_for_1_else_else_if_mul_cmp_14_z[45:24]), (Gelu_for_1_else_else_else_if_mul_cmp_14_z[45:24]),
      act_write_data_data_0_3_sva_21_0, {(~ Gelu_for_3_else_slc_32_svs) , Gelu_for_else_and_4_ssc_1
      , Gelu_for_else_or_13_nl , Gelu_for_else_else_else_and_5_ssc_1});
  assign Gelu_for_y_3_lpi_1_dfm_4_21_0_1 = MUX_v_22_2_2(22'b0000000000000000000000,
      Gelu_for_else_Gelu_for_else_mux1h_34_nl, Gelu_for_3_slc_32_1_svs);
  assign Gelu_for_else_Gelu_for_else_mux1h_18_nl = MUX1HOT_v_5_4_2((signext_5_1(Gelu_for_3_else_if_acc_itm[3])),
      (signext_5_1(Gelu_for_1_else_else_if_mul_cmp_14_z[46])), (signext_5_2(Gelu_for_y_3_sva_4_27_22_1[5:4])),
      act_write_data_data_0_3_sva_30_26, {(~ Gelu_for_3_else_slc_32_svs) , Gelu_for_else_and_4_ssc_1
      , Gelu_for_else_else_else_and_4_ssc_1 , Gelu_for_else_else_else_and_5_ssc_1});
  assign Gelu_for_y_3_lpi_1_dfm_4_30_26 = Gelu_for_else_Gelu_for_else_mux1h_18_nl
      & (signext_5_1(~ Gelu_for_else_and_34_ssc_1)) & ({{4{Gelu_for_3_slc_32_1_svs}},
      Gelu_for_3_slc_32_1_svs});
  assign Gelu_for_else_Gelu_for_else_mux1h_50_nl = MUX1HOT_s_1_4_2((Gelu_for_3_else_if_acc_itm[3]),
      (Gelu_for_1_else_else_if_mul_cmp_14_z[46]), (Gelu_for_y_3_sva_4_27_22_1[3]),
      act_write_data_data_0_3_sva_25, {(~ Gelu_for_3_else_slc_32_svs) , Gelu_for_else_and_4_ssc_1
      , Gelu_for_else_else_else_and_4_ssc_1 , Gelu_for_else_else_else_and_5_ssc_1});
  assign Gelu_for_y_3_lpi_1_dfm_4_25 = Gelu_for_else_Gelu_for_else_mux1h_50_nl &
      (~ Gelu_for_else_and_34_ssc_1) & Gelu_for_3_slc_32_1_svs;
  assign Gelu_for_else_Gelu_for_else_mux1h_66_nl = MUX1HOT_v_3_5_2((Gelu_for_3_else_if_acc_itm[2:0]),
      (signext_3_1(Gelu_for_1_else_else_if_mul_cmp_14_z[46])), (Gelu_for_1_else_else_else_if_mul_cmp_14_z[48:46]),
      (Gelu_for_y_3_sva_4_27_22_1[2:0]), act_write_data_data_0_3_sva_24_22, {(~ Gelu_for_3_else_slc_32_svs)
      , Gelu_for_else_and_4_ssc_1 , Gelu_for_else_and_34_ssc_1 , Gelu_for_else_else_else_and_4_ssc_1
      , Gelu_for_else_else_else_and_5_ssc_1});
  assign Gelu_for_y_3_lpi_1_dfm_4_24_22 = MUX_v_3_2_2(3'b000, Gelu_for_else_Gelu_for_else_mux1h_66_nl,
      Gelu_for_3_slc_32_1_svs);
  assign Gelu_for_else_Gelu_for_else_mux1h_1_nl = MUX1HOT_s_1_3_2((Gelu_for_2_else_if_acc_itm[3]),
      (Gelu_for_1_else_else_if_mul_cmp_15_z[46]), (Gelu_for_y_2_sva_4_27_22_1[5]),
      {(~ Gelu_for_2_else_slc_32_svs) , Gelu_for_else_and_2_ssc_1 , Gelu_for_else_else_else_and_2_ssc_1});
  assign Gelu_for_y_2_lpi_1_dfm_4_31_1 = Gelu_for_else_Gelu_for_else_mux1h_1_nl &
      (~(Gelu_for_else_and_33_ssc_1 | Gelu_for_else_else_else_and_3_ssc_1)) & Gelu_for_2_slc_32_1_svs;
  assign Gelu_for_else_or_14_nl = Gelu_for_else_and_33_ssc_1 | Gelu_for_else_else_else_and_2_ssc_1;
  assign Gelu_for_else_Gelu_for_else_mux1h_33_nl = MUX1HOT_v_22_4_2(reg_Silu_for_11_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1,
      (Gelu_for_1_else_else_if_mul_cmp_15_z[45:24]), (Gelu_for_1_else_else_else_if_mul_cmp_15_z[45:24]),
      act_write_data_data_0_2_sva_21_0, {(~ Gelu_for_2_else_slc_32_svs) , Gelu_for_else_and_2_ssc_1
      , Gelu_for_else_or_14_nl , Gelu_for_else_else_else_and_3_ssc_1});
  assign Gelu_for_y_2_lpi_1_dfm_4_21_0_1 = MUX_v_22_2_2(22'b0000000000000000000000,
      Gelu_for_else_Gelu_for_else_mux1h_33_nl, Gelu_for_2_slc_32_1_svs);
  assign Gelu_for_else_Gelu_for_else_mux1h_17_nl = MUX1HOT_v_5_4_2((signext_5_1(Gelu_for_2_else_if_acc_itm[3])),
      (signext_5_1(Gelu_for_1_else_else_if_mul_cmp_15_z[46])), (signext_5_2(Gelu_for_y_2_sva_4_27_22_1[5:4])),
      act_write_data_data_0_2_sva_30_26, {(~ Gelu_for_2_else_slc_32_svs) , Gelu_for_else_and_2_ssc_1
      , Gelu_for_else_else_else_and_2_ssc_1 , Gelu_for_else_else_else_and_3_ssc_1});
  assign Gelu_for_y_2_lpi_1_dfm_4_30_26 = Gelu_for_else_Gelu_for_else_mux1h_17_nl
      & (signext_5_1(~ Gelu_for_else_and_33_ssc_1)) & ({{4{Gelu_for_2_slc_32_1_svs}},
      Gelu_for_2_slc_32_1_svs});
  assign Gelu_for_else_Gelu_for_else_mux1h_49_nl = MUX1HOT_s_1_4_2((Gelu_for_2_else_if_acc_itm[3]),
      (Gelu_for_1_else_else_if_mul_cmp_15_z[46]), (Gelu_for_y_2_sva_4_27_22_1[3]),
      act_write_data_data_0_2_sva_25, {(~ Gelu_for_2_else_slc_32_svs) , Gelu_for_else_and_2_ssc_1
      , Gelu_for_else_else_else_and_2_ssc_1 , Gelu_for_else_else_else_and_3_ssc_1});
  assign Gelu_for_y_2_lpi_1_dfm_4_25 = Gelu_for_else_Gelu_for_else_mux1h_49_nl &
      (~ Gelu_for_else_and_33_ssc_1) & Gelu_for_2_slc_32_1_svs;
  assign Gelu_for_else_Gelu_for_else_mux1h_65_nl = MUX1HOT_v_3_5_2((Gelu_for_2_else_if_acc_itm[2:0]),
      (signext_3_1(Gelu_for_1_else_else_if_mul_cmp_15_z[46])), (Gelu_for_1_else_else_else_if_mul_cmp_15_z[48:46]),
      (Gelu_for_y_2_sva_4_27_22_1[2:0]), act_write_data_data_0_2_sva_24_22, {(~ Gelu_for_2_else_slc_32_svs)
      , Gelu_for_else_and_2_ssc_1 , Gelu_for_else_and_33_ssc_1 , Gelu_for_else_else_else_and_2_ssc_1
      , Gelu_for_else_else_else_and_3_ssc_1});
  assign Gelu_for_y_2_lpi_1_dfm_4_24_22 = MUX_v_3_2_2(3'b000, Gelu_for_else_Gelu_for_else_mux1h_65_nl,
      Gelu_for_2_slc_32_1_svs);
  assign Gelu_for_else_Gelu_for_else_mux1h_nl = MUX1HOT_s_1_3_2((Gelu_for_1_else_if_acc_itm[3]),
      (Gelu_for_1_else_else_if_mul_cmp_z[46]), (Gelu_for_y_1_sva_4_27_22_1[5]), {(~
      Gelu_for_1_else_slc_32_svs) , Gelu_for_else_and_ssc_1 , Gelu_for_else_else_else_and_ssc_1});
  assign Gelu_for_y_1_lpi_1_dfm_4_31_1 = Gelu_for_else_Gelu_for_else_mux1h_nl & (~(Gelu_for_else_and_32_ssc_1
      | Gelu_for_else_else_else_and_1_ssc_1)) & Gelu_for_1_slc_32_1_svs;
  assign Gelu_for_else_or_15_nl = Gelu_for_else_and_32_ssc_1 | Gelu_for_else_else_else_and_ssc_1;
  assign Gelu_for_else_Gelu_for_else_mux1h_32_nl = MUX1HOT_v_22_4_2(reg_Silu_for_10_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1,
      (Gelu_for_1_else_else_if_mul_cmp_z[45:24]), (Gelu_for_1_else_else_else_if_mul_cmp_z[45:24]),
      act_write_data_data_0_0_sva_21_0, {(~ Gelu_for_1_else_slc_32_svs) , Gelu_for_else_and_ssc_1
      , Gelu_for_else_or_15_nl , Gelu_for_else_else_else_and_1_ssc_1});
  assign Gelu_for_y_1_lpi_1_dfm_4_21_0_1 = MUX_v_22_2_2(22'b0000000000000000000000,
      Gelu_for_else_Gelu_for_else_mux1h_32_nl, Gelu_for_1_slc_32_1_svs);
  assign Gelu_for_else_Gelu_for_else_mux1h_16_nl = MUX1HOT_v_5_4_2((signext_5_1(Gelu_for_1_else_if_acc_itm[3])),
      (signext_5_1(Gelu_for_1_else_else_if_mul_cmp_z[46])), (signext_5_2(Gelu_for_y_1_sva_4_27_22_1[5:4])),
      act_write_data_data_0_0_sva_30_26, {(~ Gelu_for_1_else_slc_32_svs) , Gelu_for_else_and_ssc_1
      , Gelu_for_else_else_else_and_ssc_1 , Gelu_for_else_else_else_and_1_ssc_1});
  assign Gelu_for_y_1_lpi_1_dfm_4_30_26 = Gelu_for_else_Gelu_for_else_mux1h_16_nl
      & (signext_5_1(~ Gelu_for_else_and_32_ssc_1)) & ({{4{Gelu_for_1_slc_32_1_svs}},
      Gelu_for_1_slc_32_1_svs});
  assign Gelu_for_else_Gelu_for_else_mux1h_48_nl = MUX1HOT_s_1_4_2((Gelu_for_1_else_if_acc_itm[3]),
      (Gelu_for_1_else_else_if_mul_cmp_z[46]), (Gelu_for_y_1_sva_4_27_22_1[3]), reg_act_write_data_data_0_0_2_ftd,
      {(~ Gelu_for_1_else_slc_32_svs) , Gelu_for_else_and_ssc_1 , Gelu_for_else_else_else_and_ssc_1
      , Gelu_for_else_else_else_and_1_ssc_1});
  assign Gelu_for_y_1_lpi_1_dfm_4_25 = Gelu_for_else_Gelu_for_else_mux1h_48_nl &
      (~ Gelu_for_else_and_32_ssc_1) & Gelu_for_1_slc_32_1_svs;
  assign Gelu_for_else_Gelu_for_else_mux1h_64_nl = MUX1HOT_v_3_5_2((Gelu_for_1_else_if_acc_itm[2:0]),
      (signext_3_1(Gelu_for_1_else_else_if_mul_cmp_z[46])), (Gelu_for_1_else_else_else_if_mul_cmp_z[48:46]),
      (Gelu_for_y_1_sva_4_27_22_1[2:0]), reg_act_write_data_data_0_0_2_ftd_1, {(~
      Gelu_for_1_else_slc_32_svs) , Gelu_for_else_and_ssc_1 , Gelu_for_else_and_32_ssc_1
      , Gelu_for_else_else_else_and_ssc_1 , Gelu_for_else_else_else_and_1_ssc_1});
  assign Gelu_for_y_1_lpi_1_dfm_4_24_22 = MUX_v_3_2_2(3'b000, Gelu_for_else_Gelu_for_else_mux1h_64_nl,
      Gelu_for_1_slc_32_1_svs);
  assign Silu_for_else_and_16_ssc_1 = (~ Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign Silu_for_else_else_else_and_17_ssc_1 = Gelu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
      & Gelu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Silu_for_else_and_17_m1c_mx1;
  assign Silu_for_else_and_18_ssc_1 = (~ Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign Silu_for_else_else_else_and_19_ssc_1 = Gelu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
      & Gelu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Silu_for_else_and_19_m1c_mx1;
  assign Silu_for_else_and_20_ssc_1 = (~ Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign Silu_for_else_else_else_and_21_ssc_1 = Gelu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
      & Gelu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Silu_for_else_and_21_m1c_mx1;
  assign Silu_for_else_and_22_ssc_1 = (~ Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign Silu_for_else_else_else_and_23_ssc_1 = Gelu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
      & Gelu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Silu_for_else_and_23_m1c_mx1;
  assign Silu_for_else_and_24_ssc_1 = (~ Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign Silu_for_else_else_else_and_25_ssc_1 = Gelu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
      & Gelu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Silu_for_else_and_25_m1c_mx1;
  assign Silu_for_else_and_26_ssc_1 = (~ Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign Silu_for_else_else_else_and_27_ssc_1 = Gelu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
      & Gelu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Silu_for_else_and_27_m1c_mx1;
  assign Silu_for_else_and_28_ssc_1 = (~ Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign Silu_for_else_else_else_and_29_ssc_1 = Gelu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
      & Gelu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Silu_for_else_and_29_m1c_mx1;
  assign Silu_for_else_and_30_ssc_1 = (~ Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs;
  assign Silu_for_else_else_else_and_31_ssc_1 = Gelu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
      & Gelu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Silu_for_else_and_31_m1c_mx1;
  assign Silu_for_else_and_47_ssc_1 = (~ Gelu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs)
      & Silu_for_else_and_31_m1c_mx1;
  assign Silu_for_else_else_else_and_30_ssc_1 = (~ Gelu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      & Gelu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Silu_for_else_and_31_m1c_mx1;
  assign Silu_for_else_and_46_ssc_1 = (~ Gelu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs)
      & Silu_for_else_and_29_m1c_mx1;
  assign Silu_for_else_else_else_and_28_ssc_1 = (~ Gelu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      & Gelu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Silu_for_else_and_29_m1c_mx1;
  assign Silu_for_else_and_45_ssc_1 = (~ Gelu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs)
      & Silu_for_else_and_27_m1c_mx1;
  assign Silu_for_else_else_else_and_26_ssc_1 = (~ Gelu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      & Gelu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Silu_for_else_and_27_m1c_mx1;
  assign Silu_for_else_and_44_ssc_1 = (~ Gelu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs)
      & Silu_for_else_and_25_m1c_mx1;
  assign Silu_for_else_else_else_and_24_ssc_1 = (~ Gelu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      & Gelu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Silu_for_else_and_25_m1c_mx1;
  assign Silu_for_else_and_43_ssc_1 = (~ Gelu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs)
      & Silu_for_else_and_23_m1c_mx1;
  assign Silu_for_else_else_else_and_22_ssc_1 = (~ Gelu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      & Gelu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Silu_for_else_and_23_m1c_mx1;
  assign Silu_for_else_and_42_ssc_1 = (~ Gelu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs)
      & Silu_for_else_and_21_m1c_mx1;
  assign Silu_for_else_else_else_and_20_ssc_1 = (~ Gelu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      & Gelu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Silu_for_else_and_21_m1c_mx1;
  assign Silu_for_else_and_41_ssc_1 = (~ Gelu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs)
      & Silu_for_else_and_19_m1c_mx1;
  assign Silu_for_else_else_else_and_18_ssc_1 = (~ Gelu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      & Gelu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Silu_for_else_and_19_m1c_mx1;
  assign Silu_for_else_and_40_ssc_1 = (~ Gelu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs)
      & Silu_for_else_and_17_m1c_mx1;
  assign Silu_for_else_else_else_and_16_ssc_1 = (~ Gelu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      & Gelu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Silu_for_else_and_17_m1c_mx1;
  assign nl_Gelu_for_y_1_sva_4_27_22_1 = conv_u2s_5_6(Gelu_for_1_else_else_else_if_mul_cmp_z[50:46])
      + 6'b111111;
  assign Gelu_for_y_1_sva_4_27_22_1 = nl_Gelu_for_y_1_sva_4_27_22_1[5:0];
  assign nl_Gelu_for_y_2_sva_4_27_22_1 = conv_u2s_5_6(Gelu_for_1_else_else_else_if_mul_cmp_15_z[50:46])
      + 6'b111111;
  assign Gelu_for_y_2_sva_4_27_22_1 = nl_Gelu_for_y_2_sva_4_27_22_1[5:0];
  assign nl_Gelu_for_y_3_sva_4_27_22_1 = conv_u2s_5_6(Gelu_for_1_else_else_else_if_mul_cmp_14_z[50:46])
      + 6'b111111;
  assign Gelu_for_y_3_sva_4_27_22_1 = nl_Gelu_for_y_3_sva_4_27_22_1[5:0];
  assign nl_Gelu_for_y_4_sva_4_27_22_1 = conv_u2s_5_6(Gelu_for_1_else_else_else_if_mul_cmp_13_z[50:46])
      + 6'b111111;
  assign Gelu_for_y_4_sva_4_27_22_1 = nl_Gelu_for_y_4_sva_4_27_22_1[5:0];
  assign nl_Gelu_for_y_5_sva_4_27_22_1 = conv_u2s_5_6(Gelu_for_1_else_else_else_if_mul_cmp_12_z[50:46])
      + 6'b111111;
  assign Gelu_for_y_5_sva_4_27_22_1 = nl_Gelu_for_y_5_sva_4_27_22_1[5:0];
  assign nl_Gelu_for_y_6_sva_4_27_22_1 = conv_u2s_5_6(Gelu_for_1_else_else_else_if_mul_cmp_11_z[50:46])
      + 6'b111111;
  assign Gelu_for_y_6_sva_4_27_22_1 = nl_Gelu_for_y_6_sva_4_27_22_1[5:0];
  assign nl_Gelu_for_y_7_sva_4_27_22_1 = conv_u2s_5_6(Gelu_for_1_else_else_else_if_mul_cmp_10_z[50:46])
      + 6'b111111;
  assign Gelu_for_y_7_sva_4_27_22_1 = nl_Gelu_for_y_7_sva_4_27_22_1[5:0];
  assign nl_Gelu_for_y_8_sva_4_27_22_1 = conv_u2s_5_6(Gelu_for_1_else_else_else_if_mul_cmp_9_z[50:46])
      + 6'b111111;
  assign Gelu_for_y_8_sva_4_27_22_1 = nl_Gelu_for_y_8_sva_4_27_22_1[5:0];
  assign nl_Gelu_for_y_9_sva_4_27_22_1 = conv_u2s_5_6(Gelu_for_1_else_else_else_if_mul_cmp_8_z[50:46])
      + 6'b111111;
  assign Gelu_for_y_9_sva_4_27_22_1 = nl_Gelu_for_y_9_sva_4_27_22_1[5:0];
  assign nl_Gelu_for_y_10_sva_4_27_22_1 = conv_u2s_5_6(Gelu_for_1_else_else_else_if_mul_cmp_7_z[50:46])
      + 6'b111111;
  assign Gelu_for_y_10_sva_4_27_22_1 = nl_Gelu_for_y_10_sva_4_27_22_1[5:0];
  assign nl_Gelu_for_y_11_sva_4_27_22_1 = conv_u2s_5_6(Gelu_for_1_else_else_else_if_mul_cmp_6_z[50:46])
      + 6'b111111;
  assign Gelu_for_y_11_sva_4_27_22_1 = nl_Gelu_for_y_11_sva_4_27_22_1[5:0];
  assign nl_Gelu_for_y_12_sva_4_27_22_1 = conv_u2s_5_6(Gelu_for_1_else_else_else_if_mul_cmp_5_z[50:46])
      + 6'b111111;
  assign Gelu_for_y_12_sva_4_27_22_1 = nl_Gelu_for_y_12_sva_4_27_22_1[5:0];
  assign nl_Gelu_for_y_13_sva_4_27_22_1 = conv_u2s_5_6(Gelu_for_1_else_else_else_if_mul_cmp_4_z[50:46])
      + 6'b111111;
  assign Gelu_for_y_13_sva_4_27_22_1 = nl_Gelu_for_y_13_sva_4_27_22_1[5:0];
  assign nl_Gelu_for_y_14_sva_4_27_22_1 = conv_u2s_5_6(Gelu_for_1_else_else_else_if_mul_cmp_3_z[50:46])
      + 6'b111111;
  assign Gelu_for_y_14_sva_4_27_22_1 = nl_Gelu_for_y_14_sva_4_27_22_1[5:0];
  assign nl_Gelu_for_y_15_sva_4_27_22_1 = conv_u2s_5_6(Gelu_for_1_else_else_else_if_mul_cmp_2_z[50:46])
      + 6'b111111;
  assign Gelu_for_y_15_sva_4_27_22_1 = nl_Gelu_for_y_15_sva_4_27_22_1[5:0];
  assign nl_Gelu_for_y_sva_4_27_22_1 = conv_u2s_5_6(Gelu_for_1_else_else_else_if_mul_cmp_1_z[50:46])
      + 6'b111111;
  assign Gelu_for_y_sva_4_27_22_1 = nl_Gelu_for_y_sva_4_27_22_1[5:0];
  assign Gelu_for_else_and_30_ssc_1 = (~ Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & Gelu_for_16_else_slc_32_svs;
  assign Gelu_for_else_else_else_and_30_ssc_1 = (~ Gelu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      & Gelu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_else_and_31_m1c_mx1;
  assign Gelu_for_else_and_47_ssc_1 = (~ Gelu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs)
      & Gelu_for_else_and_31_m1c_mx1;
  assign Gelu_for_else_else_else_and_31_ssc_1 = Gelu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
      & Gelu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_else_and_31_m1c_mx1;
  assign Gelu_for_else_and_28_ssc_1 = (~ Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & Gelu_for_15_else_slc_32_svs;
  assign Gelu_for_else_else_else_and_28_ssc_1 = (~ Gelu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      & Gelu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_else_and_29_m1c_mx1;
  assign Gelu_for_else_and_46_ssc_1 = (~ Gelu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs)
      & Gelu_for_else_and_29_m1c_mx1;
  assign Gelu_for_else_else_else_and_29_ssc_1 = Gelu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
      & Gelu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_else_and_29_m1c_mx1;
  assign Gelu_for_else_and_26_ssc_1 = (~ Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & Gelu_for_14_else_slc_32_svs;
  assign Gelu_for_else_else_else_and_26_ssc_1 = (~ Gelu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      & Gelu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_else_and_27_m1c_mx1;
  assign Gelu_for_else_and_45_ssc_1 = (~ Gelu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs)
      & Gelu_for_else_and_27_m1c_mx1;
  assign Gelu_for_else_else_else_and_27_ssc_1 = Gelu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
      & Gelu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_else_and_27_m1c_mx1;
  assign Gelu_for_else_and_24_ssc_1 = (~ Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & Gelu_for_13_else_slc_32_svs;
  assign Gelu_for_else_else_else_and_24_ssc_1 = (~ Gelu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      & Gelu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_else_and_25_m1c_mx1;
  assign Gelu_for_else_and_44_ssc_1 = (~ Gelu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs)
      & Gelu_for_else_and_25_m1c_mx1;
  assign Gelu_for_else_else_else_and_25_ssc_1 = Gelu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
      & Gelu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_else_and_25_m1c_mx1;
  assign Gelu_for_else_and_22_ssc_1 = (~ Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & Gelu_for_12_else_slc_32_svs;
  assign Gelu_for_else_else_else_and_22_ssc_1 = (~ Gelu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      & Gelu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_else_and_23_m1c_mx1;
  assign Gelu_for_else_and_43_ssc_1 = (~ Gelu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs)
      & Gelu_for_else_and_23_m1c_mx1;
  assign Gelu_for_else_else_else_and_23_ssc_1 = Gelu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
      & Gelu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_else_and_23_m1c_mx1;
  assign Gelu_for_else_and_20_ssc_1 = (~ Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & Gelu_for_11_else_slc_32_svs;
  assign Gelu_for_else_else_else_and_20_ssc_1 = (~ Gelu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      & Gelu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_else_and_21_m1c_mx1;
  assign Gelu_for_else_and_42_ssc_1 = (~ Gelu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs)
      & Gelu_for_else_and_21_m1c_mx1;
  assign Gelu_for_else_else_else_and_21_ssc_1 = Gelu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
      & Gelu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_else_and_21_m1c_mx1;
  assign Gelu_for_else_and_18_ssc_1 = (~ Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & Gelu_for_10_else_slc_32_svs;
  assign Gelu_for_else_else_else_and_18_ssc_1 = (~ Gelu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      & Gelu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_else_and_19_m1c_mx1;
  assign Gelu_for_else_and_41_ssc_1 = (~ Gelu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs)
      & Gelu_for_else_and_19_m1c_mx1;
  assign Gelu_for_else_else_else_and_19_ssc_1 = Gelu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
      & Gelu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_else_and_19_m1c_mx1;
  assign Gelu_for_else_and_16_ssc_1 = (~ Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
      & Gelu_for_9_else_slc_32_svs;
  assign Gelu_for_else_else_else_and_16_ssc_1 = (~ Gelu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      & Gelu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_else_and_17_m1c_mx1;
  assign Gelu_for_else_and_40_ssc_1 = (~ Gelu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs)
      & Gelu_for_else_and_17_m1c_mx1;
  assign Gelu_for_else_else_else_and_17_ssc_1 = Gelu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
      & Gelu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_else_and_17_m1c_mx1;
  assign Gelu_for_else_and_14_ssc_1 = (~ Gelu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs)
      & Gelu_for_8_else_slc_32_svs;
  assign Gelu_for_else_else_else_and_14_ssc_1 = (~ Gelu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      & Gelu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_else_and_15_m1c_mx1;
  assign Gelu_for_else_and_39_ssc_1 = (~ Gelu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs)
      & Gelu_for_else_and_15_m1c_mx1;
  assign Gelu_for_else_else_else_and_15_ssc_1 = Gelu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
      & Gelu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_else_and_15_m1c_mx1;
  assign Gelu_for_else_and_12_ssc_1 = (~ Gelu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs)
      & Gelu_for_7_else_slc_32_svs;
  assign Gelu_for_else_else_else_and_12_ssc_1 = (~ Gelu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      & Gelu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_else_and_13_m1c_mx1;
  assign Gelu_for_else_and_38_ssc_1 = (~ Gelu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs)
      & Gelu_for_else_and_13_m1c_mx1;
  assign Gelu_for_else_else_else_and_13_ssc_1 = Gelu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
      & Gelu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_else_and_13_m1c_mx1;
  assign Gelu_for_else_and_10_ssc_1 = (~ Gelu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs)
      & Gelu_for_6_else_slc_32_svs;
  assign Gelu_for_else_else_else_and_10_ssc_1 = (~ Gelu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      & Gelu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_else_and_11_m1c_mx1;
  assign Gelu_for_else_and_37_ssc_1 = (~ Gelu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs)
      & Gelu_for_else_and_11_m1c_mx1;
  assign Gelu_for_else_else_else_and_11_ssc_1 = Gelu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
      & Gelu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_else_and_11_m1c_mx1;
  assign Gelu_for_else_and_8_ssc_1 = (~ Gelu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs)
      & Gelu_for_5_else_slc_32_svs;
  assign Gelu_for_else_else_else_and_8_ssc_1 = (~ Gelu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      & Gelu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_else_and_9_m1c_mx1;
  assign Gelu_for_else_and_36_ssc_1 = (~ Gelu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs)
      & Gelu_for_else_and_9_m1c_mx1;
  assign Gelu_for_else_else_else_and_9_ssc_1 = Gelu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
      & Gelu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_else_and_9_m1c_mx1;
  assign Gelu_for_else_and_6_ssc_1 = (~ Gelu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs)
      & Gelu_for_4_else_slc_32_svs;
  assign Gelu_for_else_else_else_and_6_ssc_1 = (~ Gelu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      & Gelu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_else_and_7_m1c_mx1;
  assign Gelu_for_else_and_35_ssc_1 = (~ Gelu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs)
      & Gelu_for_else_and_7_m1c_mx1;
  assign Gelu_for_else_else_else_and_7_ssc_1 = Gelu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
      & Gelu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_else_and_7_m1c_mx1;
  assign Gelu_for_else_and_4_ssc_1 = (~ Gelu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs)
      & Gelu_for_3_else_slc_32_svs;
  assign Gelu_for_else_else_else_and_4_ssc_1 = (~ Gelu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      & Gelu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_else_and_5_m1c_mx1;
  assign Gelu_for_else_and_34_ssc_1 = (~ Gelu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs)
      & Gelu_for_else_and_5_m1c_mx1;
  assign Gelu_for_else_else_else_and_5_ssc_1 = Gelu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
      & Gelu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_else_and_5_m1c_mx1;
  assign Gelu_for_else_and_2_ssc_1 = (~ Gelu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs)
      & Gelu_for_2_else_slc_32_svs;
  assign Gelu_for_else_else_else_and_2_ssc_1 = (~ Gelu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      & Gelu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_else_and_3_m1c_mx1;
  assign Gelu_for_else_and_33_ssc_1 = (~ Gelu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs)
      & Gelu_for_else_and_3_m1c_mx1;
  assign Gelu_for_else_else_else_and_3_ssc_1 = Gelu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
      & Gelu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_else_and_3_m1c_mx1;
  assign Gelu_for_else_and_ssc_1 = (~ Gelu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs)
      & Gelu_for_1_else_slc_32_svs;
  assign Gelu_for_else_else_else_and_ssc_1 = (~ Gelu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs)
      & Gelu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_else_and_1_m1c_mx1;
  assign Gelu_for_else_and_32_ssc_1 = (~ Gelu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs)
      & Gelu_for_else_and_1_m1c_mx1;
  assign Gelu_for_else_else_else_and_1_ssc_1 = Gelu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
      & Gelu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
      & Gelu_for_else_and_1_m1c_mx1;
  assign while_nand_112_ssc_1 = ~(is_start_sva & while_nor_48_itm);
  assign ActUnit_RunInst_switch_lp_and_801_ssc_1 = ActUnit_CheckStart_start_reg_sva
      & ActUnit_RunInst_switch_lp_equal_tmp_2 & is_start_sva;
  assign ActUnit_RunInst_switch_lp_and_545_ssc_1 = reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_2_cse
      & ActUnit_RunInst_switch_lp_equal_tmp_4 & is_start_sva;
  assign ActUnit_RunInst_switch_lp_and_547_ssc_1 = reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_2_cse
      & ActUnit_RunInst_switch_lp_equal_tmp_5 & is_start_sva;
  assign ActUnit_RunInst_switch_lp_and_551_ssc_1 = reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_2_cse
      & ActUnit_RunInst_switch_lp_equal_tmp_7 & is_start_sva;
  assign ActUnit_RunInst_switch_lp_and_553_ssc_1 = Gelu_for_and_2_cse_sva & ActUnit_RunInst_switch_lp_equal_tmp_8
      & is_start_sva;
  assign ActUnit_RunInst_switch_lp_and_549_ssc_1 = reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_2_cse
      & ActUnit_RunInst_switch_lp_equal_tmp_6 & is_start_sva;
  assign while_nand_96_ssc_1 = ~(is_start_sva & while_nor_32_itm);
  assign ActUnit_RunInst_switch_lp_and_769_ssc_1 = ActUnit_RunInst_switch_lp_and_32_tmp
      & ActUnit_RunInst_switch_lp_equal_tmp_2 & is_start_sva;
  assign ActUnit_RunInst_switch_lp_and_385_ssc_1 = reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_cse
      & ActUnit_RunInst_switch_lp_equal_tmp_4 & is_start_sva;
  assign ActUnit_RunInst_switch_lp_and_387_ssc_1 = reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_cse
      & ActUnit_RunInst_switch_lp_equal_tmp_5 & is_start_sva;
  assign ActUnit_RunInst_switch_lp_and_391_ssc_1 = reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_cse
      & ActUnit_RunInst_switch_lp_equal_tmp_7 & is_start_sva;
  assign ActUnit_RunInst_switch_lp_and_393_ssc_1 = reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_cse
      & ActUnit_RunInst_switch_lp_equal_tmp_8 & is_start_sva;
  assign ActUnit_RunInst_switch_lp_and_389_ssc_1 = reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_cse
      & ActUnit_RunInst_switch_lp_equal_tmp_6 & is_start_sva;
  assign while_nand_80_ssc_1 = ~(is_start_sva & while_nor_16_itm);
  assign ActUnit_RunInst_switch_lp_and_737_ssc_1 = ActUnit_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva
      & ActUnit_RunInst_switch_lp_equal_tmp_2 & is_start_sva;
  assign ActUnit_RunInst_switch_lp_and_225_ssc_1 = reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_1_cse
      & ActUnit_RunInst_switch_lp_equal_tmp_4 & is_start_sva;
  assign ActUnit_RunInst_switch_lp_and_227_ssc_1 = reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_1_cse
      & ActUnit_RunInst_switch_lp_equal_tmp_5 & is_start_sva;
  assign ActUnit_RunInst_switch_lp_and_231_ssc_1 = reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_1_cse
      & ActUnit_RunInst_switch_lp_equal_tmp_7 & is_start_sva;
  assign ActUnit_RunInst_switch_lp_and_233_ssc_1 = ActUnit_PushOutput_if_for_and_stg_2_7_sva
      & ActUnit_RunInst_switch_lp_equal_tmp_8 & is_start_sva;
  assign ActUnit_RunInst_switch_lp_and_229_ssc_1 = reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_1_cse
      & ActUnit_RunInst_switch_lp_equal_tmp_6 & is_start_sva;
  assign while_nand_64_ssc_1 = ~(is_start_sva & while_nor_itm);
  assign ActUnit_RunInst_switch_lp_and_704_ssc_1 = ActUnit_RunInst_switch_lp_and_tmp
      & ActUnit_RunInst_switch_lp_equal_tmp_2 & is_start_sva;
  assign ActUnit_RunInst_switch_lp_and_65_ssc_1 = reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_nor_cse
      & ActUnit_RunInst_switch_lp_equal_tmp_4 & is_start_sva;
  assign ActUnit_RunInst_switch_lp_and_67_ssc_1 = reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_nor_cse
      & ActUnit_RunInst_switch_lp_equal_tmp_5 & is_start_sva;
  assign ActUnit_RunInst_switch_lp_and_71_ssc_1 = reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_nor_cse
      & ActUnit_RunInst_switch_lp_equal_tmp_7 & is_start_sva;
  assign ActUnit_RunInst_switch_lp_and_73_ssc_1 = reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_nor_cse
      & ActUnit_RunInst_switch_lp_equal_tmp_8 & is_start_sva;
  assign ActUnit_RunInst_switch_lp_and_69_ssc_1 = reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_nor_cse
      & ActUnit_RunInst_switch_lp_equal_tmp_6 & is_start_sva;
  assign ActUnit_PushOutput_if_for_and_27_seb_1 = ActUnit_PushOutput_if_for_and_stg_2_7_sva
      & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign nvhls_get_slc_2U_NVUINT8_return_3_sva_1 = MUX_v_2_32_2((act_config_inst_regs_0_sva_dfm_5[3:2]),
      (act_config_inst_regs_1_sva_dfm_5[3:2]), (act_config_inst_regs_2_sva_dfm_5[3:2]),
      (act_config_inst_regs_3_sva_dfm_5[3:2]), (act_config_inst_regs_4_sva_dfm_5[3:2]),
      (act_config_inst_regs_5_sva_dfm_5[3:2]), (act_config_inst_regs_6_sva_dfm_5[3:2]),
      (act_config_inst_regs_7_sva_dfm_5[3:2]), (act_config_inst_regs_8_sva_dfm_5[3:2]),
      (act_config_inst_regs_9_sva_dfm_5[3:2]), (act_config_inst_regs_10_sva_dfm_5[3:2]),
      (act_config_inst_regs_11_sva_dfm_5[3:2]), (act_config_inst_regs_12_sva_dfm_5[3:2]),
      (act_config_inst_regs_13_sva_dfm_5[3:2]), (act_config_inst_regs_14_sva_dfm_5[3:2]),
      (act_config_inst_regs_15_sva_dfm_5[3:2]), (act_config_inst_regs_16_sva_dfm_6[3:2]),
      (act_config_inst_regs_17_sva_dfm_6[3:2]), (act_config_inst_regs_18_sva_dfm_6[3:2]),
      (act_config_inst_regs_19_sva_dfm_6[3:2]), (act_config_inst_regs_20_sva_dfm_6[3:2]),
      (act_config_inst_regs_21_sva_dfm_6[3:2]), (act_config_inst_regs_22_sva_dfm_6[3:2]),
      (act_config_inst_regs_23_sva_dfm_6[3:2]), (act_config_inst_regs_24_sva_dfm_6[3:2]),
      (act_config_inst_regs_25_sva_dfm_6[3:2]), (act_config_inst_regs_26_sva_dfm_6[3:2]),
      (act_config_inst_regs_27_sva_dfm_6[3:2]), (act_config_inst_regs_28_sva_dfm_6[3:2]),
      (act_config_inst_regs_29_sva_dfm_6[3:2]), (act_config_inst_regs_30_sva_dfm_6[3:2]),
      (act_config_inst_regs_31_sva_dfm_6[3:2]), act_config_inst_counter_sva_dfm_3);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289 = ~((nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b11));
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_291 = (nvhls_get_slc_2U_NVUINT8_return_3_sva_1!=2'b00);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293 = ~((nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b10));
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295 = ~((nvhls_get_slc_2U_NVUINT8_return_3_sva_1==2'b01));
  assign ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1
      = MUX_v_32_16_2(act_port_read_out_data_0_0_sva_dfm, act_port_read_out_data_0_1_sva_dfm,
      act_port_read_out_data_0_2_sva_dfm, act_port_read_out_data_0_3_sva_dfm, act_port_read_out_data_0_4_sva_dfm,
      act_port_read_out_data_0_5_sva_dfm, act_port_read_out_data_0_6_sva_dfm, act_port_read_out_data_0_7_sva_dfm,
      act_port_read_out_data_0_8_sva_dfm, act_port_read_out_data_0_9_sva_dfm, act_port_read_out_data_0_10_sva_dfm,
      act_port_read_out_data_0_11_sva_dfm, act_port_read_out_data_0_12_sva_dfm, act_port_read_out_data_0_13_sva_dfm,
      act_port_read_out_data_0_14_sva_dfm, act_port_read_out_data_0_15_sva_dfm, ActUnit_PushOutput_if_for_i_4_0_sva_3_0);
  assign act_config_InstIncr_if_act_config_InstIncr_if_if_nor_tmp = ~((({reg_act_config_output_counter_sva_dfm_3_ftd
      , reg_act_config_output_counter_sva_dfm_3_ftd_1_3 , reg_act_config_output_counter_sva_dfm_3_ftd_1_2_0})
      != (operator_8_false_acc_sdt_sva_1[7:0])) | (operator_8_false_acc_sdt_sva_1[8]));
  assign nl_operator_8_false_acc_sdt_sva_1 = conv_u2s_8_9(act_config_num_output_sva)
      + 9'b111111111;
  assign operator_8_false_acc_sdt_sva_1 = nl_operator_8_false_acc_sdt_sva_1[8:0];
  assign nl_operator_6_false_acc_tmp = conv_u2s_6_7(act_config_num_inst_sva) + 7'b1111111;
  assign operator_6_false_acc_tmp = nl_operator_6_false_acc_tmp[6:0];
  assign while_nand_ssc_1 = ~(is_start_sva & w_load_lpi_1_dfm_1);
  assign ActUnit_RunLoad_and_ssc_1 = act_config_is_zero_first_sva_dfm_4 & w_load_lpi_1_dfm_1
      & is_start_sva;
  assign ActUnit_RunLoad_and_1_ssc_1 = (~ act_config_is_zero_first_sva_dfm_4) & w_load_lpi_1_dfm_1
      & is_start_sva;
  assign ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_and_1_nl
      = MUX_v_5_2_2(5'b00000, act_write_addrs_lpi_1_dfm_5, ActUnit_RunInst_switch_lp_and_32_tmp);
  assign while_mux_55_tmp = MUX_v_5_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_2_mx0w2,
      ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_and_1_nl,
      is_start_sva);
  assign nor_215_cse = ~((fsm_output[1:0]!=2'b00));
  assign and_dcpl_7 = is_start_sva & (act_config_in_InstFetch_return_sva_7_2[4]);
  assign and_dcpl_9 = and_dcpl_7 & (act_config_in_InstFetch_return_sva_7_2[3]) &
      (act_config_in_InstFetch_return_sva_7_2[5]) & ActUnit_RunInst_switch_lp_equal_tmp_7;
  assign and_dcpl_40 = ActUnit_RunInst_switch_lp_equal_tmp_7 & (~ (act_config_in_InstFetch_return_sva_7_2[2]));
  assign and_dcpl_43 = and_dcpl_7 & (act_config_in_InstFetch_return_sva_7_2[3]) &
      (act_config_in_InstFetch_return_sva_7_2[5]);
  assign or_tmp = reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_nor_cse
      | reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_1_cse | reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_cse
      | reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_2_cse;
  assign or_dcpl_28 = ActUnit_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva
      | is_start_sva;
  assign and_dcpl_78 = (act_config_in_InstFetch_mux_tmp[6]) & (act_config_in_InstFetch_mux_tmp[4]);
  assign and_dcpl_83 = is_start_sva & (act_config_in_InstFetch_mux_tmp[7]);
  assign and_dcpl_84 = and_dcpl_83 & (act_config_in_InstFetch_mux_tmp[5]);
  assign and_dcpl_86 = (act_config_in_InstFetch_mux_tmp[6]) & (~ (act_config_in_InstFetch_mux_tmp[4]));
  assign and_dcpl_117 = and_dcpl_84 & and_dcpl_86;
  assign and_dcpl_331 = and_2371_cse & nor_1441_cse;
  assign nor_222_cse = ~((~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[8])) | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11:9]!=3'b100));
  assign nor_221_nl = ~(is_start_sva | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[8]))
      | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11:9]!=3'b100));
  assign or_356_nl = is_start_sva | nor_222_cse;
  assign mux_101_nl = MUX_s_1_2_2(nor_221_nl, or_356_nl, ActUnit_RunInst_switch_lp_and_32_tmp);
  assign and_dcpl_332 = mux_101_nl & and_dcpl_331;
  assign and_dcpl_333 = is_start_sva & w_load_lpi_1_dfm_1;
  assign or_tmp_146 = is_start_sva | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[8]))
      | rva_in_PopNB_mioi_data_rw_rsc_z_mxwt | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11:9]!=3'b100);
  assign nor_224_nl = ~((~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[8])) | rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11:9]!=3'b100));
  assign mux_114_nl = MUX_s_1_2_2(nor_224_nl, ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_2_tmp,
      is_start_sva);
  assign not_tmp_237 = MUX_s_1_2_2(mux_114_nl, (~ or_tmp_146), ActUnit_RunInst_switch_lp_and_32_tmp);
  assign and_dcpl_337 = not_tmp_237 & and_dcpl_331;
  assign or_tmp_158 = (act_config_in_InstFetch_return_sva_7_2[2]) | ActUnit_RunInst_switch_lp_equal_tmp_7;
  assign mux_tmp_108 = MUX_s_1_2_2(ActUnit_RunInst_switch_lp_equal_tmp_7, ActUnit_RunInst_switch_lp_equal_tmp_8,
      act_config_in_InstFetch_return_sva_7_2[2]);
  assign and_dcpl_469 = is_start_sva & ActUnit_RunInst_switch_lp_equal_tmp_3;
  assign or_tmp_397 = is_start_sva | (~ ActUnit_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva);
  assign or_dcpl_450 = (act_config_in_InstFetch_mux_tmp[4]) | (~ is_start_sva);
  assign and_dcpl_846 = (fsm_output[1:0]==2'b01);
  assign and_dcpl_847 = and_dcpl_846 & nor_1441_cse;
  assign and_dcpl_848 = (fsm_output[1:0]==2'b10);
  assign and_dcpl_849 = and_dcpl_848 & nor_1441_cse;
  assign and_dcpl_852 = (fsm_output[0]) & (~ (act_config_in_InstFetch_return_sva_7_2[2]))
      & (fsm_output[1]) & nor_1441_cse;
  assign and_dcpl_855 = (fsm_output[0]) & (act_config_in_InstFetch_return_sva_7_2[2])
      & (fsm_output[1]) & nor_1441_cse;
  assign or_dcpl_457 = (fsm_output[3:2]!=2'b00);
  assign and_dcpl_856 = is_start_sva & (~ (fsm_output[3]));
  assign or_tmp_409 = (~ (fsm_output[0])) | (fsm_output[2]);
  assign or_870_nl = operator_32_8_true_AC_TRN_AC_WRAP_1_less_14_tmp | (~ operator_32_8_true_AC_TRN_AC_WRAP_less_14_tmp)
      | (act_config_in_InstFetch_mux_tmp[7:5]!=3'b111) | (fsm_output[2]);
  assign or_869_nl = Gelu_for_else_if_less_15_tmp | (~ Gelu_for_if_less_15_tmp) |
      (act_config_in_InstFetch_mux_tmp[7:5]!=3'b111) | (fsm_output[2]);
  assign mux_tmp_315 = MUX_s_1_2_2(or_870_nl, or_869_nl, act_config_in_InstFetch_mux_tmp[4]);
  assign mux_332_nl = MUX_s_1_2_2((~ (fsm_output[2])), mux_tmp_315, fsm_output[0]);
  assign mux_tmp_317 = MUX_s_1_2_2(mux_332_nl, or_tmp_409, fsm_output[1]);
  assign nand_22_nl = ~((fsm_output[0]) & (~ mux_tmp_315));
  assign mux_tmp_318 = MUX_s_1_2_2(nand_22_nl, or_tmp_409, fsm_output[1]);
  assign nand_tmp_23 = (fsm_output[1:0]!=2'b01) | mux_tmp_315;
  assign or_875_nl = operator_32_8_true_AC_TRN_AC_WRAP_1_less_13_tmp | (~ operator_32_8_true_AC_TRN_AC_WRAP_less_13_tmp)
      | (act_config_in_InstFetch_mux_tmp[7:5]!=3'b111) | (fsm_output[2]);
  assign or_874_nl = Gelu_for_else_if_less_13_tmp | (~ Gelu_for_if_less_13_tmp) |
      (act_config_in_InstFetch_mux_tmp[7:5]!=3'b111) | (fsm_output[2]);
  assign mux_tmp_325 = MUX_s_1_2_2(or_875_nl, or_874_nl, act_config_in_InstFetch_mux_tmp[4]);
  assign mux_342_nl = MUX_s_1_2_2((~ (fsm_output[2])), mux_tmp_325, fsm_output[0]);
  assign mux_tmp_327 = MUX_s_1_2_2(mux_342_nl, or_tmp_409, fsm_output[1]);
  assign nand_24_nl = ~((fsm_output[0]) & (~ mux_tmp_325));
  assign mux_tmp_328 = MUX_s_1_2_2(nand_24_nl, or_tmp_409, fsm_output[1]);
  assign nand_tmp_25 = (fsm_output[1:0]!=2'b01) | mux_tmp_325;
  assign or_880_nl = operator_32_8_true_AC_TRN_AC_WRAP_1_less_12_tmp | (~ operator_32_8_true_AC_TRN_AC_WRAP_less_12_tmp)
      | (act_config_in_InstFetch_mux_tmp[7:5]!=3'b111) | (fsm_output[2]);
  assign or_879_nl = Gelu_for_else_if_less_12_tmp | (~ Gelu_for_if_less_12_tmp) |
      (act_config_in_InstFetch_mux_tmp[7:5]!=3'b111) | (fsm_output[2]);
  assign mux_tmp_335 = MUX_s_1_2_2(or_880_nl, or_879_nl, act_config_in_InstFetch_mux_tmp[4]);
  assign mux_352_nl = MUX_s_1_2_2((~ (fsm_output[2])), mux_tmp_335, fsm_output[0]);
  assign mux_tmp_337 = MUX_s_1_2_2(mux_352_nl, or_tmp_409, fsm_output[1]);
  assign nand_26_nl = ~((fsm_output[0]) & (~ mux_tmp_335));
  assign mux_tmp_338 = MUX_s_1_2_2(nand_26_nl, or_tmp_409, fsm_output[1]);
  assign nand_tmp_27 = (fsm_output[1:0]!=2'b01) | mux_tmp_335;
  assign or_885_nl = operator_32_8_true_AC_TRN_AC_WRAP_1_less_11_tmp | (~ operator_32_8_true_AC_TRN_AC_WRAP_less_11_tmp)
      | (act_config_in_InstFetch_mux_tmp[7:5]!=3'b111) | (fsm_output[2]);
  assign or_884_nl = Gelu_for_else_if_less_11_tmp | (~ Gelu_for_if_less_11_tmp) |
      (act_config_in_InstFetch_mux_tmp[7:5]!=3'b111) | (fsm_output[2]);
  assign mux_tmp_345 = MUX_s_1_2_2(or_885_nl, or_884_nl, act_config_in_InstFetch_mux_tmp[4]);
  assign mux_362_nl = MUX_s_1_2_2((~ (fsm_output[2])), mux_tmp_345, fsm_output[0]);
  assign mux_tmp_347 = MUX_s_1_2_2(mux_362_nl, or_tmp_409, fsm_output[1]);
  assign nand_28_nl = ~((fsm_output[0]) & (~ mux_tmp_345));
  assign mux_tmp_348 = MUX_s_1_2_2(nand_28_nl, or_tmp_409, fsm_output[1]);
  assign nand_tmp_29 = (fsm_output[1:0]!=2'b01) | mux_tmp_345;
  assign or_890_nl = operator_32_8_true_AC_TRN_AC_WRAP_1_less_10_tmp | (~ operator_32_8_true_AC_TRN_AC_WRAP_less_10_tmp)
      | (act_config_in_InstFetch_mux_tmp[7:5]!=3'b111) | (fsm_output[2]);
  assign or_889_nl = Gelu_for_else_if_less_10_tmp | (~ Gelu_for_if_less_10_tmp) |
      (act_config_in_InstFetch_mux_tmp[7:5]!=3'b111) | (fsm_output[2]);
  assign mux_tmp_355 = MUX_s_1_2_2(or_890_nl, or_889_nl, act_config_in_InstFetch_mux_tmp[4]);
  assign mux_372_nl = MUX_s_1_2_2((~ (fsm_output[2])), mux_tmp_355, fsm_output[0]);
  assign mux_tmp_357 = MUX_s_1_2_2(mux_372_nl, or_tmp_409, fsm_output[1]);
  assign nand_30_nl = ~((fsm_output[0]) & (~ mux_tmp_355));
  assign mux_tmp_358 = MUX_s_1_2_2(nand_30_nl, or_tmp_409, fsm_output[1]);
  assign nand_tmp_31 = (fsm_output[1:0]!=2'b01) | mux_tmp_355;
  assign or_895_nl = operator_32_8_true_AC_TRN_AC_WRAP_1_less_9_tmp | (~ operator_32_8_true_AC_TRN_AC_WRAP_less_9_tmp)
      | (act_config_in_InstFetch_mux_tmp[7:5]!=3'b111) | (fsm_output[2]);
  assign or_894_nl = Gelu_for_else_if_less_9_tmp | (~ Gelu_for_if_less_9_tmp) | (act_config_in_InstFetch_mux_tmp[7:5]!=3'b111)
      | (fsm_output[2]);
  assign mux_tmp_365 = MUX_s_1_2_2(or_895_nl, or_894_nl, act_config_in_InstFetch_mux_tmp[4]);
  assign mux_382_nl = MUX_s_1_2_2((~ (fsm_output[2])), mux_tmp_365, fsm_output[0]);
  assign mux_tmp_367 = MUX_s_1_2_2(mux_382_nl, or_tmp_409, fsm_output[1]);
  assign nand_32_nl = ~((fsm_output[0]) & (~ mux_tmp_365));
  assign mux_tmp_368 = MUX_s_1_2_2(nand_32_nl, or_tmp_409, fsm_output[1]);
  assign nand_tmp_33 = (fsm_output[1:0]!=2'b01) | mux_tmp_365;
  assign or_900_nl = operator_32_8_true_AC_TRN_AC_WRAP_1_less_8_tmp | (~ operator_32_8_true_AC_TRN_AC_WRAP_less_8_tmp)
      | (act_config_in_InstFetch_mux_tmp[7:5]!=3'b111) | (fsm_output[2]);
  assign or_899_nl = Gelu_for_else_if_less_8_tmp | (~ Gelu_for_if_less_8_tmp) | (act_config_in_InstFetch_mux_tmp[7:5]!=3'b111)
      | (fsm_output[2]);
  assign mux_tmp_375 = MUX_s_1_2_2(or_900_nl, or_899_nl, act_config_in_InstFetch_mux_tmp[4]);
  assign mux_392_nl = MUX_s_1_2_2((~ (fsm_output[2])), mux_tmp_375, fsm_output[0]);
  assign mux_tmp_377 = MUX_s_1_2_2(mux_392_nl, or_tmp_409, fsm_output[1]);
  assign nand_34_nl = ~((fsm_output[0]) & (~ mux_tmp_375));
  assign mux_tmp_378 = MUX_s_1_2_2(nand_34_nl, or_tmp_409, fsm_output[1]);
  assign nand_tmp_35 = (fsm_output[1:0]!=2'b01) | mux_tmp_375;
  assign or_905_nl = operator_32_8_true_AC_TRN_AC_WRAP_1_less_15_tmp | (~ operator_32_8_true_AC_TRN_AC_WRAP_less_15_tmp)
      | (act_config_in_InstFetch_mux_tmp[7:5]!=3'b111) | (fsm_output[2]);
  assign or_904_nl = Gelu_for_else_if_less_14_tmp | (~ Gelu_for_if_less_14_tmp) |
      (act_config_in_InstFetch_mux_tmp[7:5]!=3'b111) | (fsm_output[2]);
  assign mux_tmp_385 = MUX_s_1_2_2(or_905_nl, or_904_nl, act_config_in_InstFetch_mux_tmp[4]);
  assign mux_402_nl = MUX_s_1_2_2((~ (fsm_output[2])), mux_tmp_385, fsm_output[0]);
  assign mux_tmp_387 = MUX_s_1_2_2(mux_402_nl, or_tmp_409, fsm_output[1]);
  assign nand_36_nl = ~((fsm_output[0]) & (~ mux_tmp_385));
  assign mux_tmp_388 = MUX_s_1_2_2(nand_36_nl, or_tmp_409, fsm_output[1]);
  assign nand_tmp_37 = (fsm_output[1:0]!=2'b01) | mux_tmp_385;
  assign and_dcpl_867 = is_start_sva & (act_config_in_InstFetch_return_sva_7_2[2]);
  assign not_tmp_445 = MUX_s_1_2_2(and_2371_cse, (~ or_1872_cse), fsm_output[2]);
  assign and_dcpl_872 = not_tmp_445 & and_1648_cse;
  assign and_dcpl_953 = (act_config_in_InstFetch_return_sva_7_2[3]) & (act_config_in_InstFetch_return_sva_7_2[5])
      & and_dcpl_867;
  assign and_dcpl_1048 = (fsm_output[2:1]==2'b01);
  assign and_dcpl_1051 = is_start_sva & (~ (fsm_output[0]));
  assign and_dcpl_1056 = (fsm_output[2:1]==2'b11);
  assign and_dcpl_1061 = (fsm_output[3:2]==2'b01);
  assign and_dcpl_1062 = ~(is_start_sva | (fsm_output[0]));
  assign and_dcpl_1063 = and_dcpl_1062 & (~ (fsm_output[1]));
  assign and_dcpl_1072 = (~ is_start_sva) & (fsm_output[0]);
  assign and_dcpl_1077 = and_2371_cse & (~ (fsm_output[2]));
  assign and_dcpl_1081 = (fsm_output[3:2]==2'b10);
  assign and_dcpl_1082 = and_dcpl_1051 & (fsm_output[1]);
  assign and_dcpl_1083 = and_dcpl_1082 & and_dcpl_1081;
  assign and_dcpl_1085 = and_dcpl_1062 & (fsm_output[1]) & and_dcpl_1081;
  assign or_dcpl_462 = is_start_sva | (~ (fsm_output[0]));
  assign or_dcpl_464 = or_dcpl_462 | (~ (fsm_output[1])) | or_dcpl_457;
  assign or_dcpl_465 = (~ rva_in_PopNB_mioi_return_rsc_z_mxwt) | rva_in_PopNB_mioi_data_rw_rsc_z_mxwt;
  assign and_dcpl_1088 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11:8]==4'b1000);
  assign or_dcpl_466 = and_dcpl_1088 | or_dcpl_465;
  assign or_dcpl_468 = ~(rva_in_PopNB_mioi_return_rsc_z_mxwt & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt);
  assign or_dcpl_469 = and_dcpl_1088 | or_dcpl_468;
  assign nor_320_cse = ~((fsm_output[2:1]!=2'b00));
  assign and_dcpl_1090 = nor_320_cse & (fsm_output[3]);
  assign or_dcpl_475 = (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[8])
      | is_start_sva | (~ and_2371_cse);
  assign or_dcpl_485 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[9])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[10]) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt);
  assign or_dcpl_487 = (fsm_output[2:1]!=2'b01);
  assign or_tmp_484 = (fsm_output[1:0]!=2'b01);
  assign mux_428_nl = MUX_s_1_2_2(and_2371_cse, or_tmp_484, fsm_output[2]);
  assign mux_tmp_413 = MUX_s_1_2_2((~ mux_428_nl), or_3395_cse, fsm_output[3]);
  assign and_dcpl_1093 = and_dcpl_848 & (~ (fsm_output[2]));
  assign and_dcpl_1094 = and_dcpl_1093 & (fsm_output[3]) & w_axi_rsp_lpi_1_dfm_1
      & act_read_req_valid_lpi_1_dfm_6;
  assign and_dcpl_1096 = and_dcpl_1093 & (~(act_read_req_valid_lpi_1_dfm_6 & w_axi_rsp_lpi_1_dfm_1))
      & (fsm_output[3]);
  assign or_tmp_485 = (fsm_output[2]) | and_2371_cse;
  assign not_tmp_495 = MUX_s_1_2_2((fsm_output[2]), (~ or_3395_cse), fsm_output[3]);
  assign or_dcpl_492 = (while_mux_55_tmp[1:0]!=2'b00);
  assign or_dcpl_493 = (while_mux_55_tmp[3:2]!=2'b00);
  assign or_dcpl_494 = or_dcpl_493 | or_dcpl_492;
  assign or_dcpl_496 = or_dcpl_487 | (fsm_output[3]) | (while_mux_55_tmp[4]);
  assign mux_434_nl = MUX_s_1_2_2(nor_222_cse, ActUnit_RunInst_switch_lp_and_32_tmp,
      is_start_sva);
  assign or_dcpl_498 = ~(mux_434_nl & (fsm_output[0]));
  assign or_dcpl_500 = (while_mux_55_tmp[1:0]!=2'b01);
  assign or_dcpl_501 = or_dcpl_493 | or_dcpl_500;
  assign or_dcpl_504 = (while_mux_55_tmp[1:0]!=2'b10);
  assign or_dcpl_505 = or_dcpl_493 | or_dcpl_504;
  assign or_dcpl_508 = ~((while_mux_55_tmp[1:0]==2'b11));
  assign or_dcpl_509 = or_dcpl_493 | or_dcpl_508;
  assign or_dcpl_512 = (while_mux_55_tmp[3:2]!=2'b01);
  assign or_dcpl_513 = or_dcpl_512 | or_dcpl_492;
  assign or_dcpl_516 = or_dcpl_512 | or_dcpl_500;
  assign or_dcpl_519 = or_dcpl_512 | or_dcpl_504;
  assign or_dcpl_522 = or_dcpl_512 | or_dcpl_508;
  assign or_dcpl_525 = (while_mux_55_tmp[3:2]!=2'b10);
  assign or_dcpl_526 = or_dcpl_525 | or_dcpl_492;
  assign or_dcpl_529 = or_dcpl_525 | or_dcpl_500;
  assign or_dcpl_532 = or_dcpl_525 | or_dcpl_504;
  assign or_dcpl_535 = or_dcpl_525 | or_dcpl_508;
  assign or_dcpl_538 = ~((while_mux_55_tmp[3:2]==2'b11));
  assign or_dcpl_539 = or_dcpl_538 | or_dcpl_492;
  assign or_dcpl_542 = or_dcpl_538 | or_dcpl_500;
  assign or_dcpl_545 = or_dcpl_538 | or_dcpl_504;
  assign or_dcpl_548 = or_dcpl_538 | or_dcpl_508;
  assign or_dcpl_552 = or_dcpl_487 | (fsm_output[3]) | (~ (while_mux_55_tmp[4]));
  assign not_tmp_503 = ~((ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_23_4_mx1_tmp_7_0==8'b00000011)
      & act_config_ActConfigRead_else_unequal_tmp_1 & act_config_ActConfigRead_unequal_tmp_1
      & (~ ActUnit_DecodeAxiRead_unequal_tmp_1) & ActUnit_DecodeAxi_rva_in_reg_rw_sva_mx1
      & ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_mx1
      & (~ is_start_sva));
  assign or_dcpl_586 = (~ and_2371_cse) | (fsm_output[2]);
  assign and_dcpl_1104 = and_dcpl_848 & and_dcpl_1081;
  assign and_dcpl_1106 = (~ (fsm_output[3])) & act_read_req_valid_lpi_1_dfm_6;
  assign and_dcpl_1109 = nor_215_cse & (fsm_output[2]);
  assign and_dcpl_1112 = nor_215_cse & and_dcpl_1061;
  assign or_dcpl_593 = ~(is_start_sva & (act_config_in_InstFetch_return_sva_7_2[2]));
  assign or_dcpl_595 = ~((act_config_in_InstFetch_return_sva_7_2[4:3]==2'b11));
  assign or_dcpl_596 = or_dcpl_595 | (~ (act_config_in_InstFetch_return_sva_7_2[5]));
  assign or_dcpl_616 = or_dcpl_595 | (~((act_config_in_InstFetch_return_sva_7_2[5])
      & is_start_sva));
  assign or_dcpl_622 = ~((act_config_in_InstFetch_mux_tmp[7:5]==3'b111));
  assign or_dcpl_623 = or_dcpl_622 | or_dcpl_450;
  assign and_dcpl_1116 = and_1648_cse & and_dcpl_1051;
  assign and_dcpl_1118 = ~((act_config_in_InstFetch_return_sva_7_2[2]) | (fsm_output[1]));
  assign or_dcpl_717 = or_dcpl_622 | (~((act_config_in_InstFetch_mux_tmp[4]) & is_start_sva));
  assign and_dcpl_1143 = is_start_sva & (fsm_output[0]);
  assign and_dcpl_1144 = and_1648_cse & and_dcpl_1143;
  assign and_dcpl_1174 = (act_config_in_InstFetch_return_sva_7_2[2]) & (~ (fsm_output[1]));
  assign and_dcpl_1228 = and_dcpl_1048 & (~ (fsm_output[3]));
  assign and_dcpl_1233 = and_dcpl_1072 & (fsm_output[1]) & nor_1441_cse;
  assign and_dcpl_1235 = and_dcpl_848 & and_dcpl_1061;
  assign and_dcpl_1236 = and_2371_cse & and_dcpl_1061;
  assign or_dcpl_815 = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1:0]!=2'b00);
  assign or_dcpl_817 = or_1726_cse | or_dcpl_815;
  assign or_dcpl_822 = (~((fsm_output[1]) ^ (fsm_output[0]))) | or_dcpl_457;
  assign or_dcpl_823 = or_tmp_484 | or_dcpl_457;
  assign and_dcpl_1240 = not_tmp_445 & (~ (fsm_output[3]));
  assign or_dcpl_824 = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1:0]!=2'b10);
  assign or_dcpl_825 = ~((ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3:2]==2'b11));
  assign or_dcpl_826 = or_dcpl_825 | or_dcpl_824;
  assign or_dcpl_827 = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1:0]!=2'b01);
  assign or_dcpl_828 = or_1726_cse | or_dcpl_827;
  assign or_dcpl_829 = or_dcpl_825 | or_dcpl_827;
  assign or_dcpl_830 = or_1726_cse | or_dcpl_824;
  assign or_dcpl_831 = or_dcpl_825 | or_dcpl_815;
  assign or_dcpl_833 = or_1726_cse | nand_533_cse;
  assign or_dcpl_835 = or_1738_cse | nand_533_cse;
  assign or_dcpl_836 = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3:2]!=2'b01);
  assign or_dcpl_837 = or_dcpl_836 | or_dcpl_815;
  assign or_dcpl_838 = or_1738_cse | or_dcpl_824;
  assign or_dcpl_839 = or_dcpl_836 | or_dcpl_827;
  assign or_dcpl_840 = or_1738_cse | or_dcpl_827;
  assign or_dcpl_841 = or_dcpl_836 | or_dcpl_824;
  assign or_dcpl_842 = or_1738_cse | or_dcpl_815;
  assign or_dcpl_843 = or_dcpl_836 | nand_533_cse;
  assign and_dcpl_1244 = and_dcpl_846 & and_dcpl_1061;
  assign and_dcpl_1246 = and_dcpl_846 & and_dcpl_1081;
  assign and_dcpl_1257 = (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7:0]==8'b00000010);
  assign and_dcpl_1262 = (or_dcpl_468 | is_start_sva) & (fsm_output[0]) & and_dcpl_1228;
  assign nand_252_nl = ~((fsm_output[2]) & or_1872_cse);
  assign mux_448_itm = MUX_s_1_2_2(nand_252_nl, or_3395_cse, fsm_output[3]);
  assign mux_tmp_433 = MUX_s_1_2_2((~ and_dcpl_1056), or_3395_cse, fsm_output[3]);
  assign or_dcpl_846 = ~((ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2:1]==2'b11));
  assign or_dcpl_847 = or_dcpl_846 | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]));
  assign or_dcpl_848 = ~((nvhls_get_slc_2U_NVUINT8_return_3_sva==2'b11));
  assign or_dcpl_849 = or_dcpl_848 | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]));
  assign or_dcpl_850 = or_dcpl_849 | or_dcpl_847;
  assign or_dcpl_851 = or_dcpl_846 | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]);
  assign or_dcpl_852 = or_dcpl_849 | or_dcpl_851;
  assign or_dcpl_853 = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2:1]!=2'b10);
  assign or_dcpl_854 = or_dcpl_853 | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]));
  assign or_dcpl_855 = or_dcpl_849 | or_dcpl_854;
  assign or_dcpl_856 = or_dcpl_853 | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]);
  assign or_dcpl_857 = or_dcpl_849 | or_dcpl_856;
  assign or_dcpl_858 = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2:1]!=2'b01);
  assign or_dcpl_859 = or_dcpl_858 | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]));
  assign or_dcpl_860 = or_dcpl_849 | or_dcpl_859;
  assign or_dcpl_861 = or_dcpl_858 | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]);
  assign or_dcpl_862 = or_dcpl_849 | or_dcpl_861;
  assign or_dcpl_863 = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2:1]!=2'b00);
  assign or_dcpl_864 = or_dcpl_863 | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]));
  assign or_dcpl_865 = or_dcpl_849 | or_dcpl_864;
  assign or_dcpl_866 = or_dcpl_863 | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]);
  assign or_dcpl_867 = or_dcpl_849 | or_dcpl_866;
  assign or_dcpl_868 = or_dcpl_848 | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign or_dcpl_869 = or_dcpl_868 | or_dcpl_847;
  assign or_dcpl_870 = or_dcpl_868 | or_dcpl_851;
  assign or_dcpl_871 = or_dcpl_868 | or_dcpl_854;
  assign or_dcpl_872 = or_dcpl_868 | or_dcpl_856;
  assign or_dcpl_873 = or_dcpl_868 | or_dcpl_859;
  assign or_dcpl_874 = or_dcpl_868 | or_dcpl_861;
  assign or_dcpl_875 = or_dcpl_868 | or_dcpl_864;
  assign or_tmp_490 = (fsm_output[2:0]!=3'b000);
  assign nand_39_nl = ~((fsm_output[2]) & (~ and_2371_cse));
  assign mux_450_itm = MUX_s_1_2_2(nand_39_nl, or_tmp_490, fsm_output[3]);
  assign and_dcpl_1264 = ~((ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2:1]!=2'b00));
  assign and_dcpl_1265 = and_dcpl_1264 & (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]));
  assign and_dcpl_1266 = (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]) & (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]));
  assign and_dcpl_1267 = (~ act_config_is_zero_first_sva_dfm_4) & (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]);
  assign and_dcpl_1270 = ~((~(or_dcpl_868 | or_dcpl_866)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1271 = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2:1]==2'b11);
  assign and_dcpl_1272 = and_dcpl_1271 & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]);
  assign and_dcpl_1274 = ~(act_config_is_zero_first_sva_dfm_4 | (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]));
  assign and_dcpl_1275 = and_dcpl_1274 & (nvhls_get_slc_2U_NVUINT8_return_3_sva[1])
      & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign or_dcpl_877 = (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b10);
  assign or_dcpl_878 = or_dcpl_877 | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]));
  assign and_dcpl_1277 = ~((~(or_dcpl_878 | or_dcpl_847)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1278 = and_dcpl_1271 & (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]));
  assign and_dcpl_1280 = ~((~(or_dcpl_878 | or_dcpl_851)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1281 = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2:1]==2'b10);
  assign and_dcpl_1282 = and_dcpl_1281 & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]);
  assign and_dcpl_1284 = ~((~(or_dcpl_878 | or_dcpl_854)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1285 = and_dcpl_1281 & (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]));
  assign and_dcpl_1287 = ~((~(or_dcpl_878 | or_dcpl_856)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1288 = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2:1]==2'b01);
  assign and_dcpl_1289 = and_dcpl_1288 & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]);
  assign and_dcpl_1291 = ~((~(or_dcpl_878 | or_dcpl_859)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1292 = and_dcpl_1288 & (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]));
  assign and_dcpl_1294 = ~((~(or_dcpl_878 | or_dcpl_861)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1295 = and_dcpl_1264 & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0]);
  assign and_dcpl_1297 = ~((~(or_dcpl_878 | or_dcpl_864)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1299 = ~((~(or_dcpl_878 | or_dcpl_866)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1300 = and_dcpl_1274 & and_dcpl_1266;
  assign or_dcpl_887 = or_dcpl_877 | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign and_dcpl_1302 = ~((~(or_dcpl_887 | or_dcpl_847)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1304 = ~((~(or_dcpl_887 | or_dcpl_851)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1306 = ~((~(or_dcpl_887 | or_dcpl_854)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1308 = ~((~(or_dcpl_887 | or_dcpl_856)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1310 = ~((~(or_dcpl_887 | or_dcpl_859)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1312 = ~((~(or_dcpl_887 | or_dcpl_861)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1314 = ~((~(or_dcpl_887 | or_dcpl_864)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1316 = ~((~(or_dcpl_887 | or_dcpl_866)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1317 = (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[1])) & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign and_dcpl_1318 = and_dcpl_1267 & and_dcpl_1317;
  assign or_dcpl_896 = (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b01);
  assign or_dcpl_897 = or_dcpl_896 | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]));
  assign and_dcpl_1320 = ~((~(or_dcpl_897 | or_dcpl_847)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1322 = ~((~(or_dcpl_897 | or_dcpl_851)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1324 = ~((~(or_dcpl_897 | or_dcpl_854)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1326 = ~((~(or_dcpl_897 | or_dcpl_856)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1328 = ~((~(or_dcpl_897 | or_dcpl_859)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1330 = ~((~(or_dcpl_897 | or_dcpl_861)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1332 = ~((~(or_dcpl_897 | or_dcpl_864)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1334 = ~((~(or_dcpl_897 | or_dcpl_866)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1335 = ~((nvhls_get_slc_2U_NVUINT8_return_3_sva[1]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]));
  assign and_dcpl_1336 = and_dcpl_1267 & and_dcpl_1335;
  assign or_dcpl_906 = or_dcpl_896 | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign and_dcpl_1338 = ~((~(or_dcpl_906 | or_dcpl_847)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1340 = ~((~(or_dcpl_906 | or_dcpl_851)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1342 = ~((~(or_dcpl_906 | or_dcpl_854)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1344 = ~((~(or_dcpl_906 | or_dcpl_856)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1346 = ~((~(or_dcpl_906 | or_dcpl_859)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1348 = ~((~(or_dcpl_906 | or_dcpl_861)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1350 = ~((~(or_dcpl_906 | or_dcpl_864)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1352 = ~((~(or_dcpl_906 | or_dcpl_866)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1353 = and_dcpl_1274 & and_dcpl_1317;
  assign or_dcpl_915 = (nvhls_get_slc_2U_NVUINT8_return_3_sva!=2'b00);
  assign or_dcpl_916 = or_dcpl_915 | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]));
  assign and_dcpl_1355 = ~((~(or_dcpl_916 | or_dcpl_847)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1357 = ~((~(or_dcpl_916 | or_dcpl_851)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1359 = ~((~(or_dcpl_916 | or_dcpl_854)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1361 = ~((~(or_dcpl_916 | or_dcpl_856)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1363 = ~((~(or_dcpl_916 | or_dcpl_859)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1365 = ~((~(or_dcpl_916 | or_dcpl_861)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1367 = ~((~(or_dcpl_916 | or_dcpl_864)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1369 = ~((~(or_dcpl_916 | or_dcpl_866)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1370 = and_dcpl_1274 & and_dcpl_1335;
  assign or_dcpl_925 = or_dcpl_915 | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign and_dcpl_1372 = ~((~(or_dcpl_925 | or_dcpl_847)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1374 = ~((~(or_dcpl_925 | or_dcpl_851)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1376 = ~((~(or_dcpl_925 | or_dcpl_854)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1378 = ~((~(or_dcpl_925 | or_dcpl_856)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1380 = ~((~(or_dcpl_925 | or_dcpl_859)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1382 = ~((~(or_dcpl_925 | or_dcpl_861)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1384 = ~((~(or_dcpl_925 | or_dcpl_864)) | act_config_is_zero_first_sva_dfm_4);
  assign and_dcpl_1386 = ~((~(or_dcpl_925 | or_dcpl_866)) | act_config_is_zero_first_sva_dfm_4);
  assign not_tmp_620 = ~((fsm_output[2]) & or_tmp_484);
  assign and_dcpl_1388 = ~((ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3:2]!=2'b00));
  assign and_dcpl_1390 = and_dcpl_1235 & and_dcpl_1388 & nor_1553_cse;
  assign and_dcpl_1391 = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1:0]==2'b01);
  assign and_dcpl_1393 = and_dcpl_1235 & and_dcpl_1388 & and_dcpl_1391;
  assign and_dcpl_1395 = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1:0]==2'b10);
  assign and_dcpl_1396 = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3:2]==2'b10);
  assign and_dcpl_1402 = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3:2]==2'b11);
  assign not_tmp_640 = MUX_s_1_2_2(and_dcpl_1056, (~ or_tmp_490), fsm_output[3]);
  assign or_dcpl_934 = (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign or_dcpl_936 = or_2265_cse | or_dcpl_934;
  assign or_dcpl_945 = (nvhls_get_slc_2U_NVUINT8_return_3_sva[1]) | (~ (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]));
  assign or_dcpl_946 = or_2265_cse | or_dcpl_945;
  assign or_dcpl_955 = (z_out[4]) | (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[0]));
  assign or_dcpl_956 = or_dcpl_955 | or_dcpl_934;
  assign or_dcpl_965 = or_dcpl_955 | or_dcpl_945;
  assign or_dcpl_974 = (~ (nvhls_get_slc_2U_NVUINT8_return_3_sva[1])) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign or_dcpl_975 = or_2265_cse | or_dcpl_974;
  assign or_dcpl_984 = ~((nvhls_get_slc_2U_NVUINT8_return_3_sva[1]) & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]));
  assign or_dcpl_985 = or_2265_cse | or_dcpl_984;
  assign or_dcpl_994 = or_dcpl_955 | or_dcpl_974;
  assign or_dcpl_1003 = or_dcpl_955 | or_dcpl_984;
  assign rva_out_reg_data_39_32_sva_dfm_6_mx0c0 = MUX_s_1_2_2(or_tmp_485, (~ or_3395_cse),
      fsm_output[3]);
  assign mux_435_nl = MUX_s_1_2_2((~ and_2371_cse), (fsm_output[0]), fsm_output[2]);
  assign act_config_output_counter_sva_mx0c0 = ~(mux_435_nl | (fsm_output[3]));
  assign act_config_output_counter_sva_mx0c1 = and_dcpl_1077 & (fsm_output[3]) &
      ActUnit_CheckStart_start_reg_sva;
  assign act_config_output_counter_sva_mx0c2 = and_dcpl_1077 & (fsm_output[3]) &
      (~ ActUnit_CheckStart_start_reg_sva);
  assign act_config_inst_counter_sva_mx0c1 = and_dcpl_1104 & (~(is_start_sva & is_incr_lpi_1_dfm_1));
  assign ActUnit_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva_mx0c4
      = nor_215_cse & and_dcpl_1081;
  assign nor_451_nl = ~((fsm_output[2]) | (fsm_output[0]));
  assign mux_446_nl = MUX_s_1_2_2((fsm_output[0]), nor_451_nl, fsm_output[3]);
  assign ActUnit_PushOutput_if_for_i_4_0_sva_3_0_mx0c0 = mux_446_nl & (~ (fsm_output[1]));
  assign act_regs_data_and_2749_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_0_13_sva_8_30_26_enexo_1
      | reg_is_start_enexo_174 | reg_act_config_is_zero_first_sva_dfm_4_enexo_174
      | reg_ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_1_30_26_enexo
      | reg_w_load_lpi_1_dfm_1_enexo_174 | reg_act_regs_data_0_13_sva_dfm_2_30_26_enexo);
  assign act_regs_data_and_2750_enex5 = act_regs_data_and_ssc & (reg_is_start_enexo_175
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_175 | reg_ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_1_25_22_enexo
      | reg_act_regs_data_0_13_sva_dfm_2_25_22_enexo | reg_act_regs_data_0_13_sva_8_25_22_enexo_1
      | reg_w_load_lpi_1_dfm_1_enexo_175);
  assign act_regs_data_and_2751_enex5 = act_regs_data_and_ssc & (reg_act_config_is_zero_first_sva_dfm_4_enexo_176
      | reg_Silu_for_16_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo
      | reg_act_regs_data_0_13_sva_8_21_0_enexo_1 | reg_act_regs_data_0_13_sva_dfm_2_21_0_enexo
      | reg_w_load_lpi_1_dfm_1_enexo_176 | reg_is_start_enexo_176);
  assign act_regs_data_and_2752_enex5 = act_regs_data_and_ssc & (reg_w_load_lpi_1_dfm_1_enexo_177
      | reg_ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_1_30_26_enexo
      | reg_act_regs_data_0_12_sva_8_30_26_enexo_1 | reg_is_start_enexo_177 | reg_act_config_is_zero_first_sva_dfm_4_enexo_177
      | reg_act_regs_data_0_12_sva_dfm_2_30_26_enexo);
  assign act_regs_data_and_2753_enex5 = act_regs_data_and_ssc & (reg_w_load_lpi_1_dfm_1_enexo_178
      | reg_ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_1_25_22_enexo
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_178 | reg_act_regs_data_0_12_sva_8_25_22_enexo_1
      | reg_act_regs_data_0_12_sva_dfm_2_25_22_enexo | reg_is_start_enexo_178);
  assign act_regs_data_and_2754_enex5 = act_regs_data_and_ssc & (reg_w_load_lpi_1_dfm_1_enexo_179
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_179 | reg_Silu_for_15_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo
      | reg_act_regs_data_0_12_sva_dfm_2_21_0_enexo | reg_is_start_enexo_179 | reg_act_regs_data_0_12_sva_8_21_0_enexo_1);
  assign act_regs_data_and_2755_enex5 = act_regs_data_and_ssc & (reg_ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_1_30_26_enexo
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_180 | reg_act_regs_data_0_11_sva_dfm_2_30_26_enexo
      | reg_is_start_enexo_180 | reg_w_load_lpi_1_dfm_1_enexo_180 | reg_act_regs_data_0_11_sva_8_30_26_enexo_1);
  assign act_regs_data_and_2756_enex5 = act_regs_data_and_ssc & (reg_is_start_enexo_181
      | reg_act_regs_data_0_11_sva_dfm_2_25_22_enexo | reg_ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_1_25_22_enexo
      | reg_w_load_lpi_1_dfm_1_enexo_181 | reg_act_config_is_zero_first_sva_dfm_4_enexo_181
      | reg_act_regs_data_0_11_sva_8_25_22_enexo_1);
  assign act_regs_data_and_2757_enex5 = act_regs_data_and_ssc & (reg_w_load_lpi_1_dfm_1_enexo_182
      | reg_act_regs_data_0_11_sva_dfm_2_21_0_enexo | reg_act_regs_data_0_11_sva_8_21_0_enexo_1
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_182 | reg_is_start_enexo_182
      | reg_Silu_for_14_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo);
  assign act_regs_data_and_2758_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_0_10_sva_dfm_2_30_26_enexo
      | reg_ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_1_30_26_enexo
      | reg_is_start_enexo_183 | reg_act_regs_data_0_10_sva_8_30_26_enexo_1 | reg_act_config_is_zero_first_sva_dfm_4_enexo_183
      | reg_w_load_lpi_1_dfm_1_enexo_183);
  assign act_regs_data_and_2759_enex5 = act_regs_data_and_ssc & (reg_is_start_enexo_184
      | reg_w_load_lpi_1_dfm_1_enexo_184 | reg_act_regs_data_0_10_sva_dfm_2_25_22_enexo
      | reg_act_regs_data_0_10_sva_8_25_22_enexo_1 | reg_act_config_is_zero_first_sva_dfm_4_enexo_184
      | reg_ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_1_25_22_enexo);
  assign act_regs_data_and_2760_enex5 = act_regs_data_and_ssc & (reg_Silu_for_13_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo
      | reg_w_load_lpi_1_dfm_1_enexo_185 | reg_act_regs_data_0_10_sva_dfm_2_21_0_enexo
      | reg_act_regs_data_0_10_sva_8_21_0_enexo_1 | reg_act_config_is_zero_first_sva_dfm_4_enexo_185
      | reg_is_start_enexo_185);
  assign act_regs_data_and_2761_enex5 = act_regs_data_and_ssc & (reg_act_regs_data_0_1_sva_dfm_2_30_26_enexo
      | reg_is_start_enexo_186 | reg_rva_out_reg_data_71_64_sva_dfm_6_1_enexo | reg_act_regs_data_0_1_sva_8_30_26_enexo_1
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_186 | reg_w_load_lpi_1_dfm_1_enexo_186);
  assign act_regs_data_and_2762_enex5 = act_regs_data_and_ssc & (reg_act_config_is_zero_first_sva_dfm_4_enexo_187
      | reg_rva_out_reg_data_39_32_sva_dfm_6_1_enexo | reg_act_regs_data_0_1_sva_dfm_2_25_22_enexo
      | reg_w_load_lpi_1_dfm_1_enexo_187 | reg_act_regs_data_0_1_sva_8_25_22_enexo_1
      | reg_is_start_enexo_187);
  assign act_regs_data_and_2763_enex5 = act_regs_data_and_ssc & (reg_is_start_enexo_188
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_188 | reg_w_load_lpi_1_dfm_1_enexo_188
      | reg_Silu_for_12_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo
      | reg_act_regs_data_0_1_sva_8_21_0_enexo_1 | reg_act_regs_data_0_1_sva_dfm_2_21_0_enexo);
  assign act_regs_data_and_2764_enex5 = act_regs_data_and_ssc & (reg_ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_1_30_26_enexo
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_189 | reg_act_regs_data_0_0_sva_8_30_26_enexo_1
      | reg_act_regs_data_0_0_sva_dfm_2_30_26_enexo | reg_w_load_lpi_1_dfm_1_enexo_189
      | reg_is_start_enexo_189);
  assign act_regs_data_and_2765_enex5 = act_regs_data_and_ssc & (reg_is_start_enexo_190
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_190 | reg_rva_out_reg_data_29_24_sva_dfm_6_1_enexo
      | reg_act_regs_data_0_0_sva_8_25_22_enexo_1 | reg_act_regs_data_0_0_sva_dfm_2_25_22_enexo
      | reg_w_load_lpi_1_dfm_1_enexo_190);
  assign act_regs_data_and_2766_enex5 = act_regs_data_and_ssc & (reg_Silu_for_11_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo
      | reg_act_regs_data_0_0_sva_dfm_2_21_0_enexo | reg_act_regs_data_0_0_sva_8_21_0_enexo_1
      | reg_act_config_is_zero_first_sva_dfm_4_enexo_191 | reg_w_load_lpi_1_dfm_1_enexo_191
      | reg_is_start_enexo_191);
  assign ActUnit_RunInst_switch_lp_and_816_enex5 = operator_32_8_true_AC_TRN_AC_WRAP_2_and_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_177 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_177
      | reg_act_regs_data_2_0_2_enexo_5 | reg_act_regs_data_3_0_2_enexo_5 | reg_act_config_inst_counter_enexo_177
      | reg_act_regs_data_1_0_2_enexo_5 | reg_act_regs_data_0_0_2_enexo_5);
  assign ActUnit_RunInst_switch_lp_and_817_enex5 = operator_32_8_true_AC_TRN_AC_WRAP_2_and_cse
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_178 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_178
      | reg_act_regs_data_2_0_3_enexo_5 | reg_act_regs_data_0_0_3_enexo_5 | reg_act_regs_data_1_0_3_enexo_5
      | reg_act_regs_data_3_0_3_enexo_5 | reg_act_config_inst_counter_enexo_178);
  assign ActUnit_RunInst_switch_lp_and_818_enex5 = operator_32_8_true_AC_TRN_AC_WRAP_2_and_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_179 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_179
      | reg_act_regs_data_3_0_1_enexo_5 | reg_act_regs_data_2_0_1_enexo_5 | reg_act_regs_data_0_0_1_enexo_5
      | reg_act_regs_data_1_0_1_enexo_5 | reg_act_config_inst_counter_enexo_179);
  assign nv_scvector_cctor_nv_scvector_5_for_and_enex5 = operator_32_8_true_AC_TRN_AC_WRAP_2_and_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_180 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_180
      | reg_act_config_inst_counter_enexo_180 | reg_act_regs_data_3_1_2_enexo_5 |
      reg_act_regs_data_1_1_2_enexo_5 | reg_act_regs_data_2_1_2_enexo_5 | reg_act_regs_data_0_1_2_enexo_5);
  assign nv_scvector_cctor_nv_scvector_5_for_and_15_enex5 = operator_32_8_true_AC_TRN_AC_WRAP_2_and_cse
      & (reg_act_regs_data_3_1_3_enexo_5 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_181
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_181 | reg_act_config_inst_counter_enexo_181
      | reg_act_regs_data_0_1_3_enexo_5 | reg_act_regs_data_2_1_3_enexo_5 | reg_act_regs_data_1_1_3_enexo_5);
  assign nv_scvector_cctor_nv_scvector_5_for_and_16_enex5 = operator_32_8_true_AC_TRN_AC_WRAP_2_and_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_182 | reg_act_regs_data_3_1_1_enexo_5
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_182 | reg_act_config_inst_counter_enexo_182
      | reg_act_regs_data_1_1_1_enexo_5 | reg_act_regs_data_0_1_1_enexo_5 | reg_act_regs_data_2_1_1_enexo_5);
  assign nv_scvector_cctor_nv_scvector_5_for_and_17_enex5 = operator_32_8_true_AC_TRN_AC_WRAP_2_and_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_183 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_183
      | reg_act_config_inst_counter_enexo_183 | reg_act_regs_data_0_2_2_enexo_5 |
      reg_act_regs_data_2_2_2_enexo_5 | reg_act_regs_data_3_2_2_enexo_5 | reg_act_regs_data_1_2_2_enexo_5);
  assign nv_scvector_cctor_nv_scvector_5_for_and_18_enex5 = operator_32_8_true_AC_TRN_AC_WRAP_2_and_cse
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_184 | reg_act_regs_data_1_2_3_enexo_5
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_184 | reg_act_regs_data_3_2_3_enexo_5
      | reg_act_regs_data_2_2_3_enexo_5 | reg_act_config_inst_counter_enexo_184 |
      reg_act_regs_data_0_2_3_enexo_5);
  assign nv_scvector_cctor_nv_scvector_5_for_and_19_enex5 = operator_32_8_true_AC_TRN_AC_WRAP_2_and_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_185 | reg_act_regs_data_1_2_1_enexo_5
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_185 | reg_act_regs_data_2_2_1_enexo_5
      | reg_act_regs_data_3_2_1_enexo_5 | reg_act_config_inst_counter_enexo_185 |
      reg_act_regs_data_0_2_1_enexo_5);
  assign nv_scvector_cctor_nv_scvector_5_for_and_20_enex5 = operator_32_8_true_AC_TRN_AC_WRAP_2_and_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_186 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_186
      | reg_act_regs_data_2_3_2_enexo_5 | reg_act_regs_data_3_3_2_enexo_5 | reg_act_regs_data_1_3_2_enexo_5
      | reg_act_config_inst_counter_enexo_186 | reg_act_regs_data_0_3_2_enexo_5);
  assign nv_scvector_cctor_nv_scvector_5_for_and_21_enex5 = operator_32_8_true_AC_TRN_AC_WRAP_2_and_cse
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_187 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_187
      | reg_act_regs_data_3_3_3_enexo_5 | reg_act_regs_data_1_3_3_enexo_5 | reg_act_config_inst_counter_enexo_187
      | reg_act_regs_data_2_3_3_enexo_5 | reg_act_regs_data_0_3_3_enexo_5);
  assign nv_scvector_cctor_nv_scvector_5_for_and_22_enex5 = operator_32_8_true_AC_TRN_AC_WRAP_2_and_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_188 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_188
      | reg_act_regs_data_3_3_1_enexo_5 | reg_act_regs_data_1_3_1_enexo_5 | reg_act_regs_data_2_3_1_enexo_5
      | reg_act_config_inst_counter_enexo_188 | reg_act_regs_data_0_3_1_enexo_5);
  assign nv_scvector_cctor_nv_scvector_5_for_and_23_enex5 = operator_32_8_true_AC_TRN_AC_WRAP_2_and_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_189 | reg_act_regs_data_0_4_2_enexo_5
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_189 | reg_act_config_inst_counter_enexo_189
      | reg_act_regs_data_1_4_2_enexo_5 | reg_act_regs_data_2_4_2_enexo_5 | reg_act_regs_data_3_4_2_enexo_5);
  assign nv_scvector_cctor_nv_scvector_5_for_and_24_enex5 = operator_32_8_true_AC_TRN_AC_WRAP_2_and_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_190 | reg_act_regs_data_0_4_3_enexo_5
      | reg_act_regs_data_2_4_3_enexo_5 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_190
      | reg_act_regs_data_3_4_3_enexo_5 | reg_act_regs_data_1_4_3_enexo_5 | reg_act_config_inst_counter_enexo_190);
  assign nv_scvector_cctor_nv_scvector_5_for_and_25_enex5 = operator_32_8_true_AC_TRN_AC_WRAP_2_and_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_191 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_191
      | reg_act_config_inst_counter_enexo_191 | reg_act_regs_data_2_4_1_enexo_5 |
      reg_act_regs_data_1_4_1_enexo_5 | reg_act_regs_data_0_4_1_enexo_5 | reg_act_regs_data_3_4_1_enexo_5);
  assign nv_scvector_cctor_nv_scvector_5_for_and_26_enex5 = operator_32_8_true_AC_TRN_AC_WRAP_2_and_cse
      & (reg_act_regs_data_0_5_2_enexo_5 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_192
      | reg_act_regs_data_3_5_2_enexo_5 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_192
      | reg_act_regs_data_1_5_2_enexo_5 | reg_act_config_inst_counter_enexo_192 |
      reg_act_regs_data_2_5_2_enexo_5);
  assign nv_scvector_cctor_nv_scvector_5_for_and_27_enex5 = operator_32_8_true_AC_TRN_AC_WRAP_2_and_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_193 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_193
      | reg_act_regs_data_1_5_3_enexo_5 | reg_act_regs_data_2_5_3_enexo_5 | reg_act_config_inst_counter_enexo_193
      | reg_act_regs_data_0_5_3_enexo_5 | reg_act_regs_data_3_5_3_enexo_5);
  assign nv_scvector_cctor_nv_scvector_5_for_and_28_enex5 = operator_32_8_true_AC_TRN_AC_WRAP_2_and_cse
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_194 | reg_act_config_inst_counter_enexo_194
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_194 | reg_act_regs_data_3_5_1_enexo_5
      | reg_act_regs_data_2_5_1_enexo_5 | reg_act_regs_data_0_5_1_enexo_5 | reg_act_regs_data_1_5_1_enexo_5);
  assign nv_scvector_cctor_nv_scvector_5_for_and_29_enex5 = operator_32_8_true_AC_TRN_AC_WRAP_2_and_cse
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_195 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_195
      | reg_act_regs_data_2_6_2_enexo_5 | reg_act_regs_data_3_6_2_enexo_5 | reg_act_regs_data_0_6_2_enexo_5
      | reg_act_regs_data_1_6_2_enexo_5 | reg_act_config_inst_counter_enexo_195);
  assign nv_scvector_cctor_nv_scvector_5_for_and_30_enex5 = operator_32_8_true_AC_TRN_AC_WRAP_2_and_cse
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_196 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_196
      | reg_act_regs_data_3_6_3_enexo_5 | reg_act_regs_data_0_6_3_enexo_5 | reg_act_regs_data_1_6_3_enexo_5
      | reg_act_regs_data_2_6_3_enexo_5 | reg_act_config_inst_counter_enexo_196);
  assign nv_scvector_cctor_nv_scvector_5_for_and_31_enex5 = operator_32_8_true_AC_TRN_AC_WRAP_2_and_cse
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_197 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_197
      | reg_act_config_inst_counter_enexo_197 | reg_act_regs_data_3_6_1_enexo_5 |
      reg_act_regs_data_2_6_1_enexo_5 | reg_act_regs_data_0_6_1_enexo_5 | reg_act_regs_data_1_6_1_enexo_5);
  assign nv_scvector_cctor_nv_scvector_5_for_and_32_enex5 = operator_32_8_true_AC_TRN_AC_WRAP_2_and_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_198 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_198
      | reg_act_regs_data_1_7_2_enexo_5 | reg_act_regs_data_3_7_2_enexo_5 | reg_act_regs_data_2_7_2_enexo_5
      | reg_act_regs_data_0_7_2_enexo_5 | reg_act_config_inst_counter_enexo_198);
  assign nv_scvector_cctor_nv_scvector_5_for_and_33_enex5 = operator_32_8_true_AC_TRN_AC_WRAP_2_and_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_199 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_199
      | reg_act_regs_data_3_7_3_enexo_5 | reg_act_config_inst_counter_enexo_199 |
      reg_act_regs_data_1_7_3_enexo_5 | reg_act_regs_data_2_7_3_enexo_5 | reg_act_regs_data_0_7_3_enexo_5);
  assign nv_scvector_cctor_nv_scvector_5_for_and_34_enex5 = operator_32_8_true_AC_TRN_AC_WRAP_2_and_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_200 | reg_act_regs_data_0_7_1_enexo_5
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_200 | reg_act_regs_data_3_7_1_enexo_5
      | reg_act_config_inst_counter_enexo_200 | reg_act_regs_data_1_7_1_enexo_5 |
      reg_act_regs_data_2_7_1_enexo_5);
  assign nv_scvector_cctor_nv_scvector_5_for_and_35_enex5 = ActUnit_RunInst_switch_lp_and_802_cse
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_201 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_201
      | reg_act_regs_data_2_8_2_enexo_5 | reg_act_regs_data_3_8_2_enexo_5 | reg_act_config_inst_counter_enexo_201
      | reg_act_regs_data_1_8_2_enexo_5 | reg_act_regs_data_0_8_2_enexo_5);
  assign nv_scvector_cctor_nv_scvector_5_for_and_36_enex5 = ActUnit_RunInst_switch_lp_and_802_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_202 | reg_act_regs_data_0_8_3_enexo_5
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_202 | reg_act_regs_data_3_8_3_enexo_5
      | reg_act_regs_data_2_8_3_enexo_5 | reg_act_regs_data_1_8_3_enexo_5 | reg_act_config_inst_counter_enexo_202);
  assign nv_scvector_cctor_nv_scvector_5_for_and_37_enex5 = ActUnit_RunInst_switch_lp_and_802_cse
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_203 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_203
      | reg_act_config_inst_counter_enexo_203 | reg_act_regs_data_0_8_1_enexo_5 |
      reg_act_regs_data_3_8_1_enexo_5 | reg_act_regs_data_1_8_1_enexo_5 | reg_act_regs_data_2_8_1_enexo_5);
  assign nv_scvector_cctor_nv_scvector_5_for_and_38_enex5 = ActUnit_RunInst_switch_lp_and_802_cse
      & (reg_act_regs_data_0_9_2_enexo_5 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_204
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_204 | reg_act_config_inst_counter_enexo_204
      | reg_act_regs_data_1_9_2_enexo_5 | reg_act_regs_data_2_9_2_enexo_5 | reg_act_regs_data_3_9_2_enexo_5);
  assign nv_scvector_cctor_nv_scvector_5_for_and_39_enex5 = ActUnit_RunInst_switch_lp_and_802_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_205 | reg_act_regs_data_3_9_3_enexo_5
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_205 | reg_act_regs_data_1_9_3_enexo_5
      | reg_act_config_inst_counter_enexo_205 | reg_act_regs_data_2_9_3_enexo_5 |
      reg_act_regs_data_0_9_3_enexo_5);
  assign nv_scvector_cctor_nv_scvector_5_for_and_40_enex5 = ActUnit_RunInst_switch_lp_and_802_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_206 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_206
      | reg_act_regs_data_3_9_1_enexo_5 | reg_act_regs_data_1_9_1_enexo_5 | reg_act_config_inst_counter_enexo_206
      | reg_act_regs_data_2_9_1_enexo_5 | reg_act_regs_data_0_9_1_enexo_5);
  assign nv_scvector_cctor_nv_scvector_5_for_and_41_enex5 = ActUnit_RunInst_switch_lp_and_802_cse
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_207 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_207
      | reg_act_regs_data_1_10_2_enexo_5 | reg_act_regs_data_3_10_2_enexo_5 | reg_act_regs_data_2_10_2_enexo_5
      | reg_act_regs_data_0_10_2_enexo_5 | reg_act_config_inst_counter_enexo_207);
  assign nv_scvector_cctor_nv_scvector_5_for_and_42_enex5 = ActUnit_RunInst_switch_lp_and_802_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_208 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_208
      | reg_act_config_inst_counter_enexo_208 | reg_act_regs_data_2_10_3_enexo_5
      | reg_act_regs_data_3_10_3_enexo_5 | reg_act_regs_data_1_10_3_enexo_5 | reg_act_regs_data_0_10_3_enexo_5);
  assign nv_scvector_cctor_nv_scvector_5_for_and_43_enex5 = ActUnit_RunInst_switch_lp_and_802_cse
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_209 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_209
      | reg_act_regs_data_1_10_1_enexo_5 | reg_act_regs_data_0_10_1_enexo_5 | reg_act_regs_data_2_10_1_enexo_5
      | reg_act_regs_data_3_10_1_enexo_5 | reg_act_config_inst_counter_enexo_209);
  assign nv_scvector_cctor_nv_scvector_5_for_and_44_enex5 = ActUnit_RunInst_switch_lp_and_802_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_210 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_210
      | reg_act_regs_data_3_11_2_enexo_5 | reg_act_regs_data_2_11_2_enexo_5 | reg_act_config_inst_counter_enexo_210
      | reg_act_regs_data_0_11_2_enexo_5 | reg_act_regs_data_1_11_2_enexo_5);
  assign nv_scvector_cctor_nv_scvector_5_for_and_45_enex5 = ActUnit_RunInst_switch_lp_and_802_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_211 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_211
      | reg_act_config_inst_counter_enexo_211 | reg_act_regs_data_3_11_3_enexo_5
      | reg_act_regs_data_1_11_3_enexo_5 | reg_act_regs_data_2_11_3_enexo_5 | reg_act_regs_data_0_11_3_enexo_5);
  assign nv_scvector_cctor_nv_scvector_5_for_and_46_enex5 = ActUnit_RunInst_switch_lp_and_802_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_212 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_212
      | reg_act_config_inst_counter_enexo_212 | reg_act_regs_data_1_11_1_enexo_5
      | reg_act_regs_data_3_11_1_enexo_5 | reg_act_regs_data_2_11_1_enexo_5 | reg_act_regs_data_0_11_1_enexo_5);
  assign nv_scvector_cctor_nv_scvector_5_for_and_47_enex5 = ActUnit_RunInst_switch_lp_and_802_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_213 | reg_act_config_inst_counter_enexo_213
      | reg_act_config_inst_regs_20_sva_dfm_6_enexo_213 | reg_act_regs_data_2_12_2_enexo_5
      | reg_act_regs_data_1_12_2_enexo_5 | reg_act_regs_data_3_12_2_enexo_5 | reg_act_regs_data_0_12_2_enexo_5);
  assign nv_scvector_cctor_nv_scvector_5_for_and_48_enex5 = ActUnit_RunInst_switch_lp_and_802_cse
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_214 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_214
      | reg_act_regs_data_0_12_3_enexo_5 | reg_act_regs_data_3_12_3_enexo_5 | reg_act_regs_data_2_12_3_enexo_5
      | reg_act_config_inst_counter_enexo_214 | reg_act_regs_data_1_12_3_enexo_5);
  assign nv_scvector_cctor_nv_scvector_5_for_and_49_enex5 = ActUnit_RunInst_switch_lp_and_802_cse
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_215 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_215
      | reg_act_regs_data_0_12_1_enexo_5 | reg_act_config_inst_counter_enexo_215
      | reg_act_regs_data_3_12_1_enexo_5 | reg_act_regs_data_2_12_1_enexo_5 | reg_act_regs_data_1_12_1_enexo_5);
  assign nv_scvector_cctor_nv_scvector_5_for_and_50_enex5 = ActUnit_RunInst_switch_lp_and_802_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_216 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_216
      | reg_act_regs_data_2_13_2_enexo_5 | reg_act_regs_data_3_13_2_enexo_5 | reg_act_regs_data_1_13_2_enexo_5
      | reg_act_regs_data_0_13_2_enexo_5 | reg_act_config_inst_counter_enexo_216);
  assign nv_scvector_cctor_nv_scvector_5_for_and_51_enex5 = ActUnit_RunInst_switch_lp_and_802_cse
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_217 | reg_act_regs_data_1_13_3_enexo_5
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_217 | reg_act_regs_data_3_13_3_enexo_5
      | reg_act_config_inst_counter_enexo_217 | reg_act_regs_data_2_13_3_enexo_5
      | reg_act_regs_data_0_13_3_enexo_5);
  assign nv_scvector_cctor_nv_scvector_5_for_and_52_enex5 = ActUnit_RunInst_switch_lp_and_802_cse
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_218 | reg_act_config_inst_counter_enexo_218
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_218 | reg_act_regs_data_0_13_1_enexo_5
      | reg_act_regs_data_3_13_1_enexo_5 | reg_act_regs_data_2_13_1_enexo_5 | reg_act_regs_data_1_13_1_enexo_5);
  assign nv_scvector_cctor_nv_scvector_5_for_and_53_enex5 = ActUnit_RunInst_switch_lp_and_802_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_219 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_219
      | reg_act_config_inst_counter_enexo_219 | reg_act_regs_data_0_14_2_enexo_5
      | reg_act_regs_data_1_14_2_enexo_5 | reg_act_regs_data_2_14_2_enexo_5 | reg_act_regs_data_3_14_2_enexo_5);
  assign nv_scvector_cctor_nv_scvector_5_for_and_54_enex5 = ActUnit_RunInst_switch_lp_and_802_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_220 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_220
      | reg_act_regs_data_3_14_3_enexo_5 | reg_act_regs_data_0_14_3_enexo_5 | reg_act_regs_data_2_14_3_enexo_5
      | reg_act_regs_data_1_14_3_enexo_5 | reg_act_config_inst_counter_enexo_220);
  assign nv_scvector_cctor_nv_scvector_5_for_and_55_enex5 = ActUnit_RunInst_switch_lp_and_802_cse
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_221 | reg_act_regs_data_0_14_1_enexo_5
      | reg_act_config_inst_regs_4_sva_dfm_5_enexo_221 | reg_act_regs_data_1_14_1_enexo_5
      | reg_act_regs_data_3_14_1_enexo_5 | reg_act_regs_data_2_14_1_enexo_5 | reg_act_config_inst_counter_enexo_221);
  assign nv_scvector_cctor_nv_scvector_5_for_and_56_enex5 = ActUnit_RunInst_switch_lp_and_802_cse
      & (reg_act_config_inst_regs_4_sva_dfm_5_enexo_222 | reg_act_config_inst_regs_20_sva_dfm_6_enexo_222
      | reg_act_config_inst_counter_enexo_222 | reg_act_regs_data_3_15_2_enexo_5
      | reg_act_regs_data_1_15_2_enexo_5 | reg_act_regs_data_0_15_2_enexo_5 | reg_act_regs_data_2_15_2_enexo_5);
  assign nv_scvector_cctor_nv_scvector_5_for_and_57_enex5 = ActUnit_RunInst_switch_lp_and_802_cse
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_223 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_223
      | reg_act_config_inst_counter_enexo_223 | reg_act_regs_data_2_15_3_enexo_5
      | reg_act_regs_data_3_15_3_enexo_5 | reg_act_regs_data_1_15_3_enexo_5 | reg_act_regs_data_0_15_3_enexo_5);
  assign nv_scvector_cctor_nv_scvector_5_for_and_58_enex5 = ActUnit_RunInst_switch_lp_and_802_cse
      & (reg_act_config_inst_regs_20_sva_dfm_6_enexo_224 | reg_act_config_inst_regs_4_sva_dfm_5_enexo_224
      | reg_act_config_inst_counter_enexo_224 | reg_act_regs_data_1_15_1_enexo_5
      | reg_act_regs_data_3_15_1_enexo_5 | reg_act_regs_data_0_15_1_enexo_5 | reg_act_regs_data_2_15_1_enexo_5);
  assign nl_Silu_for_10_else_else_else_if_acc_nl = conv_u2u_25_26({reg_nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , (reg_nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:1])})
      + ({reg_nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1});
  assign Silu_for_10_else_else_else_if_acc_nl = nl_Silu_for_10_else_else_else_if_acc_nl[25:0];
  assign Silu_for_10_else_else_else_if_acc_itm_25_1_1 = readslicef_26_25_1(Silu_for_10_else_else_else_if_acc_nl);
  assign Silu_for_else_else_else_if_and_1_ssc = ActUnitRun_wen & ((act_config_in_InstFetch_return_sva_7_2[2])
      | and_dcpl_331 | and_dcpl_1235);
  assign nl_Silu_for_11_else_else_else_if_acc_nl = conv_u2u_25_26({reg_nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , (reg_nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:1])})
      + ({reg_nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1});
  assign Silu_for_11_else_else_else_if_acc_nl = nl_Silu_for_11_else_else_else_if_acc_nl[25:0];
  assign Silu_for_11_else_else_else_if_acc_itm_25_1_1 = readslicef_26_25_1(Silu_for_11_else_else_else_if_acc_nl);
  assign Silu_for_else_else_else_if_and_2_ssc = ActUnitRun_wen & ((act_config_in_InstFetch_return_sva_7_2[2])
      | and_dcpl_331 | (~ mux_tmp_433));
  assign Silu_for_else_else_else_if_or_13_rgt = and_dcpl_1112 | (~ mux_tmp_433);
  assign nl_Silu_for_12_else_else_else_if_acc_nl = conv_u2u_25_26({reg_nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , (reg_nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:1])})
      + ({reg_nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1});
  assign Silu_for_12_else_else_else_if_acc_nl = nl_Silu_for_12_else_else_else_if_acc_nl[25:0];
  assign Silu_for_12_else_else_else_if_acc_itm_25_1_1 = readslicef_26_25_1(Silu_for_12_else_else_else_if_acc_nl);
  assign Silu_for_else_else_else_if_and_3_ssc = ActUnitRun_wen & ((act_config_in_InstFetch_return_sva_7_2[2])
      | and_dcpl_331 | (~ mux_448_itm));
  assign Silu_for_else_else_else_if_or_14_cse = and_dcpl_1112 | (~ mux_448_itm);
  assign nor_1654_cse = ~(nor_320_cse | (fsm_output[3]));
  assign nl_Silu_for_13_else_else_else_if_acc_nl = conv_u2u_25_26({reg_nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , (reg_nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:1])})
      + ({reg_nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1});
  assign Silu_for_13_else_else_else_if_acc_nl = nl_Silu_for_13_else_else_else_if_acc_nl[25:0];
  assign Silu_for_13_else_else_else_if_acc_itm_25_1_1 = readslicef_26_25_1(Silu_for_13_else_else_else_if_acc_nl);
  assign nl_Silu_for_14_else_else_else_if_acc_nl = conv_u2u_25_26({reg_nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , (reg_nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:1])})
      + ({reg_nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1});
  assign Silu_for_14_else_else_else_if_acc_nl = nl_Silu_for_14_else_else_else_if_acc_nl[25:0];
  assign Silu_for_14_else_else_else_if_acc_itm_25_1_1 = readslicef_26_25_1(Silu_for_14_else_else_else_if_acc_nl);
  assign nl_Silu_for_15_else_else_else_if_acc_nl = conv_u2u_25_26({reg_nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , (reg_nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:1])})
      + ({reg_nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1});
  assign Silu_for_15_else_else_else_if_acc_nl = nl_Silu_for_15_else_else_else_if_acc_nl[25:0];
  assign Silu_for_15_else_else_else_if_acc_itm_25_1_1 = readslicef_26_25_1(Silu_for_15_else_else_else_if_acc_nl);
  assign nl_Silu_for_16_else_else_else_if_acc_nl = conv_u2u_25_26({reg_nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , (reg_nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:1])})
      + ({reg_nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
      , reg_nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1});
  assign Silu_for_16_else_else_else_if_acc_nl = nl_Silu_for_16_else_else_else_if_acc_nl[25:0];
  assign Silu_for_16_else_else_else_if_acc_itm_25_1_1 = readslicef_26_25_1(Silu_for_16_else_else_else_if_acc_nl);
  assign and_dcpl_1426 = and_dcpl_1236 & (~ nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_291);
  assign mux_459_nl = MUX_s_1_2_2(not_tmp_620, or_3395_cse, fsm_output[3]);
  assign or_dcpl_1012 = and_dcpl_1426 | mux_459_nl;
  assign or_dcpl_1013 = ~(and_dcpl_1257 | act_config_ActConfigRead_else_else_not_21);
  assign or_dcpl_1014 = and_dcpl_1262 | ActUnit_DecodeAxiRead_unequal_tmp_1;
  assign or_dcpl_1015 = and_dcpl_1426 | mux_tmp_433;
  assign nor_471_nl = ~((fsm_output[1:0]!=2'b10));
  assign nor_472_nl = ~((fsm_output[2:0]!=3'b001));
  assign not_tmp_646 = MUX_s_1_2_2(nor_471_nl, nor_472_nl, fsm_output[3]);
  assign Silu_for_else_if_and_1_cse = (~ (act_config_in_InstFetch_mux_tmp[4])) &
      and_dcpl_847;
  assign Silu_for_else_if_and_2_cse = (act_config_in_InstFetch_mux_tmp[4]) & and_dcpl_847;
  assign or_tmp_552 = (fsm_output[3:2]!=2'b01);
  assign or_tmp_555 = (fsm_output[0]) | (fsm_output[3]) | (~ (fsm_output[2]));
  assign or_tmp_653 = (~ (fsm_output[0])) | (fsm_output[3]) | (fsm_output[2]);
  assign or_tmp_871 = ActUnit_RunInst_switch_lp_equal_tmp_8 | ActUnit_RunInst_switch_lp_equal_tmp_7
      | ActUnit_RunInst_switch_lp_equal_tmp_6 | ActUnit_RunInst_switch_lp_equal_tmp_5
      | ActUnit_RunInst_switch_lp_equal_tmp_4;
  assign and_2824_cse = ActUnit_RunInst_switch_lp_equal_tmp_2 & ActUnit_RunInst_switch_lp_and_tmp;
  assign and_2825_cse = or_tmp_871 & reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_nor_cse;
  assign or_tmp_873 = and_2824_cse | and_2825_cse | while_nand_64_ssc_1;
  assign or_tmp_938 = (fsm_output[3:1]!=3'b010) | nand_543_cse;
  assign or_tmp_999 = ActUnit_RunInst_switch_lp_equal_tmp_7 | ActUnit_RunInst_switch_lp_equal_tmp_6
      | ActUnit_RunInst_switch_lp_equal_tmp_5 | ActUnit_RunInst_switch_lp_equal_tmp_4;
  assign and_2872_cse = ActUnit_RunInst_switch_lp_equal_tmp_2 & ActUnit_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva;
  assign nand_tmp_41 = ~(while_nor_16_itm & (~(and_2872_cse | (~((~(or_tmp_999 &
      reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_1_cse)) & is_start_sva
      & (~(ActUnit_RunInst_switch_lp_equal_tmp_8 & ActUnit_PushOutput_if_for_and_stg_2_7_sva)))))));
  assign or_tmp_1057 = (fsm_output[3:1]!=3'b010) | nand_583_cse;
  assign and_2936_cse = ActUnit_RunInst_switch_lp_equal_tmp_2 & ActUnit_RunInst_switch_lp_and_32_tmp;
  assign and_2937_cse = or_tmp_871 & reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_cse;
  assign or_tmp_1113 = and_2936_cse | and_2937_cse | while_nand_96_ssc_1;
  assign or_tmp_1178 = (fsm_output[3:1]!=3'b010) | nand_623_cse;
  assign and_2984_cse = ActUnit_RunInst_switch_lp_equal_tmp_2 & ActUnit_CheckStart_start_reg_sva;
  assign nand_tmp_73 = ~(while_nor_48_itm & (~(and_2984_cse | (~((~(or_tmp_999 &
      reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_2_cse)) & is_start_sva
      & (~(ActUnit_RunInst_switch_lp_equal_tmp_8 & Gelu_for_and_2_cse_sva)))))));
  assign or_tmp_1297 = (fsm_output[3:1]!=3'b010) | nand_663_cse;
  assign nand_tmp_104 = ~(while_nor_itm & is_start_sva & (~(and_2824_cse | and_2825_cse)));
  assign or_tmp_1408 = (fsm_output[3:1]!=3'b010) | nand_704_cse;
  assign nor_tmp_635 = ActUnit_RunInst_switch_lp_equal_tmp_8 & ActUnit_PushOutput_if_for_and_stg_2_7_sva;
  assign or_2499_nl = or_tmp_999 | nor_tmp_635;
  assign mux_1050_nl = MUX_s_1_2_2(nor_tmp_635, or_2499_nl, reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_1_cse);
  assign nand_tmp_120 = ~(while_nor_16_itm & is_start_sva & (~(and_2872_cse | mux_1050_nl)));
  assign or_tmp_1529 = (fsm_output[3:1]!=3'b010) | nand_744_cse;
  assign nand_tmp_136 = ~(while_nor_32_itm & is_start_sva & (~(and_2936_cse | and_2937_cse)));
  assign or_tmp_1648 = (fsm_output[3:1]!=3'b010) | nand_784_cse;
  assign nor_tmp_771 = ActUnit_RunInst_switch_lp_equal_tmp_8 & Gelu_for_and_2_cse_sva;
  assign or_2739_nl = or_tmp_999 | nor_tmp_771;
  assign mux_1178_nl = MUX_s_1_2_2(nor_tmp_771, or_2739_nl, reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_2_cse);
  assign nand_tmp_152 = ~(while_nor_48_itm & is_start_sva & (~(and_2984_cse | mux_1178_nl)));
  assign or_tmp_1769 = (fsm_output[3:1]!=3'b010) | nand_824_cse;
  assign not_tmp_2198 = ~((ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]) & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[0])
      & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[1]));
  assign or_dcpl = and_dcpl_1426 | and_dcpl_1244;
  assign is_start_and_tmp = ActUnitRun_wen & (and_dcpl_1083 | and_dcpl_1085);
  assign mux_1248_nl = MUX_s_1_2_2(or_tmp_1769, (~ mux_1180_cse), and_2533_cse);
  assign mux_1249_nl = MUX_s_1_2_2(mux_1248_nl, or_tmp_1769, z_out[4]);
  assign and_2189_tmp = (~ mux_1249_nl) & ActUnitRun_wen;
  assign w_load_and_tmp = ActUnitRun_wen & ((is_start_sva & (~ or_dcpl_822)) | and_dcpl_847)
      & or_243_cse;
  assign mux_1243_nl = MUX_s_1_2_2(or_tmp_1769, (~ mux_1180_cse), and_2494_cse);
  assign mux_1244_nl = MUX_s_1_2_2(mux_1243_nl, or_tmp_1769, or_2371_cse);
  assign and_2187_tmp = (~ mux_1244_nl) & ActUnitRun_wen;
  assign mux_1238_nl = MUX_s_1_2_2(or_tmp_1769, (~ mux_1180_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_1239_nl = MUX_s_1_2_2(mux_1238_nl, or_tmp_1769, or_2364_cse);
  assign and_2185_tmp = (~ mux_1239_nl) & ActUnitRun_wen;
  assign mux_1233_nl = MUX_s_1_2_2(or_tmp_1769, (~ mux_1180_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_1234_nl = MUX_s_1_2_2(mux_1233_nl, or_tmp_1769, or_2357_cse);
  assign and_2183_tmp = (~ mux_1234_nl) & ActUnitRun_wen;
  assign mux_1228_nl = MUX_s_1_2_2(or_tmp_1769, (~ mux_1180_cse), and_2484_cse);
  assign mux_1229_nl = MUX_s_1_2_2(mux_1228_nl, or_tmp_1769, or_2350_cse);
  assign and_2181_tmp = (~ mux_1229_nl) & ActUnitRun_wen;
  assign mux_1223_nl = MUX_s_1_2_2(or_tmp_1769, (~ mux_1180_cse), and_2484_cse);
  assign mux_1224_nl = MUX_s_1_2_2(mux_1223_nl, or_tmp_1769, or_2343_cse);
  assign and_2179_tmp = (~ mux_1224_nl) & ActUnitRun_wen;
  assign mux_1218_nl = MUX_s_1_2_2(or_tmp_1769, (~ mux_1180_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_1219_nl = MUX_s_1_2_2(mux_1218_nl, or_tmp_1769, or_2336_cse);
  assign and_2177_tmp = (~ mux_1219_nl) & ActUnitRun_wen;
  assign mux_1213_nl = MUX_s_1_2_2(or_tmp_1769, (~ mux_1180_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_1214_nl = MUX_s_1_2_2(mux_1213_nl, or_tmp_1769, or_2329_cse);
  assign and_2175_tmp = (~ mux_1214_nl) & ActUnitRun_wen;
  assign mux_1209_nl = MUX_s_1_2_2(mux_1180_cse, nor_1610_cse, nand_685_cse);
  assign and_2173_tmp = mux_1209_nl & ActUnitRun_wen;
  assign mux_1205_nl = MUX_s_1_2_2(mux_1180_cse, nor_1610_cse, or_2315_cse);
  assign and_2171_tmp = mux_1205_nl & ActUnitRun_wen;
  assign mux_1201_nl = MUX_s_1_2_2(mux_1180_cse, nor_1610_cse, or_2308_cse);
  assign and_2169_tmp = mux_1201_nl & ActUnitRun_wen;
  assign mux_1197_nl = MUX_s_1_2_2(mux_1180_cse, nor_1610_cse, or_2301_cse);
  assign and_2167_tmp = mux_1197_nl & ActUnitRun_wen;
  assign mux_1193_nl = MUX_s_1_2_2(mux_1180_cse, nor_1610_cse, or_2294_cse);
  assign and_2165_tmp = mux_1193_nl & ActUnitRun_wen;
  assign mux_1189_nl = MUX_s_1_2_2(mux_1180_cse, nor_1610_cse, or_2287_cse);
  assign and_2163_tmp = mux_1189_nl & ActUnitRun_wen;
  assign mux_1185_nl = MUX_s_1_2_2(mux_1180_cse, nor_1610_cse, or_2280_cse);
  assign and_2161_tmp = mux_1185_nl & ActUnitRun_wen;
  assign mux_1181_nl = MUX_s_1_2_2(mux_1180_cse, nor_1610_cse, or_2273_cse);
  assign and_2159_tmp = mux_1181_nl & ActUnitRun_wen;
  assign mux_1176_nl = MUX_s_1_2_2(or_tmp_1648, (~ mux_1123_cse), and_2497_cse);
  assign mux_1177_nl = MUX_s_1_2_2(mux_1176_nl, or_tmp_1648, or_2265_cse);
  assign and_2157_tmp = (~ mux_1177_nl) & ActUnitRun_wen;
  assign mux_1172_nl = MUX_s_1_2_2(or_tmp_1648, (~ mux_1123_cse), and_2494_cse);
  assign mux_1173_nl = MUX_s_1_2_2(mux_1172_nl, or_tmp_1648, or_2257_cse);
  assign and_2155_tmp = (~ mux_1173_nl) & ActUnitRun_wen;
  assign mux_1168_nl = MUX_s_1_2_2(or_tmp_1648, (~ mux_1123_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_1169_nl = MUX_s_1_2_2(mux_1168_nl, or_tmp_1648, or_2249_cse);
  assign and_2153_tmp = (~ mux_1169_nl) & ActUnitRun_wen;
  assign mux_1164_nl = MUX_s_1_2_2(or_tmp_1648, (~ mux_1123_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_1165_nl = MUX_s_1_2_2(mux_1164_nl, or_tmp_1648, or_2241_cse);
  assign and_2151_tmp = (~ mux_1165_nl) & ActUnitRun_wen;
  assign mux_1160_nl = MUX_s_1_2_2(or_tmp_1648, (~ mux_1123_cse), and_2484_cse);
  assign mux_1161_nl = MUX_s_1_2_2(mux_1160_nl, or_tmp_1648, or_2233_cse);
  assign and_2149_tmp = (~ mux_1161_nl) & ActUnitRun_wen;
  assign mux_1156_nl = MUX_s_1_2_2(or_tmp_1648, (~ mux_1123_cse), and_2484_cse);
  assign mux_1157_nl = MUX_s_1_2_2(mux_1156_nl, or_tmp_1648, or_2225_cse);
  assign and_2147_tmp = (~ mux_1157_nl) & ActUnitRun_wen;
  assign mux_1152_nl = MUX_s_1_2_2(or_tmp_1648, (~ mux_1123_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_1153_nl = MUX_s_1_2_2(mux_1152_nl, or_tmp_1648, or_2217_cse);
  assign and_2145_tmp = (~ mux_1153_nl) & ActUnitRun_wen;
  assign mux_1148_nl = MUX_s_1_2_2(or_tmp_1648, (~ mux_1123_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_1149_nl = MUX_s_1_2_2(mux_1148_nl, or_tmp_1648, or_2209_cse);
  assign and_2143_tmp = (~ mux_1149_nl) & ActUnitRun_wen;
  assign mux_1145_nl = MUX_s_1_2_2(mux_1123_cse, nor_1602_cse, or_2201_cse);
  assign and_2141_tmp = mux_1145_nl & ActUnitRun_wen;
  assign mux_1142_nl = MUX_s_1_2_2(mux_1123_cse, nor_1602_cse, or_2193_cse);
  assign and_2139_tmp = mux_1142_nl & ActUnitRun_wen;
  assign mux_1139_nl = MUX_s_1_2_2(mux_1123_cse, nor_1602_cse, or_2185_cse);
  assign and_2137_tmp = mux_1139_nl & ActUnitRun_wen;
  assign mux_1136_nl = MUX_s_1_2_2(mux_1123_cse, nor_1602_cse, or_2177_cse);
  assign and_2135_tmp = mux_1136_nl & ActUnitRun_wen;
  assign mux_1133_nl = MUX_s_1_2_2(mux_1123_cse, nor_1602_cse, or_2169_cse);
  assign and_2133_tmp = mux_1133_nl & ActUnitRun_wen;
  assign mux_1130_nl = MUX_s_1_2_2(mux_1123_cse, nor_1602_cse, or_2161_cse);
  assign and_2131_tmp = mux_1130_nl & ActUnitRun_wen;
  assign mux_1127_nl = MUX_s_1_2_2(mux_1123_cse, nor_1602_cse, or_2153_cse);
  assign and_2129_tmp = mux_1127_nl & ActUnitRun_wen;
  assign mux_1124_nl = MUX_s_1_2_2(mux_1123_cse, nor_1602_cse, or_2145_cse);
  assign and_2127_tmp = mux_1124_nl & ActUnitRun_wen;
  assign mux_1120_nl = MUX_s_1_2_2(or_tmp_1529, (~ mux_1052_cse), and_2412_cse);
  assign mux_1121_nl = MUX_s_1_2_2(mux_1120_nl, or_tmp_1529, or_2138_cse);
  assign and_2125_tmp = (~ mux_1121_nl) & ActUnitRun_wen;
  assign mux_1115_nl = MUX_s_1_2_2(or_tmp_1529, (~ mux_1052_cse), and_2412_cse);
  assign mux_1116_nl = MUX_s_1_2_2(mux_1115_nl, or_tmp_1529, or_2131_cse);
  assign and_2123_tmp = (~ mux_1116_nl) & ActUnitRun_wen;
  assign mux_1110_nl = MUX_s_1_2_2(or_tmp_1529, (~ mux_1052_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_1111_nl = MUX_s_1_2_2(mux_1110_nl, or_tmp_1529, or_2124_cse);
  assign and_2121_tmp = (~ mux_1111_nl) & ActUnitRun_wen;
  assign mux_1105_nl = MUX_s_1_2_2(or_tmp_1529, (~ mux_1052_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_1106_nl = MUX_s_1_2_2(mux_1105_nl, or_tmp_1529, or_2117_cse);
  assign and_2119_tmp = (~ mux_1106_nl) & ActUnitRun_wen;
  assign mux_1100_nl = MUX_s_1_2_2(or_tmp_1529, (~ mux_1052_cse), and_2412_cse);
  assign mux_1101_nl = MUX_s_1_2_2(mux_1100_nl, or_tmp_1529, or_2110_cse);
  assign and_2117_tmp = (~ mux_1101_nl) & ActUnitRun_wen;
  assign mux_1095_nl = MUX_s_1_2_2(or_tmp_1529, (~ mux_1052_cse), and_2412_cse);
  assign mux_1096_nl = MUX_s_1_2_2(mux_1095_nl, or_tmp_1529, or_2103_cse);
  assign and_2115_tmp = (~ mux_1096_nl) & ActUnitRun_wen;
  assign mux_1090_nl = MUX_s_1_2_2(or_tmp_1529, (~ mux_1052_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_1091_nl = MUX_s_1_2_2(mux_1090_nl, or_tmp_1529, or_2096_cse);
  assign and_2113_tmp = (~ mux_1091_nl) & ActUnitRun_wen;
  assign mux_1085_nl = MUX_s_1_2_2(or_tmp_1529, (~ mux_1052_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_1086_nl = MUX_s_1_2_2(mux_1085_nl, or_tmp_1529, or_2089_cse);
  assign and_2111_tmp = (~ mux_1086_nl) & ActUnitRun_wen;
  assign mux_1081_nl = MUX_s_1_2_2(mux_1052_cse, nor_1594_cse, or_2082_cse);
  assign and_2109_tmp = mux_1081_nl & ActUnitRun_wen;
  assign mux_1077_nl = MUX_s_1_2_2(mux_1052_cse, nor_1594_cse, or_2075_cse);
  assign and_2107_tmp = mux_1077_nl & ActUnitRun_wen;
  assign mux_1073_nl = MUX_s_1_2_2(mux_1052_cse, nor_1594_cse, or_2068_cse);
  assign and_2105_tmp = mux_1073_nl & ActUnitRun_wen;
  assign mux_1069_nl = MUX_s_1_2_2(mux_1052_cse, nor_1594_cse, or_2061_cse);
  assign and_2103_tmp = mux_1069_nl & ActUnitRun_wen;
  assign mux_1065_nl = MUX_s_1_2_2(mux_1052_cse, nor_1594_cse, or_2054_cse);
  assign and_2101_tmp = mux_1065_nl & ActUnitRun_wen;
  assign mux_1061_nl = MUX_s_1_2_2(mux_1052_cse, nor_1594_cse, or_2047_cse);
  assign and_2099_tmp = mux_1061_nl & ActUnitRun_wen;
  assign mux_1057_nl = MUX_s_1_2_2(mux_1052_cse, nor_1594_cse, or_2040_cse);
  assign and_2097_tmp = mux_1057_nl & ActUnitRun_wen;
  assign mux_1053_nl = MUX_s_1_2_2(mux_1052_cse, nor_1594_cse, or_2033_cse);
  assign and_2095_tmp = mux_1053_nl & ActUnitRun_wen;
  assign mux_1048_nl = MUX_s_1_2_2(or_tmp_1408, (~ mux_995_cse), and_2412_cse);
  assign mux_1049_nl = MUX_s_1_2_2(mux_1048_nl, or_tmp_1408, or_2025_cse);
  assign and_2093_tmp = (~ mux_1049_nl) & ActUnitRun_wen;
  assign mux_757_nl = MUX_s_1_2_2(mux_438_cse, and_2364_cse, or_1702_cse);
  assign and_1891_tmp = mux_757_nl & (~ (fsm_output[3])) & ActUnitRun_wen;
  assign nand_532_nl = ~((fsm_output[2:1]==2'b11) & or_1702_cse);
  assign mux_731_nl = MUX_s_1_2_2(nand_532_nl, or_3395_cse, fsm_output[3]);
  assign mux_732_nl = MUX_s_1_2_2(mux_731_nl, or_1831_cse, fsm_output[0]);
  assign and_1867_tmp = mux_732_nl & ActUnitRun_wen;
  assign and_1933_tmp = (and_2354_cse | (fsm_output[1:0]!=2'b10)) & (fsm_output[3:2]==2'b01)
      & ActUnitRun_wen;
  assign mux_1044_nl = MUX_s_1_2_2(or_tmp_1408, (~ mux_995_cse), and_2412_cse);
  assign mux_1045_nl = MUX_s_1_2_2(mux_1044_nl, or_tmp_1408, or_2017_cse);
  assign and_2091_tmp = (~ mux_1045_nl) & ActUnitRun_wen;
  assign mux_755_nl = MUX_s_1_2_2(mux_438_cse, and_2364_cse, nand_cse);
  assign and_1889_tmp = mux_755_nl & (~ (fsm_output[3])) & ActUnitRun_wen;
  assign or_1838_nl = (fsm_output[2:0]!=3'b110) | and_2354_cse;
  assign mux_730_nl = MUX_s_1_2_2(or_1838_nl, or_3395_cse, fsm_output[3]);
  assign and_1865_tmp = mux_730_nl & ActUnitRun_wen;
  assign mux_1024_nl = MUX_s_1_2_2(or_tmp_1408, (~ mux_995_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_1025_nl = MUX_s_1_2_2(mux_1024_nl, or_tmp_1408, or_1977_cse);
  assign and_2081_tmp = (~ mux_1025_nl) & ActUnitRun_wen;
  assign mux_1020_nl = MUX_s_1_2_2(or_tmp_1408, (~ mux_995_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_1021_nl = MUX_s_1_2_2(mux_1020_nl, or_tmp_1408, or_1969_cse);
  assign and_2079_tmp = (~ mux_1021_nl) & ActUnitRun_wen;
  assign nand_538_nl = ~((fsm_output[2:1]==2'b11) & ((ActUnit_PushOutput_if_for_i_4_0_sva_3_0!=4'b1001)));
  assign mux_741_nl = MUX_s_1_2_2(nand_538_nl, or_3395_cse, fsm_output[3]);
  assign mux_742_nl = MUX_s_1_2_2(mux_741_nl, or_1831_cse, fsm_output[0]);
  assign and_1877_tmp = mux_742_nl & ActUnitRun_wen;
  assign mux_1017_nl = MUX_s_1_2_2(mux_995_cse, nor_1586_cse, or_1961_cse);
  assign and_2077_tmp = mux_1017_nl & ActUnitRun_wen;
  assign mux_769_nl = MUX_s_1_2_2(mux_746_cse, and_2364_cse, or_1810_cse);
  assign and_1903_tmp = mux_769_nl & (~ (fsm_output[3])) & ActUnitRun_wen;
  assign nand_530_nl = ~((fsm_output[2:1]==2'b11) & or_1810_cse);
  assign mux_728_nl = MUX_s_1_2_2(nand_530_nl, or_3395_cse, fsm_output[3]);
  assign mux_729_nl = MUX_s_1_2_2(mux_728_nl, or_1831_cse, fsm_output[0]);
  assign and_1864_tmp = mux_729_nl & ActUnitRun_wen;
  assign mux_1014_nl = MUX_s_1_2_2(mux_995_cse, nor_1586_cse, or_1953_cse);
  assign and_2075_tmp = mux_1014_nl & ActUnitRun_wen;
  assign and_2387_nl = (ActUnit_PushOutput_if_for_i_4_0_sva_3_0==4'b0111);
  assign mux_767_nl = MUX_s_1_2_2(and_2364_cse, mux_438_cse, and_2387_nl);
  assign and_1901_tmp = mux_767_nl & (~ (fsm_output[3])) & ActUnitRun_wen;
  assign and_1878_nl = (fsm_output[2]) & ((ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3:2]!=2'b01)
      | nand_533_cse);
  assign mux_743_nl = MUX_s_1_2_2((fsm_output[2]), and_1878_nl, fsm_output[1]);
  assign mux_744_nl = MUX_s_1_2_2((~ mux_743_nl), or_3395_cse, fsm_output[3]);
  assign mux_745_nl = MUX_s_1_2_2(mux_744_nl, or_1831_cse, fsm_output[0]);
  assign and_1879_tmp = mux_745_nl & ActUnitRun_wen;
  assign mux_1011_nl = MUX_s_1_2_2(mux_995_cse, nor_1586_cse, or_1945_cse);
  assign and_2073_tmp = mux_1011_nl & ActUnitRun_wen;
  assign mux_765_nl = MUX_s_1_2_2(mux_438_cse, and_2364_cse, or_1798_cse);
  assign and_1899_tmp = mux_765_nl & (~ (fsm_output[3])) & ActUnitRun_wen;
  assign nand_537_nl = ~((fsm_output[2:1]==2'b11) & or_1798_cse);
  assign mux_739_nl = MUX_s_1_2_2(nand_537_nl, or_3395_cse, fsm_output[3]);
  assign mux_740_nl = MUX_s_1_2_2(mux_739_nl, or_1831_cse, fsm_output[0]);
  assign and_1875_tmp = mux_740_nl & ActUnitRun_wen;
  assign mux_1008_nl = MUX_s_1_2_2(mux_995_cse, nor_1586_cse, or_1937_cse);
  assign and_2071_tmp = mux_1008_nl & ActUnitRun_wen;
  assign nor_511_nl = ~((ActUnit_PushOutput_if_for_i_4_0_sva_3_0!=4'b0101));
  assign mux_763_nl = MUX_s_1_2_2(and_2364_cse, mux_438_cse, nor_511_nl);
  assign and_1897_tmp = mux_763_nl & (~ (fsm_output[3])) & ActUnitRun_wen;
  assign nand_536_nl = ~((fsm_output[2:1]==2'b11) & ((ActUnit_PushOutput_if_for_i_4_0_sva_3_0!=4'b0101)));
  assign mux_737_nl = MUX_s_1_2_2(nand_536_nl, or_3395_cse, fsm_output[3]);
  assign mux_738_nl = MUX_s_1_2_2(mux_737_nl, or_1831_cse, fsm_output[0]);
  assign and_1873_tmp = mux_738_nl & ActUnitRun_wen;
  assign mux_1005_nl = MUX_s_1_2_2(mux_995_cse, nor_1586_cse, or_1929_cse);
  assign and_2069_tmp = mux_1005_nl & ActUnitRun_wen;
  assign mux_761_nl = MUX_s_1_2_2(mux_438_cse, and_2364_cse, or_1750_cse);
  assign and_1895_tmp = mux_761_nl & (~ (fsm_output[3])) & ActUnitRun_wen;
  assign nand_535_nl = ~((fsm_output[2:1]==2'b11) & or_1750_cse);
  assign mux_735_nl = MUX_s_1_2_2(nand_535_nl, or_3395_cse, fsm_output[3]);
  assign mux_736_nl = MUX_s_1_2_2(mux_735_nl, or_1831_cse, fsm_output[0]);
  assign and_1871_tmp = mux_736_nl & ActUnitRun_wen;
  assign mux_1002_nl = MUX_s_1_2_2(mux_995_cse, nor_1586_cse, or_1921_cse);
  assign and_2067_tmp = mux_1002_nl & ActUnitRun_wen;
  assign nor_506_nl = ~((ActUnit_PushOutput_if_for_i_4_0_sva_3_0!=4'b0011));
  assign mux_759_nl = MUX_s_1_2_2(and_2364_cse, mux_438_cse, nor_506_nl);
  assign and_1893_tmp = mux_759_nl & (~ (fsm_output[3])) & ActUnitRun_wen;
  assign nand_534_nl = ~((fsm_output[2:1]==2'b11) & ((ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3:2]!=2'b00)
      | nand_533_cse));
  assign mux_733_nl = MUX_s_1_2_2(nand_534_nl, or_3395_cse, fsm_output[3]);
  assign mux_734_nl = MUX_s_1_2_2(mux_733_nl, or_1831_cse, fsm_output[0]);
  assign and_1869_tmp = mux_734_nl & ActUnitRun_wen;
  assign act_config_inst_counter_and_tmp = ActUnitRun_wen & ((and_dcpl_1082 & and_dcpl_1081
      & is_incr_lpi_1_dfm_1) | act_config_inst_counter_sva_mx0c1);
  assign or_943_nl = (fsm_output[1:0]!=2'b10);
  assign mux_447_nl = MUX_s_1_2_2(or_943_nl, or_tmp_484, fsm_output[3]);
  assign ActUnit_PushOutput_if_for_i_and_tmp = ActUnitRun_wen & ((~((z_out[4]) |
      and_dcpl_1112)) | ActUnit_PushOutput_if_for_i_4_0_sva_3_0_mx0c0 | (~(mux_447_nl
      | (fsm_output[2]))) | and_dcpl_331);
  assign ActUnit_RunLoad_if_a2_and_tmp = ActUnitRun_wen & (~ and_dcpl_1090) & and_dcpl_333
      & (~(act_config_is_zero_first_sva | act_config_is_zero_first_sva_dfm_4));
  assign and_1927_tmp = (and_2372_cse | (fsm_output[1:0]!=2'b10)) & (fsm_output[3:2]==2'b01)
      & ActUnitRun_wen;
  assign mux_1040_nl = MUX_s_1_2_2(or_tmp_1408, (~ mux_995_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_1041_nl = MUX_s_1_2_2(mux_1040_nl, or_tmp_1408, or_2009_cse);
  assign and_2089_tmp = (~ mux_1041_nl) & ActUnitRun_wen;
  assign mux_753_nl = MUX_s_1_2_2(and_2364_cse, mux_438_cse, and_2372_cse);
  assign and_1887_tmp = mux_753_nl & (~ (fsm_output[3])) & ActUnitRun_wen;
  assign and_2822_nl = (fsm_output[3:1]==3'b011) & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0==4'b1101);
  assign mux_1493_nl = MUX_s_1_2_2(and_2822_nl, nor_1654_cse, fsm_output[0]);
  assign or_3389_nl = (fsm_output[3:2]!=2'b01) | and_2372_cse;
  assign mux_1491_nl = MUX_s_1_2_2(or_1579_cse, or_3389_nl, fsm_output[1]);
  assign mux_1492_nl = MUX_s_1_2_2(mux_1491_nl, or_1831_cse, fsm_output[0]);
  assign mux_1494_nl = MUX_s_1_2_2(mux_1493_nl, mux_1492_nl, act_config_in_InstFetch_return_sva_7_2[2]);
  assign and_2328_tmp = mux_1494_nl & ActUnitRun_wen;
  assign and_1921_tmp = ((nor_1553_cse & (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3:2]==2'b11))
      | (fsm_output[1:0]!=2'b10)) & (fsm_output[3:2]==2'b01) & ActUnitRun_wen;
  assign mux_1036_nl = MUX_s_1_2_2(or_tmp_1408, (~ mux_995_cse), ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]);
  assign mux_1037_nl = MUX_s_1_2_2(mux_1036_nl, or_tmp_1408, or_2001_cse);
  assign and_2087_tmp = (~ mux_1037_nl) & ActUnitRun_wen;
  assign mux_751_nl = MUX_s_1_2_2(mux_746_cse, and_2364_cse, or_1714_cse);
  assign and_1885_tmp = mux_751_nl & (~ (fsm_output[3])) & ActUnitRun_wen;
  assign nor_1665_nl = ~((fsm_output[3:1]!=3'b011) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0!=4'b1100));
  assign mux_1489_nl = MUX_s_1_2_2(nor_1665_nl, nor_1654_cse, fsm_output[0]);
  assign or_3380_nl = (fsm_output[3:2]!=2'b01) | (~((ActUnit_PushOutput_if_for_i_4_0_sva_3_0!=4'b1100)));
  assign mux_1487_nl = MUX_s_1_2_2(or_1579_cse, or_3380_nl, fsm_output[1]);
  assign mux_1488_nl = MUX_s_1_2_2(mux_1487_nl, or_1831_cse, fsm_output[0]);
  assign mux_1490_nl = MUX_s_1_2_2(mux_1489_nl, mux_1488_nl, act_config_in_InstFetch_return_sva_7_2[2]);
  assign and_2327_tmp = mux_1490_nl & ActUnitRun_wen;
  assign and_1915_tmp = (and_2367_cse | (fsm_output[1:0]!=2'b10)) & (fsm_output[3:2]==2'b01)
      & ActUnitRun_wen;
  assign mux_1032_nl = MUX_s_1_2_2(or_tmp_1408, (~ mux_995_cse), and_2412_cse);
  assign mux_1033_nl = MUX_s_1_2_2(mux_1032_nl, or_tmp_1408, or_1993_cse);
  assign and_2085_tmp = (~ mux_1033_nl) & ActUnitRun_wen;
  assign mux_749_nl = MUX_s_1_2_2(and_2364_cse, mux_746_cse, and_2367_cse);
  assign and_1883_tmp = mux_749_nl & (~ (fsm_output[3])) & ActUnitRun_wen;
  assign nor_1661_nl = ~((fsm_output[3:1]!=3'b011) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2])
      | not_tmp_2198);
  assign mux_1485_nl = MUX_s_1_2_2(nor_1661_nl, nor_1654_cse, fsm_output[0]);
  assign or_3370_nl = (fsm_output[3:2]!=2'b01) | (~((ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2])
      | not_tmp_2198));
  assign mux_1483_nl = MUX_s_1_2_2(or_1579_cse, or_3370_nl, fsm_output[1]);
  assign mux_1484_nl = MUX_s_1_2_2(mux_1483_nl, or_1831_cse, fsm_output[0]);
  assign mux_1486_nl = MUX_s_1_2_2(mux_1485_nl, mux_1484_nl, act_config_in_InstFetch_return_sva_7_2[2]);
  assign and_2326_tmp = mux_1486_nl & ActUnitRun_wen;
  assign and_1909_tmp = (((ActUnit_PushOutput_if_for_i_4_0_sva_3_0==4'b1010)) | (fsm_output[1:0]!=2'b10))
      & (fsm_output[3:2]==2'b01) & ActUnitRun_wen;
  assign mux_1028_nl = MUX_s_1_2_2(or_tmp_1408, (~ mux_995_cse), and_2412_cse);
  assign mux_1029_nl = MUX_s_1_2_2(mux_1028_nl, or_tmp_1408, or_1985_cse);
  assign and_2083_tmp = (~ mux_1029_nl) & ActUnitRun_wen;
  assign mux_747_nl = MUX_s_1_2_2(mux_746_cse, and_2364_cse, or_1762_cse);
  assign and_1881_tmp = mux_747_nl & (~ (fsm_output[3])) & ActUnitRun_wen;
  assign nor_1657_nl = ~((fsm_output[3:1]!=3'b011) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0!=4'b1010));
  assign mux_1481_nl = MUX_s_1_2_2(nor_1657_nl, nor_1654_cse, fsm_output[0]);
  assign or_3360_nl = (fsm_output[3:2]!=2'b01) | (~((ActUnit_PushOutput_if_for_i_4_0_sva_3_0!=4'b1010)));
  assign mux_1479_nl = MUX_s_1_2_2(or_1579_cse, or_3360_nl, fsm_output[1]);
  assign mux_1480_nl = MUX_s_1_2_2(mux_1479_nl, or_1831_cse, fsm_output[0]);
  assign mux_1482_nl = MUX_s_1_2_2(mux_1481_nl, mux_1480_nl, act_config_in_InstFetch_return_sva_7_2[2]);
  assign and_2325_tmp = mux_1482_nl & ActUnitRun_wen;
  assign and_2329_nl = (fsm_output[2]) & ((fsm_output[1:0]!=2'b10) | nor_1406_cse);
  assign mux_590_nl = MUX_s_1_2_2(and_2329_nl, nor_1405_cse, fsm_output[3]);
  assign and_1803_tmp = mux_590_nl & ActUnitRun_wen;
  assign mux_999_nl = MUX_s_1_2_2(mux_995_cse, nor_1586_cse, or_1913_cse);
  assign and_2065_tmp = mux_999_nl & ActUnitRun_wen;
  assign nor_1404_nl = ~((fsm_output[2:1]!=2'b11) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0!=4'b0001));
  assign mux_588_nl = MUX_s_1_2_2(nor_1404_nl, or_3395_cse, fsm_output[0]);
  assign mux_589_nl = MUX_s_1_2_2(mux_588_nl, nor_1405_cse, fsm_output[3]);
  assign and_1801_tmp = mux_589_nl & ActUnitRun_wen;
  assign nor_1653_nl = ~((fsm_output[3:1]!=3'b011) | (ActUnit_PushOutput_if_for_i_4_0_sva_3_0!=4'b0001));
  assign mux_1477_nl = MUX_s_1_2_2(nor_1653_nl, nor_1654_cse, fsm_output[0]);
  assign or_3350_nl = (fsm_output[3:2]!=2'b01) | nor_1406_cse;
  assign mux_1475_nl = MUX_s_1_2_2(or_1579_cse, or_3350_nl, fsm_output[1]);
  assign mux_1476_nl = MUX_s_1_2_2(mux_1475_nl, or_1831_cse, fsm_output[0]);
  assign mux_1478_nl = MUX_s_1_2_2(mux_1477_nl, mux_1476_nl, act_config_in_InstFetch_return_sva_7_2[2]);
  assign and_2324_tmp = mux_1478_nl & ActUnitRun_wen;
  assign mux_625_nl = MUX_s_1_2_2((~ (fsm_output[2])), (fsm_output[2]), fsm_output[3]);
  assign mux_626_nl = MUX_s_1_2_2(mux_625_nl, or_tmp_552, fsm_output[0]);
  assign mux_627_nl = MUX_s_1_2_2(or_tmp_555, mux_626_nl, fsm_output[1]);
  assign mux_623_nl = MUX_s_1_2_2(or_1579_cse, or_tmp_552, fsm_output[0]);
  assign mux_624_nl = MUX_s_1_2_2(or_tmp_555, mux_623_nl, fsm_output[1]);
  assign mux_628_nl = MUX_s_1_2_2(mux_627_nl, mux_624_nl, or_1427_cse);
  assign and_1808_tmp = (~ mux_628_nl) & ActUnitRun_wen;
  assign mux_996_nl = MUX_s_1_2_2(mux_995_cse, nor_1586_cse, or_1905_cse);
  assign and_2063_tmp = mux_996_nl & ActUnitRun_wen;
  assign or_1429_nl = (fsm_output[2:0]!=3'b100);
  assign mux_453_nl = MUX_s_1_2_2(or_1429_nl, or_3395_cse, fsm_output[3]);
  assign or_1428_nl = (~ (fsm_output[2])) | (fsm_output[0]);
  assign mux_452_nl = MUX_s_1_2_2(or_1428_nl, or_3395_cse, fsm_output[3]);
  assign mux_454_nl = MUX_s_1_2_2(mux_453_nl, mux_452_nl, or_1427_cse);
  assign rva_out_reg_data_and_61_tmp = rva_out_reg_data_and_ssc & mux_454_nl;
  assign Silu_for_else_else_else_if_and_tmp = Silu_for_else_else_else_if_and_2_ssc
      & (and_dcpl_1112 | and_dcpl_1390 | and_dcpl_1236 | (~ Silu_for_else_else_else_if_or_13_rgt));
  assign nl_Silu_for_12_else_else_else_else_if_acc_sdt = ({reg_nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1})
      + 4'b1111;
  assign Silu_for_12_else_else_else_else_if_acc_sdt = nl_Silu_for_12_else_else_else_else_if_acc_sdt[3:0];
  assign nl_Silu_for_13_else_else_else_else_if_acc_sdt = ({reg_nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1})
      + 4'b1111;
  assign Silu_for_13_else_else_else_else_if_acc_sdt = nl_Silu_for_13_else_else_else_else_if_acc_sdt[3:0];
  assign and_1715_ssc = and_dcpl_1236 & (~ or_1527_tmp);
  assign nl_Silu_for_14_else_else_else_else_if_acc_sdt = ({reg_nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1})
      + 4'b1111;
  assign Silu_for_14_else_else_else_else_if_acc_sdt = nl_Silu_for_14_else_else_else_else_if_acc_sdt[3:0];
  assign nl_Silu_for_15_else_else_else_else_if_acc_sdt = ({reg_nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1})
      + 4'b1111;
  assign Silu_for_15_else_else_else_else_if_acc_sdt = nl_Silu_for_15_else_else_else_else_if_acc_sdt[3:0];
  assign nl_Silu_for_16_else_else_else_else_if_acc_sdt = ({reg_nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1})
      + 4'b1111;
  assign Silu_for_16_else_else_else_else_if_acc_sdt = nl_Silu_for_16_else_else_else_else_if_acc_sdt[3:0];
  assign nl_Silu_for_1_else_else_else_else_if_acc_sdt = ({reg_ActUnit_RunInst_case_14_nv_scvector_cctor_data_0_1_ftd_rsp_0
      , reg_ActUnit_RunInst_case_14_nv_scvector_cctor_data_0_1_ftd_rsp_1}) + 4'b1111;
  assign Silu_for_1_else_else_else_else_if_acc_sdt = nl_Silu_for_1_else_else_else_else_if_acc_sdt[3:0];
  assign nl_Silu_for_2_else_else_else_else_if_acc_sdt = ({reg_nv_scvector_cctor_nv_scvector_5_for_2_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_2_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1})
      + 4'b1111;
  assign Silu_for_2_else_else_else_else_if_acc_sdt = nl_Silu_for_2_else_else_else_else_if_acc_sdt[3:0];
  assign nl_Silu_for_3_else_else_else_else_if_acc_sdt = ({reg_nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1})
      + 4'b1111;
  assign Silu_for_3_else_else_else_else_if_acc_sdt = nl_Silu_for_3_else_else_else_else_if_acc_sdt[3:0];
  assign nl_Silu_for_4_else_else_else_else_if_acc_sdt = ({reg_nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1})
      + 4'b1111;
  assign Silu_for_4_else_else_else_else_if_acc_sdt = nl_Silu_for_4_else_else_else_else_if_acc_sdt[3:0];
  assign nl_Silu_for_5_else_else_else_else_if_acc_sdt = ({reg_nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1})
      + 4'b1111;
  assign Silu_for_5_else_else_else_else_if_acc_sdt = nl_Silu_for_5_else_else_else_else_if_acc_sdt[3:0];
  assign nl_Silu_for_6_else_else_else_else_if_acc_sdt = ({reg_nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1})
      + 4'b1111;
  assign Silu_for_6_else_else_else_else_if_acc_sdt = nl_Silu_for_6_else_else_else_else_if_acc_sdt[3:0];
  assign nl_Silu_for_7_else_else_else_else_if_acc_sdt = ({reg_nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1})
      + 4'b1111;
  assign Silu_for_7_else_else_else_else_if_acc_sdt = nl_Silu_for_7_else_else_else_else_if_acc_sdt[3:0];
  assign nl_Silu_for_8_else_else_else_else_if_acc_sdt = ({reg_nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1})
      + 4'b1111;
  assign Silu_for_8_else_else_else_else_if_acc_sdt = nl_Silu_for_8_else_else_else_else_if_acc_sdt[3:0];
  assign nl_Silu_for_9_else_else_else_else_if_acc_sdt = ({reg_nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1})
      + 4'b1111;
  assign Silu_for_9_else_else_else_else_if_acc_sdt = nl_Silu_for_9_else_else_else_else_if_acc_sdt[3:0];
  assign nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      = MUX_s_1_4_2(reg_act_regs_data_0_0_ftd_2_3, act_regs_data_1_0_sva_25, act_regs_data_2_0_sva_25,
      act_regs_data_3_0_sva_25, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      = MUX_v_3_4_2(reg_act_regs_data_0_0_ftd_2_2_0, act_regs_data_1_0_sva_24_22,
      act_regs_data_2_0_sva_24_22, act_regs_data_3_0_sva_24_22, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      = MUX_s_1_4_2(reg_act_regs_data_0_1_ftd_2_3, act_regs_data_1_1_sva_25, act_regs_data_2_1_sva_25,
      act_regs_data_3_1_sva_25, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      = MUX_v_3_4_2(reg_act_regs_data_0_1_ftd_2_2_0, act_regs_data_1_1_sva_24_22,
      act_regs_data_2_1_sva_24_22, act_regs_data_3_1_sva_24_22, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      = MUX_s_1_4_2(act_regs_data_0_2_sva_25, act_regs_data_1_2_sva_25, act_regs_data_2_2_sva_25,
      act_regs_data_3_2_sva_25, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      = MUX_v_3_4_2(act_regs_data_0_2_sva_24_22, act_regs_data_1_2_sva_24_22, act_regs_data_2_2_sva_24_22,
      act_regs_data_3_2_sva_24_22, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      = MUX_s_1_4_2(act_regs_data_0_3_sva_25, act_regs_data_1_3_sva_25, act_regs_data_2_3_sva_25,
      act_regs_data_3_3_sva_25, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      = MUX_v_3_4_2(act_regs_data_0_3_sva_24_22, act_regs_data_1_3_sva_24_22, act_regs_data_2_3_sva_24_22,
      act_regs_data_3_3_sva_24_22, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      = MUX_s_1_4_2(act_regs_data_0_4_sva_25, act_regs_data_1_4_sva_25, act_regs_data_2_4_sva_25,
      act_regs_data_3_4_sva_25, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      = MUX_v_3_4_2(act_regs_data_0_4_sva_24_22, act_regs_data_1_4_sva_24_22, act_regs_data_2_4_sva_24_22,
      act_regs_data_3_4_sva_24_22, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      = MUX_s_1_4_2(act_regs_data_0_5_sva_25, act_regs_data_1_5_sva_25, act_regs_data_2_5_sva_25,
      act_regs_data_3_5_sva_25, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      = MUX_v_3_4_2(act_regs_data_0_5_sva_24_22, act_regs_data_1_5_sva_24_22, act_regs_data_2_5_sva_24_22,
      act_regs_data_3_5_sva_24_22, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      = MUX_s_1_4_2(act_regs_data_0_6_sva_25, act_regs_data_1_6_sva_25, act_regs_data_2_6_sva_25,
      act_regs_data_3_6_sva_25, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      = MUX_v_3_4_2(act_regs_data_0_6_sva_24_22, act_regs_data_1_6_sva_24_22, act_regs_data_2_6_sva_24_22,
      act_regs_data_3_6_sva_24_22, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      = MUX_s_1_4_2(act_regs_data_0_7_sva_25, act_regs_data_1_7_sva_25, act_regs_data_2_7_sva_25,
      act_regs_data_3_7_sva_25, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      = MUX_v_3_4_2(act_regs_data_0_7_sva_24_22, act_regs_data_1_7_sva_24_22, act_regs_data_2_7_sva_24_22,
      act_regs_data_3_7_sva_24_22, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      = MUX_s_1_4_2(act_regs_data_0_8_sva_25, act_regs_data_1_8_sva_25, act_regs_data_2_8_sva_25,
      act_regs_data_3_8_sva_25, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      = MUX_v_3_4_2(act_regs_data_0_8_sva_24_22, act_regs_data_1_8_sva_24_22, act_regs_data_2_8_sva_24_22,
      act_regs_data_3_8_sva_24_22, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      = MUX_s_1_4_2(act_regs_data_0_9_sva_25, act_regs_data_1_9_sva_25, act_regs_data_2_9_sva_25,
      act_regs_data_3_9_sva_25, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      = MUX_v_3_4_2(act_regs_data_0_9_sva_24_22, act_regs_data_1_9_sva_24_22, act_regs_data_2_9_sva_24_22,
      act_regs_data_3_9_sva_24_22, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      = MUX_s_1_4_2(reg_act_regs_data_0_10_ftd_2_3, act_regs_data_1_10_sva_25, act_regs_data_2_10_sva_25,
      act_regs_data_3_10_sva_25, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      = MUX_v_3_4_2(reg_act_regs_data_0_10_ftd_2_2_0, act_regs_data_1_10_sva_24_22,
      act_regs_data_2_10_sva_24_22, act_regs_data_3_10_sva_24_22, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      = MUX_s_1_4_2(reg_act_regs_data_0_11_ftd_2_3, act_regs_data_1_11_sva_25, act_regs_data_2_11_sva_25,
      act_regs_data_3_11_sva_25, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      = MUX_v_3_4_2(reg_act_regs_data_0_11_ftd_2_2_0, act_regs_data_1_11_sva_24_22,
      act_regs_data_2_11_sva_24_22, act_regs_data_3_11_sva_24_22, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      = MUX_s_1_4_2(reg_act_regs_data_0_12_ftd_2_3, act_regs_data_1_12_sva_25, act_regs_data_2_12_sva_25,
      act_regs_data_3_12_sva_25, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      = MUX_v_3_4_2(reg_act_regs_data_0_12_ftd_2_2_0, act_regs_data_1_12_sva_24_22,
      act_regs_data_2_12_sva_24_22, act_regs_data_3_12_sva_24_22, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      = MUX_s_1_4_2(reg_act_regs_data_0_13_ftd_2_3, act_regs_data_1_13_sva_25, act_regs_data_2_13_sva_25,
      act_regs_data_3_13_sva_25, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      = MUX_v_3_4_2(reg_act_regs_data_0_13_ftd_2_2_0, act_regs_data_1_13_sva_24_22,
      act_regs_data_2_13_sva_24_22, act_regs_data_3_13_sva_24_22, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      = MUX_s_1_4_2(act_regs_data_0_14_sva_25, act_regs_data_1_14_sva_25, act_regs_data_2_14_sva_25,
      act_regs_data_3_14_sva_25, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      = MUX_v_3_4_2(act_regs_data_0_14_sva_24_22, act_regs_data_1_14_sva_24_22, act_regs_data_2_14_sva_24_22,
      act_regs_data_3_14_sva_24_22, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
      = MUX_s_1_4_2(act_regs_data_0_15_sva_25, act_regs_data_1_15_sva_25, act_regs_data_2_15_sva_25,
      act_regs_data_3_15_sva_25, act_config_in_InstFetch_mux_tmp[3:2]);
  assign nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
      = MUX_v_3_4_2(act_regs_data_0_15_sva_24_22, act_regs_data_1_15_sva_24_22, act_regs_data_2_15_sva_24_22,
      act_regs_data_3_15_sva_24_22, act_config_in_InstFetch_mux_tmp[3:2]);
  assign ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_25 = MUX_s_1_64_2(reg_act_regs_data_0_0_ftd_2_3,
      reg_act_regs_data_0_1_ftd_2_3, act_regs_data_0_2_sva_25, act_regs_data_0_3_sva_25,
      act_regs_data_0_4_sva_25, act_regs_data_0_5_sva_25, act_regs_data_0_6_sva_25,
      act_regs_data_0_7_sva_25, act_regs_data_0_8_sva_25, act_regs_data_0_9_sva_25,
      reg_act_regs_data_0_10_ftd_2_3, reg_act_regs_data_0_11_ftd_2_3, reg_act_regs_data_0_12_ftd_2_3,
      reg_act_regs_data_0_13_ftd_2_3, act_regs_data_0_14_sva_25, act_regs_data_0_15_sva_25,
      act_regs_data_1_0_sva_25, act_regs_data_1_1_sva_25, act_regs_data_1_2_sva_25,
      act_regs_data_1_3_sva_25, act_regs_data_1_4_sva_25, act_regs_data_1_5_sva_25,
      act_regs_data_1_6_sva_25, act_regs_data_1_7_sva_25, act_regs_data_1_8_sva_25,
      act_regs_data_1_9_sva_25, act_regs_data_1_10_sva_25, act_regs_data_1_11_sva_25,
      act_regs_data_1_12_sva_25, act_regs_data_1_13_sva_25, act_regs_data_1_14_sva_25,
      act_regs_data_1_15_sva_25, act_regs_data_2_0_sva_25, act_regs_data_2_1_sva_25,
      act_regs_data_2_2_sva_25, act_regs_data_2_3_sva_25, act_regs_data_2_4_sva_25,
      act_regs_data_2_5_sva_25, act_regs_data_2_6_sva_25, act_regs_data_2_7_sva_25,
      act_regs_data_2_8_sva_25, act_regs_data_2_9_sva_25, act_regs_data_2_10_sva_25,
      act_regs_data_2_11_sva_25, act_regs_data_2_12_sva_25, act_regs_data_2_13_sva_25,
      act_regs_data_2_14_sva_25, act_regs_data_2_15_sva_25, act_regs_data_3_0_sva_25,
      act_regs_data_3_1_sva_25, act_regs_data_3_2_sva_25, act_regs_data_3_3_sva_25,
      act_regs_data_3_4_sva_25, act_regs_data_3_5_sva_25, act_regs_data_3_6_sva_25,
      act_regs_data_3_7_sva_25, act_regs_data_3_8_sva_25, act_regs_data_3_9_sva_25,
      act_regs_data_3_10_sva_25, act_regs_data_3_11_sva_25, act_regs_data_3_12_sva_25,
      act_regs_data_3_13_sva_25, act_regs_data_3_14_sva_25, act_regs_data_3_15_sva_25,
      {(act_config_in_InstFetch_return_sva_7_2[1:0]) , ActUnit_PushOutput_if_for_i_4_0_sva_3_0});
  assign ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_24_22
      = MUX_v_3_64_2(reg_act_regs_data_0_0_ftd_2_2_0, reg_act_regs_data_0_1_ftd_2_2_0,
      act_regs_data_0_2_sva_24_22, act_regs_data_0_3_sva_24_22, act_regs_data_0_4_sva_24_22,
      act_regs_data_0_5_sva_24_22, act_regs_data_0_6_sva_24_22, act_regs_data_0_7_sva_24_22,
      act_regs_data_0_8_sva_24_22, act_regs_data_0_9_sva_24_22, reg_act_regs_data_0_10_ftd_2_2_0,
      reg_act_regs_data_0_11_ftd_2_2_0, reg_act_regs_data_0_12_ftd_2_2_0, reg_act_regs_data_0_13_ftd_2_2_0,
      act_regs_data_0_14_sva_24_22, act_regs_data_0_15_sva_24_22, act_regs_data_1_0_sva_24_22,
      act_regs_data_1_1_sva_24_22, act_regs_data_1_2_sva_24_22, act_regs_data_1_3_sva_24_22,
      act_regs_data_1_4_sva_24_22, act_regs_data_1_5_sva_24_22, act_regs_data_1_6_sva_24_22,
      act_regs_data_1_7_sva_24_22, act_regs_data_1_8_sva_24_22, act_regs_data_1_9_sva_24_22,
      act_regs_data_1_10_sva_24_22, act_regs_data_1_11_sva_24_22, act_regs_data_1_12_sva_24_22,
      act_regs_data_1_13_sva_24_22, act_regs_data_1_14_sva_24_22, act_regs_data_1_15_sva_24_22,
      act_regs_data_2_0_sva_24_22, act_regs_data_2_1_sva_24_22, act_regs_data_2_2_sva_24_22,
      act_regs_data_2_3_sva_24_22, act_regs_data_2_4_sva_24_22, act_regs_data_2_5_sva_24_22,
      act_regs_data_2_6_sva_24_22, act_regs_data_2_7_sva_24_22, act_regs_data_2_8_sva_24_22,
      act_regs_data_2_9_sva_24_22, act_regs_data_2_10_sva_24_22, act_regs_data_2_11_sva_24_22,
      act_regs_data_2_12_sva_24_22, act_regs_data_2_13_sva_24_22, act_regs_data_2_14_sva_24_22,
      act_regs_data_2_15_sva_24_22, act_regs_data_3_0_sva_24_22, act_regs_data_3_1_sva_24_22,
      act_regs_data_3_2_sva_24_22, act_regs_data_3_3_sva_24_22, act_regs_data_3_4_sva_24_22,
      act_regs_data_3_5_sva_24_22, act_regs_data_3_6_sva_24_22, act_regs_data_3_7_sva_24_22,
      act_regs_data_3_8_sva_24_22, act_regs_data_3_9_sva_24_22, act_regs_data_3_10_sva_24_22,
      act_regs_data_3_11_sva_24_22, act_regs_data_3_12_sva_24_22, act_regs_data_3_13_sva_24_22,
      act_regs_data_3_14_sva_24_22, act_regs_data_3_15_sva_24_22, {(act_config_in_InstFetch_return_sva_7_2[1:0])
      , ActUnit_PushOutput_if_for_i_4_0_sva_3_0});
  assign ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_25_22_mx0w2_3
      = MUX_s_1_64_2(act_regs_data_0_0_sva_dfm_2_25_22_rsp_0, act_regs_data_0_1_sva_dfm_2_25_22_rsp_0,
      act_regs_data_0_2_sva_dfm_2_25_22_rsp_0, act_regs_data_0_3_sva_dfm_2_25_22_rsp_0,
      act_regs_data_0_4_sva_dfm_2_25_22_rsp_0, act_regs_data_0_5_sva_dfm_2_25_22_rsp_0,
      act_regs_data_0_6_sva_dfm_2_25_22_rsp_0, act_regs_data_0_7_sva_dfm_2_25_22_rsp_0,
      act_regs_data_0_8_sva_dfm_2_25_22_rsp_0, act_regs_data_0_9_sva_dfm_2_25_22_rsp_0,
      act_regs_data_0_10_sva_dfm_2_25_22_rsp_0, act_regs_data_0_11_sva_dfm_2_25_22_rsp_0,
      act_regs_data_0_12_sva_dfm_2_25_22_rsp_0, act_regs_data_0_13_sva_dfm_2_25_22_rsp_0,
      act_regs_data_0_14_sva_dfm_2_25_22_rsp_0, act_regs_data_0_15_sva_dfm_2_25_22_rsp_0,
      act_regs_data_1_0_sva_dfm_2_25_22_rsp_0, act_regs_data_1_1_sva_dfm_2_25_22_rsp_0,
      act_regs_data_1_2_sva_dfm_2_25_22_rsp_0, act_regs_data_1_3_sva_dfm_2_25_22_rsp_0,
      act_regs_data_1_4_sva_dfm_2_25_22_rsp_0, act_regs_data_1_5_sva_dfm_2_25_22_rsp_0,
      act_regs_data_1_6_sva_dfm_2_25_22_rsp_0, act_regs_data_1_7_sva_dfm_2_25_22_rsp_0,
      act_regs_data_1_8_sva_dfm_2_25_22_rsp_0, act_regs_data_1_9_sva_dfm_2_25_22_rsp_0,
      act_regs_data_1_10_sva_dfm_2_25_22_rsp_0, act_regs_data_1_11_sva_dfm_2_25_22_rsp_0,
      act_regs_data_1_12_sva_dfm_2_25_22_rsp_0, act_regs_data_1_13_sva_dfm_2_25_22_rsp_0,
      act_regs_data_1_14_sva_dfm_2_25_22_rsp_0, act_regs_data_1_15_sva_dfm_2_25_22_rsp_0,
      act_regs_data_2_0_sva_dfm_2_25_22_rsp_0, act_regs_data_2_1_sva_dfm_2_25_22_rsp_0,
      act_regs_data_2_2_sva_dfm_2_25_22_rsp_0, act_regs_data_2_3_sva_dfm_2_25_22_rsp_0,
      act_regs_data_2_4_sva_dfm_2_25_22_rsp_0, act_regs_data_2_5_sva_dfm_2_25_22_rsp_0,
      act_regs_data_2_6_sva_dfm_2_25_22_rsp_0, act_regs_data_2_7_sva_dfm_2_25_22_rsp_0,
      act_regs_data_2_8_sva_dfm_2_25_22_rsp_0, act_regs_data_2_9_sva_dfm_2_25_22_rsp_0,
      act_regs_data_2_10_sva_dfm_2_25_22_rsp_0, act_regs_data_2_11_sva_dfm_2_25_22_rsp_0,
      act_regs_data_2_12_sva_dfm_2_25_22_rsp_0, act_regs_data_2_13_sva_dfm_2_25_22_rsp_0,
      act_regs_data_2_14_sva_dfm_2_25_22_rsp_0, act_regs_data_2_15_sva_dfm_2_25_22_rsp_0,
      act_regs_data_3_0_sva_dfm_2_25_22_rsp_0, act_regs_data_3_1_sva_dfm_2_25_22_rsp_0,
      act_regs_data_3_2_sva_dfm_2_25_22_rsp_0, act_regs_data_3_3_sva_dfm_2_25_22_rsp_0,
      act_regs_data_3_4_sva_dfm_2_25_22_rsp_0, act_regs_data_3_5_sva_dfm_2_25_22_rsp_0,
      act_regs_data_3_6_sva_dfm_2_25_22_rsp_0, act_regs_data_3_7_sva_dfm_2_25_22_rsp_0,
      act_regs_data_3_8_sva_dfm_2_25_22_rsp_0, act_regs_data_3_9_sva_dfm_2_25_22_rsp_0,
      act_regs_data_3_10_sva_dfm_2_25_22_rsp_0, act_regs_data_3_11_sva_dfm_2_25_22_rsp_0,
      act_regs_data_3_12_sva_dfm_2_25_22_rsp_0, act_regs_data_3_13_sva_dfm_2_25_22_rsp_0,
      act_regs_data_3_14_sva_dfm_2_25_22_rsp_0, act_regs_data_3_15_sva_dfm_2_25_22_rsp_0,
      {nvhls_get_slc_2U_NVUINT8_return_2_sva , ActUnit_PushOutput_if_for_i_4_0_sva_3_0});
  assign ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_25_22_mx0w2_2_0
      = MUX_v_3_64_2(act_regs_data_0_0_sva_dfm_2_25_22_rsp_1, act_regs_data_0_1_sva_dfm_2_25_22_rsp_1,
      act_regs_data_0_2_sva_dfm_2_25_22_rsp_1, act_regs_data_0_3_sva_dfm_2_25_22_rsp_1,
      act_regs_data_0_4_sva_dfm_2_25_22_rsp_1, act_regs_data_0_5_sva_dfm_2_25_22_rsp_1,
      act_regs_data_0_6_sva_dfm_2_25_22_rsp_1, act_regs_data_0_7_sva_dfm_2_25_22_rsp_1,
      act_regs_data_0_8_sva_dfm_2_25_22_rsp_1, act_regs_data_0_9_sva_dfm_2_25_22_rsp_1,
      act_regs_data_0_10_sva_dfm_2_25_22_rsp_1, act_regs_data_0_11_sva_dfm_2_25_22_rsp_1,
      act_regs_data_0_12_sva_dfm_2_25_22_rsp_1, act_regs_data_0_13_sva_dfm_2_25_22_rsp_1,
      act_regs_data_0_14_sva_dfm_2_25_22_rsp_1, act_regs_data_0_15_sva_dfm_2_25_22_rsp_1,
      act_regs_data_1_0_sva_dfm_2_25_22_rsp_1, act_regs_data_1_1_sva_dfm_2_25_22_rsp_1,
      act_regs_data_1_2_sva_dfm_2_25_22_rsp_1, act_regs_data_1_3_sva_dfm_2_25_22_rsp_1,
      act_regs_data_1_4_sva_dfm_2_25_22_rsp_1, act_regs_data_1_5_sva_dfm_2_25_22_rsp_1,
      act_regs_data_1_6_sva_dfm_2_25_22_rsp_1, act_regs_data_1_7_sva_dfm_2_25_22_rsp_1,
      act_regs_data_1_8_sva_dfm_2_25_22_rsp_1, act_regs_data_1_9_sva_dfm_2_25_22_rsp_1,
      act_regs_data_1_10_sva_dfm_2_25_22_rsp_1, act_regs_data_1_11_sva_dfm_2_25_22_rsp_1,
      act_regs_data_1_12_sva_dfm_2_25_22_rsp_1, act_regs_data_1_13_sva_dfm_2_25_22_rsp_1,
      act_regs_data_1_14_sva_dfm_2_25_22_rsp_1, act_regs_data_1_15_sva_dfm_2_25_22_rsp_1,
      act_regs_data_2_0_sva_dfm_2_25_22_rsp_1, act_regs_data_2_1_sva_dfm_2_25_22_rsp_1,
      act_regs_data_2_2_sva_dfm_2_25_22_rsp_1, act_regs_data_2_3_sva_dfm_2_25_22_rsp_1,
      act_regs_data_2_4_sva_dfm_2_25_22_rsp_1, act_regs_data_2_5_sva_dfm_2_25_22_rsp_1,
      act_regs_data_2_6_sva_dfm_2_25_22_rsp_1, act_regs_data_2_7_sva_dfm_2_25_22_rsp_1,
      act_regs_data_2_8_sva_dfm_2_25_22_rsp_1, act_regs_data_2_9_sva_dfm_2_25_22_rsp_1,
      act_regs_data_2_10_sva_dfm_2_25_22_rsp_1, act_regs_data_2_11_sva_dfm_2_25_22_rsp_1,
      act_regs_data_2_12_sva_dfm_2_25_22_rsp_1, act_regs_data_2_13_sva_dfm_2_25_22_rsp_1,
      act_regs_data_2_14_sva_dfm_2_25_22_rsp_1, act_regs_data_2_15_sva_dfm_2_25_22_rsp_1,
      act_regs_data_3_0_sva_dfm_2_25_22_rsp_1, act_regs_data_3_1_sva_dfm_2_25_22_rsp_1,
      act_regs_data_3_2_sva_dfm_2_25_22_rsp_1, act_regs_data_3_3_sva_dfm_2_25_22_rsp_1,
      act_regs_data_3_4_sva_dfm_2_25_22_rsp_1, act_regs_data_3_5_sva_dfm_2_25_22_rsp_1,
      act_regs_data_3_6_sva_dfm_2_25_22_rsp_1, act_regs_data_3_7_sva_dfm_2_25_22_rsp_1,
      act_regs_data_3_8_sva_dfm_2_25_22_rsp_1, act_regs_data_3_9_sva_dfm_2_25_22_rsp_1,
      act_regs_data_3_10_sva_dfm_2_25_22_rsp_1, act_regs_data_3_11_sva_dfm_2_25_22_rsp_1,
      act_regs_data_3_12_sva_dfm_2_25_22_rsp_1, act_regs_data_3_13_sva_dfm_2_25_22_rsp_1,
      act_regs_data_3_14_sva_dfm_2_25_22_rsp_1, act_regs_data_3_15_sva_dfm_2_25_22_rsp_1,
      {nvhls_get_slc_2U_NVUINT8_return_2_sva , ActUnit_PushOutput_if_for_i_4_0_sva_3_0});
  assign Silu_for_else_Silu_for_else_mux1h_31_nl = MUX1HOT_s_1_4_2((Silu_for_y_1_sva_1_22_0_1[22]),
      (Silu_for_16_else_else_if_acc_itm[1]), ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_1_25,
      reg_nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0,
      {(~ Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_30_ssc_1 , Silu_for_else_else_else_and_30_ssc_1 , Silu_for_else_else_else_and_31_ssc_1});
  assign Silu_for_y_lpi_1_dfm_4_25 = Silu_for_else_Silu_for_else_mux1h_31_nl & (~
      Silu_for_else_and_47_ssc_1) & Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  assign Silu_for_else_Silu_for_else_mux1h_65_nl = MUX1HOT_v_3_5_2((signext_3_1(Silu_for_y_1_sva_1_22_0_1[22])),
      ({{1{Silu_for_16_else_else_if_acc_itm[1]}}, Silu_for_16_else_else_if_acc_itm}),
      reg_Silu_for_16_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd,
      ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_1_24_22, reg_nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1,
      {(~ Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_30_ssc_1 , Silu_for_else_and_47_ssc_1 , Silu_for_else_else_else_and_30_ssc_1
      , Silu_for_else_else_else_and_31_ssc_1});
  assign Silu_for_y_lpi_1_dfm_4_24_22 = MUX_v_3_2_2(3'b000, Silu_for_else_Silu_for_else_mux1h_65_nl,
      Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
  assign Silu_for_else_Silu_for_else_mux1h_30_nl = MUX1HOT_s_1_4_2((Silu_for_y_8_sva_1_22_0_1[22]),
      (Silu_for_15_else_else_if_acc_itm[1]), ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_1_25,
      reg_nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0,
      {(~ Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_28_ssc_1 , Silu_for_else_else_else_and_28_ssc_1 , Silu_for_else_else_else_and_29_ssc_1});
  assign Silu_for_y_15_lpi_1_dfm_4_25 = Silu_for_else_Silu_for_else_mux1h_30_nl &
      (~ Silu_for_else_and_46_ssc_1) & Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  assign Silu_for_else_Silu_for_else_mux1h_67_nl = MUX1HOT_v_3_5_2((signext_3_1(Silu_for_y_8_sva_1_22_0_1[22])),
      ({{1{Silu_for_15_else_else_if_acc_itm[1]}}, Silu_for_15_else_else_if_acc_itm}),
      reg_Silu_for_15_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd,
      ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_1_24_22, reg_nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1,
      {(~ Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_28_ssc_1 , Silu_for_else_and_46_ssc_1 , Silu_for_else_else_else_and_28_ssc_1
      , Silu_for_else_else_else_and_29_ssc_1});
  assign Silu_for_y_15_lpi_1_dfm_4_24_22 = MUX_v_3_2_2(3'b000, Silu_for_else_Silu_for_else_mux1h_67_nl,
      Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
  assign Silu_for_else_Silu_for_else_mux1h_29_nl = MUX1HOT_s_1_4_2((Silu_for_y_7_sva_1_22_0_1[22]),
      (Silu_for_14_else_else_if_acc_itm[1]), ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_1_25,
      reg_nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0,
      {(~ Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_26_ssc_1 , Silu_for_else_else_else_and_26_ssc_1 , Silu_for_else_else_else_and_27_ssc_1});
  assign Silu_for_y_14_lpi_1_dfm_4_25 = Silu_for_else_Silu_for_else_mux1h_29_nl &
      (~ Silu_for_else_and_45_ssc_1) & Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  assign Silu_for_else_Silu_for_else_mux1h_69_nl = MUX1HOT_v_3_5_2((signext_3_1(Silu_for_y_7_sva_1_22_0_1[22])),
      ({{1{Silu_for_14_else_else_if_acc_itm[1]}}, Silu_for_14_else_else_if_acc_itm}),
      reg_Silu_for_14_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd,
      ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_1_24_22, reg_nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1,
      {(~ Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_26_ssc_1 , Silu_for_else_and_45_ssc_1 , Silu_for_else_else_else_and_26_ssc_1
      , Silu_for_else_else_else_and_27_ssc_1});
  assign Silu_for_y_14_lpi_1_dfm_4_24_22 = MUX_v_3_2_2(3'b000, Silu_for_else_Silu_for_else_mux1h_69_nl,
      Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
  assign Silu_for_else_Silu_for_else_mux1h_28_nl = MUX1HOT_s_1_4_2((Silu_for_y_6_sva_1_22_0_1[22]),
      (Silu_for_13_else_else_if_acc_itm[1]), rva_out_reg_data_39_32_sva_dfm_6_3,
      reg_nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0,
      {(~ Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_24_ssc_1 , Silu_for_else_else_else_and_24_ssc_1 , Silu_for_else_else_else_and_25_ssc_1});
  assign Silu_for_y_13_lpi_1_dfm_4_25 = Silu_for_else_Silu_for_else_mux1h_28_nl &
      (~ Silu_for_else_and_44_ssc_1) & Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  assign Silu_for_else_Silu_for_else_mux1h_71_nl = MUX1HOT_v_3_5_2((signext_3_1(Silu_for_y_6_sva_1_22_0_1[22])),
      ({{1{Silu_for_13_else_else_if_acc_itm[1]}}, Silu_for_13_else_else_if_acc_itm}),
      reg_Silu_for_13_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd,
      rva_out_reg_data_39_32_sva_dfm_6_2_0, reg_nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1,
      {(~ Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_24_ssc_1 , Silu_for_else_and_44_ssc_1 , Silu_for_else_else_else_and_24_ssc_1
      , Silu_for_else_else_else_and_25_ssc_1});
  assign Silu_for_y_13_lpi_1_dfm_4_24_22 = MUX_v_3_2_2(3'b000, Silu_for_else_Silu_for_else_mux1h_71_nl,
      Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
  assign Silu_for_else_Silu_for_else_mux1h_27_nl = MUX1HOT_s_1_4_2((Silu_for_y_5_sva_1_22_0_1[22]),
      (Silu_for_12_else_else_if_acc_itm[1]), rva_out_reg_data_29_24_sva_dfm_6_3,
      reg_nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0,
      {(~ Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_22_ssc_1 , Silu_for_else_else_else_and_22_ssc_1 , Silu_for_else_else_else_and_23_ssc_1});
  assign Silu_for_y_12_lpi_1_dfm_4_25 = Silu_for_else_Silu_for_else_mux1h_27_nl &
      (~ Silu_for_else_and_43_ssc_1) & Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  assign Silu_for_else_Silu_for_else_mux1h_73_nl = MUX1HOT_v_3_5_2((signext_3_1(Silu_for_y_5_sva_1_22_0_1[22])),
      ({{1{Silu_for_12_else_else_if_acc_itm[1]}}, Silu_for_12_else_else_if_acc_itm}),
      reg_Silu_for_12_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd,
      rva_out_reg_data_29_24_sva_dfm_6_2_0, reg_nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1,
      {(~ Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_22_ssc_1 , Silu_for_else_and_43_ssc_1 , Silu_for_else_else_else_and_22_ssc_1
      , Silu_for_else_else_else_and_23_ssc_1});
  assign Silu_for_y_12_lpi_1_dfm_4_24_22 = MUX_v_3_2_2(3'b000, Silu_for_else_Silu_for_else_mux1h_73_nl,
      Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
  assign Silu_for_else_Silu_for_else_mux1h_26_nl = MUX1HOT_s_1_4_2((Silu_for_y_4_sva_1_22_0_1[22]),
      (Silu_for_11_else_else_if_acc_itm[1]), act_config_output_counter_sva_3, reg_nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0,
      {(~ Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_20_ssc_1 , Silu_for_else_else_else_and_20_ssc_1 , Silu_for_else_else_else_and_21_ssc_1});
  assign Silu_for_y_11_lpi_1_dfm_4_25 = Silu_for_else_Silu_for_else_mux1h_26_nl &
      (~ Silu_for_else_and_42_ssc_1) & Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  assign Silu_for_else_Silu_for_else_mux1h_75_nl = MUX1HOT_v_3_5_2((signext_3_1(Silu_for_y_4_sva_1_22_0_1[22])),
      ({{1{Silu_for_11_else_else_if_acc_itm[1]}}, Silu_for_11_else_else_if_acc_itm}),
      reg_Silu_for_11_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd,
      act_config_output_counter_sva_2_0, reg_nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1,
      {(~ Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_20_ssc_1 , Silu_for_else_and_42_ssc_1 , Silu_for_else_else_else_and_20_ssc_1
      , Silu_for_else_else_else_and_21_ssc_1});
  assign Silu_for_y_11_lpi_1_dfm_4_24_22 = MUX_v_3_2_2(3'b000, Silu_for_else_Silu_for_else_mux1h_75_nl,
      Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
  assign Silu_for_else_Silu_for_else_mux1h_25_nl = MUX1HOT_s_1_4_2((Silu_for_y_3_sva_1_22_0_1[22]),
      (Silu_for_10_else_else_if_acc_itm[1]), (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[3]),
      reg_nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0,
      {(~ Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_18_ssc_1 , Silu_for_else_else_else_and_18_ssc_1 , Silu_for_else_else_else_and_19_ssc_1});
  assign Silu_for_y_10_lpi_1_dfm_4_25 = Silu_for_else_Silu_for_else_mux1h_25_nl &
      (~ Silu_for_else_and_41_ssc_1) & Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  assign Silu_for_else_Silu_for_else_mux1h_77_nl = MUX1HOT_v_3_5_2((signext_3_1(Silu_for_y_3_sva_1_22_0_1[22])),
      ({{1{Silu_for_10_else_else_if_acc_itm[1]}}, Silu_for_10_else_else_if_acc_itm}),
      reg_Silu_for_10_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd,
      (ActUnit_PushOutput_if_for_i_4_0_sva_3_0[2:0]), reg_nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1,
      {(~ Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_18_ssc_1 , Silu_for_else_and_41_ssc_1 , Silu_for_else_else_else_and_18_ssc_1
      , Silu_for_else_else_else_and_19_ssc_1});
  assign Silu_for_y_10_lpi_1_dfm_4_24_22 = MUX_v_3_2_2(3'b000, Silu_for_else_Silu_for_else_mux1h_77_nl,
      Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
  assign Silu_for_else_Silu_for_else_mux1h_24_nl = MUX1HOT_s_1_4_2((Silu_for_y_2_sva_1_22_0_1[22]),
      (Silu_for_9_else_else_if_acc_itm[1]), ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_1_25,
      reg_nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0,
      {(~ Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_16_ssc_1 , Silu_for_else_else_else_and_16_ssc_1 , Silu_for_else_else_else_and_17_ssc_1});
  assign Silu_for_y_9_lpi_1_dfm_4_25 = Silu_for_else_Silu_for_else_mux1h_24_nl &
      (~ Silu_for_else_and_40_ssc_1) & Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
  assign Silu_for_else_Silu_for_else_mux1h_79_nl = MUX1HOT_v_3_5_2((signext_3_1(Silu_for_y_2_sva_1_22_0_1[22])),
      ({{1{Silu_for_9_else_else_if_acc_itm[1]}}, Silu_for_9_else_else_if_acc_itm}),
      Silu_for_9_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_24_22,
      ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_1_24_22, reg_nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1,
      {(~ Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_16_ssc_1 , Silu_for_else_and_40_ssc_1 , Silu_for_else_else_else_and_16_ssc_1
      , Silu_for_else_else_else_and_17_ssc_1});
  assign Silu_for_y_9_lpi_1_dfm_4_24_22 = MUX_v_3_2_2(3'b000, Silu_for_else_Silu_for_else_mux1h_79_nl,
      Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_7_cse <= 1'b0;
      reg_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_6_cse <= 1'b0;
      reg_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_5_cse <= 1'b0;
      reg_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_4_cse <= 1'b0;
      reg_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_3_cse <= 1'b0;
      reg_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_2_cse <= 1'b0;
      reg_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_1_cse <= 1'b0;
      reg_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_cse <= 1'b0;
      reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_15_cse <= 1'b0;
      reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_14_cse <= 1'b0;
      reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_13_cse <= 1'b0;
      reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_12_cse <= 1'b0;
      reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_11_cse <= 1'b0;
      reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_10_cse <= 1'b0;
      reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_9_cse <= 1'b0;
      reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_8_cse <= 1'b0;
      reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_7_cse <= 1'b0;
      reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_6_cse <= 1'b0;
      reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_5_cse <= 1'b0;
      reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_4_cse <= 1'b0;
      reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_3_cse <= 1'b0;
      reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_2_cse <= 1'b0;
      reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_1_cse <= 1'b0;
      reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_cse <= 1'b0;
      reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_15_cse <= 1'b0;
      reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_14_cse <= 1'b0;
      reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_13_cse <= 1'b0;
      reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_12_cse <= 1'b0;
      reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_11_cse <= 1'b0;
      reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_10_cse <= 1'b0;
      reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_9_cse <= 1'b0;
      reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_8_cse <= 1'b0;
      reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_7_cse <= 1'b0;
      reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_6_cse <= 1'b0;
      reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_5_cse <= 1'b0;
      reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_4_cse <= 1'b0;
      reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_3_cse <= 1'b0;
      reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_2_cse <= 1'b0;
      reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_1_cse <= 1'b0;
      reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_cse <= 1'b0;
      reg_done_Push_mioi_iswt0_cse <= 1'b0;
      reg_output_port_Push_mioi_iswt0_cse <= 1'b0;
      reg_start_PopNB_mioi_iswt0_cse <= 1'b0;
      reg_rva_out_Push_mioi_iswt0_cse <= 1'b0;
      reg_act_port_PopNB_mioi_iswt0_cse <= 1'b0;
      reg_rva_in_PopNB_mioi_iswt0_cse <= 1'b0;
      ActUnit_RunInst_switch_lp_nor_tmp <= 1'b0;
      act_write_req_valid_lpi_1_dfm_5 <= 1'b0;
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen ) begin
      reg_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_7_cse <= and_899_rmff;
      reg_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_6_cse <= and_900_rmff;
      reg_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_5_cse <= and_901_rmff;
      reg_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_4_cse <= and_902_rmff;
      reg_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_3_cse <= and_903_rmff;
      reg_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_2_cse <= and_904_rmff;
      reg_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_1_cse <= and_905_rmff;
      reg_Silu_for_1_else_if_Silu_for_else_if_mul_cmp_cgo_ir_cse <= and_906_rmff;
      reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_15_cse <= and_915_rmff;
      reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_14_cse <= and_920_rmff;
      reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_13_cse <= and_925_rmff;
      reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_12_cse <= and_930_rmff;
      reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_11_cse <= and_935_rmff;
      reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_10_cse <= and_940_rmff;
      reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_9_cse <= and_945_rmff;
      reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_8_cse <= and_950_rmff;
      reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_7_cse <= and_955_rmff;
      reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_6_cse <= and_960_rmff;
      reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_5_cse <= and_965_rmff;
      reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_4_cse <= and_970_rmff;
      reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_3_cse <= and_975_rmff;
      reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_2_cse <= and_980_rmff;
      reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_1_cse <= and_985_rmff;
      reg_Gelu_for_1_else_else_if_mul_cmp_cgo_ir_cse <= and_990_rmff;
      reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_15_cse <= and_998_rmff;
      reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_14_cse <= and_1004_rmff;
      reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_13_cse <= and_1010_rmff;
      reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_12_cse <= and_1016_rmff;
      reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_11_cse <= and_1022_rmff;
      reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_10_cse <= and_1028_rmff;
      reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_9_cse <= and_1034_rmff;
      reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_8_cse <= and_1040_rmff;
      reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_7_cse <= and_1046_rmff;
      reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_6_cse <= and_1052_rmff;
      reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_5_cse <= and_1058_rmff;
      reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_4_cse <= and_1064_rmff;
      reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_3_cse <= and_1070_rmff;
      reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_2_cse <= and_1076_rmff;
      reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_1_cse <= and_1082_rmff;
      reg_Gelu_for_1_else_else_else_if_mul_cmp_cgo_ir_cse <= and_1088_rmff;
      reg_done_Push_mioi_iswt0_cse <= and_1097_rmff;
      reg_output_port_Push_mioi_iswt0_cse <= and_1102_rmff;
      reg_start_PopNB_mioi_iswt0_cse <= and_1106_rmff;
      reg_rva_out_Push_mioi_iswt0_cse <= and_1108_rmff;
      reg_act_port_PopNB_mioi_iswt0_cse <= and_1113_rmff;
      reg_rva_in_PopNB_mioi_iswt0_cse <= and_1116_rmff;
      ActUnit_RunInst_switch_lp_nor_tmp <= ActUnit_RunInst_switch_lp_nor_tmp_mx0;
      act_write_req_valid_lpi_1_dfm_5 <= MUX_s_1_2_2(ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_7_nl,
          ActUnit_RunInst_switch_lp_and_32_tmp, is_start_sva);
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_31 <= ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_31_3;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_config_is_zero_first_sva <= 1'b0;
    end
    else if ( ActUnitRun_wen & (fsm_output[3]) ) begin
      act_config_is_zero_first_sva <= MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
          while_else_1_mux_1_itm, and_1122_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva
          <= 1'b0;
      ActUnit_DecodeAxi_rva_in_reg_rw_sva <= 1'b0;
    end
    else if ( ActUnit_DecodeAxi_if_and_37_cse ) begin
      ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva
          <= ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_mx1;
      ActUnit_DecodeAxi_rva_in_reg_rw_sva <= ActUnit_DecodeAxi_rva_in_reg_rw_sva_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      is_start_sva <= 1'b0;
    end
    else if ( is_start_and_tmp ) begin
      is_start_sva <= MUX_s_1_2_2(while_else_1_while_else_1_nand_1_nl, ActUnit_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva,
          and_dcpl_1085);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_DecodeAxiRead_else_unequal_tmp <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_466 | or_dcpl_464)) ) begin
      ActUnit_DecodeAxiRead_else_unequal_tmp <= ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_DecodeAxiWrite_else_unequal_tmp <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_469 | or_dcpl_464)) ) begin
      ActUnit_DecodeAxiWrite_else_unequal_tmp <= ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_config_inst_regs_0_sva_0 <= 1'b0;
      act_config_inst_regs_16_sva_0 <= 1'b0;
      act_config_inst_regs_1_sva_0 <= 1'b0;
      act_config_inst_regs_17_sva_0 <= 1'b0;
    end
    else if ( act_config_inst_regs_and_36_cse ) begin
      act_config_inst_regs_0_sva_0 <= act_config_inst_regs_0_sva_dfm_5[0];
      act_config_inst_regs_16_sva_0 <= act_config_inst_regs_16_sva_dfm_6[0];
      act_config_inst_regs_1_sva_0 <= act_config_inst_regs_1_sva_dfm_5[0];
      act_config_inst_regs_17_sva_0 <= act_config_inst_regs_17_sva_dfm_6[0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_config_num_inst_sva <= 6'b000001;
      act_config_num_output_sva <= 8'b00000001;
      act_config_buffer_addr_base_sva <= 5'b00000;
      act_config_output_addr_base_sva <= 8'b00000000;
    end
    else if ( act_config_num_inst_and_cse ) begin
      act_config_num_inst_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[29:24];
      act_config_num_output_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[39:32];
      act_config_buffer_addr_base_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[52:48];
      act_config_output_addr_base_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[71:64];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_config_is_valid_sva <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~(act_config_ActConfigRead_unequal_tmp_1 | ActUnit_DecodeAxiRead_unequal_tmp_1
        | or_dcpl_468 | or_dcpl_462 | or_dcpl_487 | (fsm_output[3]))) ) begin
      act_config_is_valid_sva <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_29_24_sva_dfm_6_5_4 <= 2'b00;
    end
    else if ( rva_out_reg_data_and_ssc ) begin
      rva_out_reg_data_29_24_sva_dfm_6_5_4 <= MUX_v_2_2_2((act_mem_banks_read_read_data_lpi_1_dfm_1_31_0[29:28]),
          rva_out_reg_data_29_24_sva_dfm_3_5_4, and_dcpl_1096);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_39_32_sva_dfm_6_7_4 <= 4'b0000;
    end
    else if ( ActUnitRun_wen & (rva_out_reg_data_39_32_sva_dfm_6_mx0c0 | and_dcpl_1094
        | and_dcpl_1096) ) begin
      rva_out_reg_data_39_32_sva_dfm_6_7_4 <= MUX_v_4_2_2((act_mem_banks_read_read_data_lpi_1_dfm_1_63_32[7:4]),
          rva_out_reg_data_39_32_sva_dfm_3_7_4, and_dcpl_1096);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_71_64_sva_dfm_6_7_5 <= 3'b000;
    end
    else if ( ActUnitRun_wen & (not_tmp_495 | and_dcpl_1094 | and_dcpl_1096) ) begin
      rva_out_reg_data_71_64_sva_dfm_6_7_5 <= MUX_v_3_2_2((act_mem_banks_read_read_data_lpi_1_dfm_1_95_64[7:5]),
          rva_out_reg_data_71_64_sva_dfm_3_7_5, and_dcpl_1096);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_71_64_sva_dfm_6_4_0 <= 5'b00000;
    end
    else if ( and_1803_tmp ) begin
      rva_out_reg_data_71_64_sva_dfm_6_4_0 <= MUX1HOT_v_5_3_2(and_1716_nl, (act_mem_banks_read_read_data_lpi_1_dfm_1_95_64[4:0]),
          rva_out_reg_data_71_64_sva_dfm_3_4_0, {not_tmp_495 , and_dcpl_1094 , and_dcpl_1096});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_0_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_0_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_0_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_0_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_0_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_0_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_0_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_0_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_0_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_0_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_0_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_0_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_0_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_0_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_0_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_0_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_cse ) begin
      act_mem_banks_bank_a_0_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_0_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_0_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_0_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_0_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_0_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_0_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_0_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_0_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_0_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_0_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_0_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_0_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_0_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_0_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_0_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_1_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_1_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_1_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_1_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_1_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_1_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_1_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_1_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_1_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_1_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_1_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_1_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_1_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_1_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_1_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_1_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_1_cse ) begin
      act_mem_banks_bank_a_1_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_1_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_1_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_1_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_1_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_1_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_1_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_1_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_1_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_1_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_1_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_1_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_1_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_1_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_1_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_1_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_2_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_2_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_2_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_2_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_2_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_2_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_2_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_2_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_2_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_2_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_2_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_2_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_2_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_2_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_2_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_2_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_2_cse ) begin
      act_mem_banks_bank_a_2_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_2_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_2_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_2_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_2_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_2_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_2_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_2_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_2_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_2_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_2_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_2_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_2_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_2_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_2_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_2_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_3_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_3_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_3_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_3_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_3_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_3_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_3_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_3_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_3_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_3_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_3_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_3_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_3_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_3_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_3_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_3_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_3_cse ) begin
      act_mem_banks_bank_a_3_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_3_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_3_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_3_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_3_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_3_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_3_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_3_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_3_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_3_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_3_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_3_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_3_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_3_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_3_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_3_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_4_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_4_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_4_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_4_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_4_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_4_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_4_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_4_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_4_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_4_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_4_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_4_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_4_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_4_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_4_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_4_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_4_cse ) begin
      act_mem_banks_bank_a_4_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_4_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_4_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_4_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_4_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_4_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_4_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_4_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_4_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_4_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_4_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_4_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_4_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_4_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_4_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_4_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_5_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_5_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_5_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_5_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_5_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_5_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_5_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_5_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_5_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_5_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_5_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_5_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_5_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_5_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_5_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_5_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_5_cse ) begin
      act_mem_banks_bank_a_5_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_5_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_5_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_5_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_5_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_5_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_5_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_5_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_5_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_5_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_5_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_5_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_5_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_5_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_5_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_5_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_6_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_6_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_6_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_6_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_6_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_6_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_6_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_6_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_6_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_6_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_6_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_6_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_6_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_6_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_6_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_6_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_6_cse ) begin
      act_mem_banks_bank_a_6_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_6_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_6_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_6_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_6_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_6_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_6_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_6_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_6_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_6_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_6_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_6_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_6_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_6_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_6_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_6_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_7_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_7_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_7_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_7_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_7_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_7_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_7_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_7_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_7_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_7_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_7_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_7_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_7_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_7_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_7_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_7_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_7_cse ) begin
      act_mem_banks_bank_a_7_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_7_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_7_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_7_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_7_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_7_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_7_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_7_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_7_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_7_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_7_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_7_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_7_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_7_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_7_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_7_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_8_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_8_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_8_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_8_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_8_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_8_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_8_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_8_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_8_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_8_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_8_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_8_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_8_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_8_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_8_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_8_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_8_cse ) begin
      act_mem_banks_bank_a_8_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_8_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_8_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_8_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_8_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_8_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_8_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_8_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_8_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_8_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_8_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_8_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_8_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_8_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_8_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_8_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_9_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_9_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_9_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_9_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_9_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_9_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_9_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_9_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_9_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_9_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_9_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_9_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_9_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_9_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_9_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_9_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_9_cse ) begin
      act_mem_banks_bank_a_9_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_9_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_9_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_9_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_9_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_9_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_9_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_9_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_9_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_9_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_9_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_9_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_9_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_9_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_9_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_9_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_10_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_10_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_10_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_10_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_10_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_10_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_10_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_10_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_10_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_10_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_10_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_10_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_10_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_10_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_10_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_10_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_10_cse ) begin
      act_mem_banks_bank_a_10_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_10_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_10_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_10_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_10_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_10_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_10_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_10_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_10_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_10_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_10_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_10_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_10_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_10_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_10_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_10_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_11_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_11_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_11_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_11_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_11_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_11_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_11_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_11_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_11_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_11_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_11_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_11_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_11_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_11_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_11_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_11_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_11_cse ) begin
      act_mem_banks_bank_a_11_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_11_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_11_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_11_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_11_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_11_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_11_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_11_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_11_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_11_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_11_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_11_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_11_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_11_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_11_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_11_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_12_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_12_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_12_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_12_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_12_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_12_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_12_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_12_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_12_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_12_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_12_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_12_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_12_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_12_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_12_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_12_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_12_cse ) begin
      act_mem_banks_bank_a_12_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_12_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_12_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_12_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_12_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_12_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_12_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_12_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_12_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_12_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_12_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_12_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_12_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_12_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_12_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_12_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_13_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_13_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_13_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_13_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_13_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_13_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_13_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_13_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_13_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_13_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_13_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_13_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_13_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_13_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_13_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_13_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_13_cse ) begin
      act_mem_banks_bank_a_13_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_13_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_13_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_13_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_13_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_13_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_13_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_13_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_13_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_13_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_13_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_13_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_13_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_13_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_13_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_13_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_14_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_14_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_14_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_14_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_14_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_14_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_14_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_14_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_14_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_14_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_14_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_14_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_14_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_14_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_14_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_14_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_14_cse ) begin
      act_mem_banks_bank_a_14_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_14_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_14_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_14_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_14_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_14_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_14_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_14_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_14_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_14_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_14_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_14_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_14_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_14_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_14_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_14_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_15_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_15_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_15_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_15_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_15_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_15_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_15_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_15_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_15_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_15_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_15_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_15_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_15_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_15_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_15_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_15_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_15_cse ) begin
      act_mem_banks_bank_a_15_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_15_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_15_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_15_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_15_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_15_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_15_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_15_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_15_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_15_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_15_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_15_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_15_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_15_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_15_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_15_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_16_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_16_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_16_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_16_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_16_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_16_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_16_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_16_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_16_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_16_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_16_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_16_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_16_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_16_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_16_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_16_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_16_cse ) begin
      act_mem_banks_bank_a_16_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_16_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_16_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_16_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_16_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_16_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_16_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_16_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_16_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_16_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_16_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_16_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_16_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_16_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_16_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_16_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_17_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_17_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_17_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_17_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_17_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_17_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_17_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_17_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_17_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_17_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_17_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_17_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_17_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_17_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_17_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_17_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_17_cse ) begin
      act_mem_banks_bank_a_17_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_17_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_17_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_17_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_17_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_17_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_17_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_17_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_17_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_17_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_17_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_17_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_17_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_17_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_17_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_17_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_18_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_18_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_18_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_18_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_18_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_18_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_18_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_18_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_18_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_18_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_18_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_18_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_18_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_18_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_18_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_18_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_18_cse ) begin
      act_mem_banks_bank_a_18_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_18_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_18_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_18_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_18_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_18_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_18_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_18_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_18_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_18_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_18_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_18_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_18_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_18_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_18_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_18_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_19_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_19_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_19_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_19_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_19_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_19_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_19_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_19_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_19_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_19_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_19_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_19_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_19_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_19_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_19_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_19_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_19_cse ) begin
      act_mem_banks_bank_a_19_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_19_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_19_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_19_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_19_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_19_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_19_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_19_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_19_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_19_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_19_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_19_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_19_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_19_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_19_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_19_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_20_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_20_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_20_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_20_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_20_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_20_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_20_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_20_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_20_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_20_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_20_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_20_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_20_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_20_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_20_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_20_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_20_cse ) begin
      act_mem_banks_bank_a_20_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_20_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_20_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_20_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_20_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_20_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_20_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_20_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_20_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_20_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_20_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_20_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_20_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_20_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_20_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_20_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_21_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_21_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_21_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_21_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_21_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_21_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_21_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_21_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_21_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_21_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_21_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_21_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_21_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_21_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_21_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_21_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_21_cse ) begin
      act_mem_banks_bank_a_21_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_21_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_21_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_21_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_21_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_21_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_21_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_21_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_21_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_21_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_21_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_21_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_21_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_21_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_21_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_21_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_22_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_22_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_22_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_22_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_22_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_22_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_22_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_22_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_22_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_22_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_22_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_22_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_22_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_22_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_22_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_22_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_22_cse ) begin
      act_mem_banks_bank_a_22_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_22_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_22_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_22_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_22_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_22_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_22_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_22_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_22_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_22_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_22_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_22_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_22_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_22_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_22_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_22_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_23_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_23_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_23_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_23_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_23_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_23_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_23_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_23_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_23_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_23_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_23_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_23_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_23_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_23_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_23_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_23_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_23_cse ) begin
      act_mem_banks_bank_a_23_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_23_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_23_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_23_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_23_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_23_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_23_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_23_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_23_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_23_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_23_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_23_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_23_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_23_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_23_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_23_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_24_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_24_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_24_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_24_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_24_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_24_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_24_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_24_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_24_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_24_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_24_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_24_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_24_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_24_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_24_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_24_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_24_cse ) begin
      act_mem_banks_bank_a_24_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_24_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_24_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_24_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_24_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_24_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_24_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_24_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_24_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_24_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_24_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_24_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_24_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_24_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_24_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_24_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_25_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_25_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_25_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_25_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_25_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_25_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_25_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_25_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_25_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_25_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_25_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_25_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_25_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_25_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_25_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_25_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_25_cse ) begin
      act_mem_banks_bank_a_25_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_25_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_25_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_25_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_25_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_25_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_25_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_25_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_25_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_25_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_25_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_25_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_25_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_25_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_25_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_25_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_26_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_26_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_26_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_26_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_26_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_26_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_26_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_26_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_26_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_26_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_26_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_26_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_26_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_26_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_26_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_26_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_26_cse ) begin
      act_mem_banks_bank_a_26_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_26_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_26_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_26_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_26_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_26_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_26_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_26_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_26_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_26_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_26_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_26_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_26_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_26_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_26_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_26_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_27_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_27_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_27_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_27_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_27_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_27_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_27_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_27_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_27_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_27_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_27_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_27_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_27_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_27_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_27_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_27_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_27_cse ) begin
      act_mem_banks_bank_a_27_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_27_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_27_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_27_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_27_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_27_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_27_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_27_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_27_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_27_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_27_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_27_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_27_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_27_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_27_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_27_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_28_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_28_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_28_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_28_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_28_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_28_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_28_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_28_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_28_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_28_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_28_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_28_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_28_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_28_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_28_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_28_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_28_cse ) begin
      act_mem_banks_bank_a_28_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_28_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_28_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_28_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_28_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_28_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_28_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_28_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_28_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_28_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_28_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_28_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_28_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_28_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_28_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_28_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_29_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_29_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_29_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_29_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_29_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_29_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_29_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_29_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_29_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_29_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_29_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_29_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_29_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_29_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_29_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_29_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_29_cse ) begin
      act_mem_banks_bank_a_29_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_29_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_29_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_29_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_29_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_29_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_29_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_29_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_29_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_29_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_29_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_29_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_29_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_29_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_29_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_29_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_30_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_30_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_30_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_30_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_30_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_30_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_30_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_30_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_30_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_30_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_30_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_30_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_30_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_30_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_30_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_30_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_30_cse ) begin
      act_mem_banks_bank_a_30_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_30_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_30_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_30_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_30_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_30_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_30_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_30_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_30_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_30_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_30_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_30_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_30_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_30_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_30_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_30_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_bank_a_31_31_0_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_31_63_32_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_31_95_64_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_31_127_96_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_31_159_128_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_31_191_160_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_31_223_192_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_31_255_224_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_31_287_256_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_31_319_288_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_31_351_320_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_31_383_352_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_31_415_384_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_31_447_416_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_31_479_448_sva_dfm <= 32'b00000000000000000000000000000000;
      act_mem_banks_bank_a_31_511_480_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_bank_a_and_31_cse ) begin
      act_mem_banks_bank_a_31_31_0_sva_dfm <= act_write_data_data_0_0_lpi_1_dfm_7;
      act_mem_banks_bank_a_31_63_32_sva_dfm <= act_write_data_data_0_1_lpi_1_dfm_7;
      act_mem_banks_bank_a_31_95_64_sva_dfm <= act_write_data_data_0_2_lpi_1_dfm_7;
      act_mem_banks_bank_a_31_127_96_sva_dfm <= act_write_data_data_0_3_lpi_1_dfm_7;
      act_mem_banks_bank_a_31_159_128_sva_dfm <= act_write_data_data_0_4_lpi_1_dfm_7;
      act_mem_banks_bank_a_31_191_160_sva_dfm <= act_write_data_data_0_5_lpi_1_dfm_7;
      act_mem_banks_bank_a_31_223_192_sva_dfm <= act_write_data_data_0_6_lpi_1_dfm_7;
      act_mem_banks_bank_a_31_255_224_sva_dfm <= act_write_data_data_0_7_lpi_1_dfm_7;
      act_mem_banks_bank_a_31_287_256_sva_dfm <= act_write_data_data_0_8_lpi_1_dfm_7;
      act_mem_banks_bank_a_31_319_288_sva_dfm <= act_write_data_data_0_9_lpi_1_dfm_7;
      act_mem_banks_bank_a_31_351_320_sva_dfm <= act_write_data_data_0_10_lpi_1_dfm_7;
      act_mem_banks_bank_a_31_383_352_sva_dfm <= act_write_data_data_0_11_lpi_1_dfm_7;
      act_mem_banks_bank_a_31_415_384_sva_dfm <= act_write_data_data_0_12_lpi_1_dfm_7;
      act_mem_banks_bank_a_31_447_416_sva_dfm <= act_write_data_data_0_13_lpi_1_dfm_7;
      act_mem_banks_bank_a_31_479_448_sva_dfm <= act_write_data_data_0_14_lpi_1_dfm_7;
      act_mem_banks_bank_a_31_511_480_sva_dfm <= act_write_data_data_0_15_lpi_1_dfm_7;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_config_inst_regs_16_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_17_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_18_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_19_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_20_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_21_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_22_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_23_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_24_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_25_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_26_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_27_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_28_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_29_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_30_sva_dfm_6 <= 8'b00000000;
      act_config_inst_regs_31_sva_dfm_6 <= 8'b00000000;
    end
    else if ( act_config_inst_regs_and_4_cse ) begin
      act_config_inst_regs_16_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[7:0];
      act_config_inst_regs_17_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[15:8];
      act_config_inst_regs_18_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[23:16];
      act_config_inst_regs_19_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[31:24];
      act_config_inst_regs_20_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[39:32];
      act_config_inst_regs_21_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[47:40];
      act_config_inst_regs_22_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[55:48];
      act_config_inst_regs_23_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[63:56];
      act_config_inst_regs_24_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[71:64];
      act_config_inst_regs_25_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[79:72];
      act_config_inst_regs_26_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[87:80];
      act_config_inst_regs_27_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[95:88];
      act_config_inst_regs_28_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[103:96];
      act_config_inst_regs_29_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[111:104];
      act_config_inst_regs_30_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[119:112];
      act_config_inst_regs_31_sva_dfm_6 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[127:120];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_config_inst_regs_0_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_1_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_2_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_3_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_4_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_5_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_6_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_7_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_8_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_9_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_10_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_11_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_12_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_13_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_14_sva_dfm_5 <= 8'b00000000;
      act_config_inst_regs_15_sva_dfm_5 <= 8'b00000000;
    end
    else if ( act_config_inst_regs_and_20_cse ) begin
      act_config_inst_regs_0_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[7:0];
      act_config_inst_regs_1_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[15:8];
      act_config_inst_regs_2_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[23:16];
      act_config_inst_regs_3_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[31:24];
      act_config_inst_regs_4_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[39:32];
      act_config_inst_regs_5_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[47:40];
      act_config_inst_regs_6_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[55:48];
      act_config_inst_regs_7_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[63:56];
      act_config_inst_regs_8_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[71:64];
      act_config_inst_regs_9_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[79:72];
      act_config_inst_regs_10_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[87:80];
      act_config_inst_regs_11_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[95:88];
      act_config_inst_regs_12_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[103:96];
      act_config_inst_regs_13_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[111:104];
      act_config_inst_regs_14_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[119:112];
      act_config_inst_regs_15_sva_dfm_5 <= rva_in_PopNB_mioi_data_data_rsc_z_mxwt[127:120];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_config_output_counter_sva_7_4 <= 4'b0000;
    end
    else if ( act_config_output_counter_and_ssc ) begin
      act_config_output_counter_sva_7_4 <= MUX_v_4_2_2(act_config_InstIncr_if_act_config_InstIncr_if_and_1_nl,
          reg_act_config_output_counter_sva_dfm_3_ftd, act_config_output_counter_sva_mx0c2);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_config_output_counter_sva_3 <= 1'b0;
      act_config_output_counter_sva_2_0 <= 3'b000;
    end
    else if ( act_config_output_counter_and_2_ssc ) begin
      act_config_output_counter_sva_3 <= MUX1HOT_s_1_4_2((Silu_for_11_else_else_else_else_if_acc_sdt[3]),
          ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_25_22_mx0w2_3,
          act_config_InstIncr_if_act_config_InstIncr_if_and_2_nl, reg_act_config_output_counter_sva_dfm_3_ftd_1_3,
          {act_config_output_counter_and_3_ssc , and_dcpl_1235 , act_config_output_counter_sva_mx0c1
          , act_config_output_counter_sva_mx0c2});
      act_config_output_counter_sva_2_0 <= MUX1HOT_v_3_4_2((Silu_for_11_else_else_else_else_if_acc_sdt[2:0]),
          ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_25_22_mx0w2_2_0,
          act_config_InstIncr_if_act_config_InstIncr_if_and_3_nl, reg_act_config_output_counter_sva_dfm_3_ftd_1_2_0,
          {act_config_output_counter_and_3_ssc , and_dcpl_1235 , act_config_output_counter_sva_mx0c1
          , act_config_output_counter_sva_mx0c2});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_config_inst_counter_sva <= 5'b00000;
    end
    else if ( act_config_inst_counter_and_tmp ) begin
      act_config_inst_counter_sva <= MUX_v_5_2_2(act_config_InstIncr_act_config_InstIncr_and_1_nl,
          act_config_inst_counter_sva_dfm_3, act_config_inst_counter_sva_mx0c1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_15_sva_31 <= 1'b0;
      act_regs_data_3_14_sva_31 <= 1'b0;
      act_regs_data_3_13_sva_31 <= 1'b0;
      act_regs_data_3_12_sva_31 <= 1'b0;
      act_regs_data_3_11_sva_31 <= 1'b0;
      act_regs_data_3_10_sva_31 <= 1'b0;
      act_regs_data_3_9_sva_31 <= 1'b0;
      act_regs_data_3_8_sva_31 <= 1'b0;
      act_regs_data_3_7_sva_31 <= 1'b0;
      act_regs_data_3_6_sva_31 <= 1'b0;
      act_regs_data_3_5_sva_31 <= 1'b0;
      act_regs_data_3_4_sva_31 <= 1'b0;
      act_regs_data_3_3_sva_31 <= 1'b0;
      act_regs_data_3_2_sva_31 <= 1'b0;
      act_regs_data_3_1_sva_31 <= 1'b0;
      act_regs_data_3_0_sva_31 <= 1'b0;
      act_regs_data_2_15_sva_31 <= 1'b0;
      act_regs_data_2_14_sva_31 <= 1'b0;
      act_regs_data_2_13_sva_31 <= 1'b0;
      act_regs_data_2_12_sva_31 <= 1'b0;
      act_regs_data_2_11_sva_31 <= 1'b0;
      act_regs_data_2_10_sva_31 <= 1'b0;
      act_regs_data_2_9_sva_31 <= 1'b0;
      act_regs_data_2_8_sva_31 <= 1'b0;
      act_regs_data_2_7_sva_31 <= 1'b0;
      act_regs_data_2_6_sva_31 <= 1'b0;
      act_regs_data_2_5_sva_31 <= 1'b0;
      act_regs_data_2_4_sva_31 <= 1'b0;
      act_regs_data_2_3_sva_31 <= 1'b0;
      act_regs_data_2_2_sva_31 <= 1'b0;
      act_regs_data_2_1_sva_31 <= 1'b0;
      act_regs_data_2_0_sva_31 <= 1'b0;
      act_regs_data_1_15_sva_31 <= 1'b0;
      act_regs_data_1_14_sva_31 <= 1'b0;
      act_regs_data_1_13_sva_31 <= 1'b0;
      act_regs_data_1_12_sva_31 <= 1'b0;
      act_regs_data_1_11_sva_31 <= 1'b0;
      act_regs_data_1_10_sva_31 <= 1'b0;
      act_regs_data_1_9_sva_31 <= 1'b0;
      act_regs_data_1_8_sva_31 <= 1'b0;
      act_regs_data_1_7_sva_31 <= 1'b0;
      act_regs_data_1_6_sva_31 <= 1'b0;
      act_regs_data_1_5_sva_31 <= 1'b0;
      act_regs_data_1_4_sva_31 <= 1'b0;
      act_regs_data_1_3_sva_31 <= 1'b0;
      act_regs_data_1_2_sva_31 <= 1'b0;
      act_regs_data_1_1_sva_31 <= 1'b0;
      act_regs_data_1_0_sva_31 <= 1'b0;
      act_regs_data_0_15_sva_31 <= 1'b0;
      act_regs_data_0_14_sva_31 <= 1'b0;
      act_regs_data_0_9_sva_31 <= 1'b0;
      act_regs_data_0_8_sva_31 <= 1'b0;
      act_regs_data_0_7_sva_31 <= 1'b0;
      act_regs_data_0_6_sva_31 <= 1'b0;
      act_regs_data_0_5_sva_31 <= 1'b0;
      act_regs_data_0_4_sva_31 <= 1'b0;
      act_regs_data_0_3_sva_31 <= 1'b0;
      act_regs_data_0_2_sva_31 <= 1'b0;
      reg_act_regs_data_0_13_ftd <= 1'b0;
      reg_act_regs_data_0_12_ftd <= 1'b0;
      reg_act_regs_data_0_11_ftd <= 1'b0;
      reg_act_regs_data_0_10_ftd <= 1'b0;
      reg_act_regs_data_0_1_ftd <= 1'b0;
      reg_act_regs_data_0_0_ftd <= 1'b0;
    end
    else if ( act_regs_data_and_ssc ) begin
      act_regs_data_3_15_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_3_15_sva_dfm_2_31,
          act_regs_data_2_2_sva_8_31, act_regs_data_3_15_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_3_14_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_3_14_sva_dfm_2_31,
          act_regs_data_2_15_sva_8_31, act_regs_data_3_14_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_3_13_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_3_13_sva_dfm_2_31,
          act_regs_data_2_14_sva_8_31, act_regs_data_3_13_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_3_12_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_3_12_sva_dfm_2_31,
          act_regs_data_2_13_sva_8_31, act_regs_data_3_12_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_3_11_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_3_11_sva_dfm_2_31,
          act_regs_data_2_12_sva_8_31, act_regs_data_3_11_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_3_10_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_3_10_sva_dfm_2_31,
          act_regs_data_2_11_sva_8_31, act_regs_data_3_10_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_3_9_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_3_9_sva_dfm_2_31,
          act_regs_data_3_0_sva_8_31, act_regs_data_3_9_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_3_8_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_3_8_sva_dfm_2_31,
          act_regs_data_2_9_sva_8_31, act_regs_data_3_8_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_3_7_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_3_7_sva_dfm_2_31,
          act_regs_data_2_8_sva_8_31, act_regs_data_3_7_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_3_6_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_3_6_sva_dfm_2_31,
          act_regs_data_2_7_sva_8_31, act_regs_data_3_6_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_3_5_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_3_5_sva_dfm_2_31,
          act_regs_data_2_6_sva_8_31, act_regs_data_3_5_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_3_4_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_3_4_sva_dfm_2_31,
          act_regs_data_2_5_sva_8_31, act_regs_data_3_4_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_3_3_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_3_3_sva_dfm_2_31,
          act_regs_data_2_4_sva_8_31, act_regs_data_3_3_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_3_2_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_3_2_sva_dfm_2_31,
          act_regs_data_2_3_sva_8_31, act_regs_data_3_2_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_3_1_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_3_1_sva_dfm_2_31,
          act_regs_data_2_10_sva_8_31, act_regs_data_3_1_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_3_0_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_3_0_sva_dfm_2_31,
          act_regs_data_2_1_sva_8_31, act_regs_data_3_0_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_2_15_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_2_15_sva_dfm_2_31,
          act_regs_data_1_2_sva_8_31, act_regs_data_2_15_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_2_14_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_2_14_sva_dfm_2_31,
          act_regs_data_1_15_sva_8_31, act_regs_data_2_14_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_2_13_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_2_13_sva_dfm_2_31,
          act_regs_data_1_14_sva_8_31, act_regs_data_2_13_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_2_12_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_2_12_sva_dfm_2_31,
          act_regs_data_1_13_sva_8_31, act_regs_data_2_12_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_2_11_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_2_11_sva_dfm_2_31,
          act_regs_data_1_12_sva_8_31, act_regs_data_2_11_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_2_10_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_2_10_sva_dfm_2_31,
          act_regs_data_1_11_sva_8_31, act_regs_data_2_10_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_2_9_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_2_9_sva_dfm_2_31,
          act_regs_data_2_0_sva_8_31, act_regs_data_2_9_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_2_8_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_2_8_sva_dfm_2_31,
          act_regs_data_1_9_sva_8_31, act_regs_data_2_8_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_2_7_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_2_7_sva_dfm_2_31,
          act_regs_data_1_8_sva_8_31, act_regs_data_2_7_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_2_6_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_2_6_sva_dfm_2_31,
          act_regs_data_1_7_sva_8_31, act_regs_data_2_6_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_2_5_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_2_5_sva_dfm_2_31,
          act_regs_data_1_6_sva_8_31, act_regs_data_2_5_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_2_4_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_2_4_sva_dfm_2_31,
          act_regs_data_1_5_sva_8_31, act_regs_data_2_4_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_2_3_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_2_3_sva_dfm_2_31,
          act_regs_data_1_4_sva_8_31, act_regs_data_2_3_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_2_2_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_2_2_sva_dfm_2_31,
          act_regs_data_1_3_sva_8_31, act_regs_data_2_2_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_2_1_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_2_1_sva_dfm_2_31,
          act_regs_data_1_10_sva_8_31, act_regs_data_2_1_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_2_0_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_2_0_sva_dfm_2_31,
          act_regs_data_1_1_sva_8_31, act_regs_data_2_0_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_1_15_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_1_15_sva_dfm_2_31,
          act_regs_data_0_2_sva_8_31, act_regs_data_1_15_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_1_14_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_1_14_sva_dfm_2_31,
          act_regs_data_0_15_sva_8_31, act_regs_data_1_14_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_1_13_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_1_13_sva_dfm_2_31,
          act_regs_data_0_14_sva_8_31, act_regs_data_1_13_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_1_12_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_1_12_sva_dfm_2_31,
          act_regs_data_0_13_sva_8_31, act_regs_data_1_12_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_1_11_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_1_11_sva_dfm_2_31,
          act_regs_data_0_12_sva_8_31, act_regs_data_1_11_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_1_10_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_1_10_sva_dfm_2_31,
          act_regs_data_0_11_sva_8_31, act_regs_data_1_10_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_1_9_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_1_9_sva_dfm_2_31,
          act_regs_data_1_0_sva_8_31, act_regs_data_1_9_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_1_8_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_1_8_sva_dfm_2_31,
          act_regs_data_0_9_sva_8_31, act_regs_data_1_8_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_1_7_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_1_7_sva_dfm_2_31,
          act_regs_data_0_8_sva_8_31, act_regs_data_1_7_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_1_6_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_1_6_sva_dfm_2_31,
          act_regs_data_0_7_sva_8_31, act_regs_data_1_6_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_1_5_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_1_5_sva_dfm_2_31,
          act_regs_data_0_6_sva_8_31, act_regs_data_1_5_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_1_4_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_1_4_sva_dfm_2_31,
          act_regs_data_0_5_sva_8_31, act_regs_data_1_4_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_1_3_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_1_3_sva_dfm_2_31,
          act_regs_data_0_4_sva_8_31, act_regs_data_1_3_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_1_2_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_1_2_sva_dfm_2_31,
          act_regs_data_0_3_sva_8_31, act_regs_data_1_2_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_1_1_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_1_1_sva_dfm_2_31,
          act_regs_data_0_10_sva_8_31, act_regs_data_1_1_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_1_0_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_1_0_sva_dfm_2_31,
          act_regs_data_0_1_sva_8_31, act_regs_data_1_0_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_0_15_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_0_15_sva_dfm_2_31,
          ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_1_31, act_regs_data_0_15_sva_8_31,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_0_14_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_0_14_sva_dfm_2_31,
          ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_1_31, act_regs_data_0_14_sva_8_31,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_0_9_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_0_9_sva_dfm_2_31,
          act_regs_data_0_0_sva_8_31, act_regs_data_0_9_sva_8_31, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_0_8_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_0_8_sva_dfm_2_31,
          ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_1_31, act_regs_data_0_8_sva_8_31,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_0_7_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_0_7_sva_dfm_2_31,
          ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_1_31, act_regs_data_0_7_sva_8_31,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_0_6_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_0_6_sva_dfm_2_31,
          ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_1_31, act_regs_data_0_6_sva_8_31,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_0_5_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_0_5_sva_dfm_2_31,
          ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_1_31, act_regs_data_0_5_sva_8_31,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_0_4_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_0_4_sva_dfm_2_31,
          ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_1_31, act_regs_data_0_4_sva_8_31,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_0_3_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_0_3_sva_dfm_2_31,
          ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_1_31, act_regs_data_0_3_sva_8_31,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_0_2_sva_31 <= MUX1HOT_s_1_3_2(act_regs_data_0_2_sva_dfm_2_31,
          ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_1_31, act_regs_data_0_2_sva_8_31,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      reg_act_regs_data_0_13_ftd <= MUX1HOT_s_1_3_2(act_regs_data_0_13_sva_dfm_2_31,
          ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_1_31, act_regs_data_0_13_sva_8_31,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      reg_act_regs_data_0_12_ftd <= MUX1HOT_s_1_3_2(act_regs_data_0_12_sva_dfm_2_31,
          ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_1_31, act_regs_data_0_12_sva_8_31,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      reg_act_regs_data_0_11_ftd <= MUX1HOT_s_1_3_2(act_regs_data_0_11_sva_dfm_2_31,
          ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_1_31, act_regs_data_0_11_sva_8_31,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      reg_act_regs_data_0_10_ftd <= MUX1HOT_s_1_3_2(act_regs_data_0_10_sva_dfm_2_31,
          ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_1_31, act_regs_data_0_10_sva_8_31,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      reg_act_regs_data_0_1_ftd <= MUX1HOT_s_1_3_2(act_regs_data_0_1_sva_dfm_2_31,
          ActUnit_PushOutput_if_output_port_reg_data_data_1_sva_1_31, act_regs_data_0_1_sva_8_31,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      reg_act_regs_data_0_0_ftd <= MUX1HOT_s_1_3_2(act_regs_data_0_0_sva_dfm_2_31,
          ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_1_31, act_regs_data_0_0_sva_8_31,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_15_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2530_enex5 ) begin
      act_regs_data_3_15_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_3_15_sva_dfm_2_30_26,
          act_regs_data_2_2_sva_8_30_26, act_regs_data_3_15_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_15_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2532_enex5 ) begin
      act_regs_data_3_15_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_3_15_sva_dfm_2_21_0,
          act_regs_data_2_2_sva_8_21_0, act_regs_data_3_15_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_14_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2533_enex5 ) begin
      act_regs_data_3_14_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_3_14_sva_dfm_2_30_26,
          act_regs_data_2_15_sva_8_30_26, act_regs_data_3_14_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_14_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2535_enex5 ) begin
      act_regs_data_3_14_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_3_14_sva_dfm_2_21_0,
          act_regs_data_2_15_sva_8_21_0, act_regs_data_3_14_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_13_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2536_enex5 ) begin
      act_regs_data_3_13_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_3_13_sva_dfm_2_30_26,
          act_regs_data_2_14_sva_8_30_26, act_regs_data_3_13_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_13_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2538_enex5 ) begin
      act_regs_data_3_13_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_3_13_sva_dfm_2_21_0,
          act_regs_data_2_14_sva_8_21_0, act_regs_data_3_13_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_12_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2539_enex5 ) begin
      act_regs_data_3_12_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_3_12_sva_dfm_2_30_26,
          act_regs_data_2_13_sva_8_30_26, act_regs_data_3_12_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_12_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2541_enex5 ) begin
      act_regs_data_3_12_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_3_12_sva_dfm_2_21_0,
          act_regs_data_2_13_sva_8_21_0, act_regs_data_3_12_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_11_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2542_enex5 ) begin
      act_regs_data_3_11_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_3_11_sva_dfm_2_30_26,
          act_regs_data_2_12_sva_8_30_26, act_regs_data_3_11_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_11_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2544_enex5 ) begin
      act_regs_data_3_11_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_3_11_sva_dfm_2_21_0,
          act_regs_data_2_12_sva_8_21_0, act_regs_data_3_11_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_10_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2545_enex5 ) begin
      act_regs_data_3_10_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_3_10_sva_dfm_2_30_26,
          act_regs_data_2_11_sva_8_30_26, act_regs_data_3_10_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_10_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2547_enex5 ) begin
      act_regs_data_3_10_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_3_10_sva_dfm_2_21_0,
          act_regs_data_2_11_sva_8_21_0, act_regs_data_3_10_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_9_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2548_enex5 ) begin
      act_regs_data_3_9_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_3_9_sva_dfm_2_30_26,
          act_regs_data_3_0_sva_8_30_26, act_regs_data_3_9_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_9_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2550_enex5 ) begin
      act_regs_data_3_9_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_3_9_sva_dfm_2_21_0,
          act_regs_data_3_0_sva_8_21_0, act_regs_data_3_9_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_8_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2551_enex5 ) begin
      act_regs_data_3_8_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_3_8_sva_dfm_2_30_26,
          act_regs_data_2_9_sva_8_30_26, act_regs_data_3_8_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_8_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2553_enex5 ) begin
      act_regs_data_3_8_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_3_8_sva_dfm_2_21_0,
          act_regs_data_2_9_sva_8_21_0, act_regs_data_3_8_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_7_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2554_enex5 ) begin
      act_regs_data_3_7_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_3_7_sva_dfm_2_30_26,
          act_regs_data_2_8_sva_8_30_26, act_regs_data_3_7_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_7_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2556_enex5 ) begin
      act_regs_data_3_7_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_3_7_sva_dfm_2_21_0,
          act_regs_data_2_8_sva_8_21_0, act_regs_data_3_7_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_6_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2557_enex5 ) begin
      act_regs_data_3_6_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_3_6_sva_dfm_2_30_26,
          act_regs_data_2_7_sva_8_30_26, act_regs_data_3_6_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_6_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2559_enex5 ) begin
      act_regs_data_3_6_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_3_6_sva_dfm_2_21_0,
          act_regs_data_2_7_sva_8_21_0, act_regs_data_3_6_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_5_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2560_enex5 ) begin
      act_regs_data_3_5_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_3_5_sva_dfm_2_30_26,
          act_regs_data_2_6_sva_8_30_26, act_regs_data_3_5_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_5_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2562_enex5 ) begin
      act_regs_data_3_5_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_3_5_sva_dfm_2_21_0,
          act_regs_data_2_6_sva_8_21_0, act_regs_data_3_5_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_4_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2563_enex5 ) begin
      act_regs_data_3_4_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_3_4_sva_dfm_2_30_26,
          act_regs_data_2_5_sva_8_30_26, act_regs_data_3_4_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_4_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2565_enex5 ) begin
      act_regs_data_3_4_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_3_4_sva_dfm_2_21_0,
          act_regs_data_2_5_sva_8_21_0, act_regs_data_3_4_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_3_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2566_enex5 ) begin
      act_regs_data_3_3_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_3_3_sva_dfm_2_30_26,
          act_regs_data_2_4_sva_8_30_26, act_regs_data_3_3_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_3_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2568_enex5 ) begin
      act_regs_data_3_3_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_3_3_sva_dfm_2_21_0,
          act_regs_data_2_4_sva_8_21_0, act_regs_data_3_3_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_2_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2569_enex5 ) begin
      act_regs_data_3_2_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_3_2_sva_dfm_2_30_26,
          act_regs_data_2_3_sva_8_30_26, act_regs_data_3_2_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_2_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2571_enex5 ) begin
      act_regs_data_3_2_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_3_2_sva_dfm_2_21_0,
          act_regs_data_2_3_sva_8_21_0, act_regs_data_3_2_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_1_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2572_enex5 ) begin
      act_regs_data_3_1_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_3_1_sva_dfm_2_30_26,
          act_regs_data_2_10_sva_8_30_26, act_regs_data_3_1_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_1_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2574_enex5 ) begin
      act_regs_data_3_1_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_3_1_sva_dfm_2_21_0,
          act_regs_data_2_10_sva_8_21_0, act_regs_data_3_1_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_0_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2575_enex5 ) begin
      act_regs_data_3_0_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_3_0_sva_dfm_2_30_26,
          act_regs_data_2_1_sva_8_30_26, act_regs_data_3_0_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_0_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2577_enex5 ) begin
      act_regs_data_3_0_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_3_0_sva_dfm_2_21_0,
          act_regs_data_2_1_sva_8_21_0, act_regs_data_3_0_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_15_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2578_enex5 ) begin
      act_regs_data_2_15_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_2_15_sva_dfm_2_30_26,
          act_regs_data_1_2_sva_8_30_26, act_regs_data_2_15_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_15_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2580_enex5 ) begin
      act_regs_data_2_15_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_2_15_sva_dfm_2_21_0,
          act_regs_data_1_2_sva_8_21_0, act_regs_data_2_15_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_14_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2581_enex5 ) begin
      act_regs_data_2_14_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_2_14_sva_dfm_2_30_26,
          act_regs_data_1_15_sva_8_30_26, act_regs_data_2_14_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_14_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2583_enex5 ) begin
      act_regs_data_2_14_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_2_14_sva_dfm_2_21_0,
          act_regs_data_1_15_sva_8_21_0, act_regs_data_2_14_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_13_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2584_enex5 ) begin
      act_regs_data_2_13_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_2_13_sva_dfm_2_30_26,
          act_regs_data_1_14_sva_8_30_26, act_regs_data_2_13_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_13_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2586_enex5 ) begin
      act_regs_data_2_13_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_2_13_sva_dfm_2_21_0,
          act_regs_data_1_14_sva_8_21_0, act_regs_data_2_13_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_12_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2587_enex5 ) begin
      act_regs_data_2_12_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_2_12_sva_dfm_2_30_26,
          act_regs_data_1_13_sva_8_30_26, act_regs_data_2_12_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_12_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2589_enex5 ) begin
      act_regs_data_2_12_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_2_12_sva_dfm_2_21_0,
          act_regs_data_1_13_sva_8_21_0, act_regs_data_2_12_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_11_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2590_enex5 ) begin
      act_regs_data_2_11_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_2_11_sva_dfm_2_30_26,
          act_regs_data_1_12_sva_8_30_26, act_regs_data_2_11_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_11_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2592_enex5 ) begin
      act_regs_data_2_11_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_2_11_sva_dfm_2_21_0,
          act_regs_data_1_12_sva_8_21_0, act_regs_data_2_11_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_10_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2593_enex5 ) begin
      act_regs_data_2_10_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_2_10_sva_dfm_2_30_26,
          act_regs_data_1_11_sva_8_30_26, act_regs_data_2_10_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_10_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2595_enex5 ) begin
      act_regs_data_2_10_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_2_10_sva_dfm_2_21_0,
          act_regs_data_1_11_sva_8_21_0, act_regs_data_2_10_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_9_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2596_enex5 ) begin
      act_regs_data_2_9_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_2_9_sva_dfm_2_30_26,
          act_regs_data_2_0_sva_8_30_26, act_regs_data_2_9_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_9_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2598_enex5 ) begin
      act_regs_data_2_9_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_2_9_sva_dfm_2_21_0,
          act_regs_data_2_0_sva_8_21_0, act_regs_data_2_9_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_8_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2599_enex5 ) begin
      act_regs_data_2_8_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_2_8_sva_dfm_2_30_26,
          act_regs_data_1_9_sva_8_30_26, act_regs_data_2_8_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_8_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2601_enex5 ) begin
      act_regs_data_2_8_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_2_8_sva_dfm_2_21_0,
          act_regs_data_1_9_sva_8_21_0, act_regs_data_2_8_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_7_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2602_enex5 ) begin
      act_regs_data_2_7_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_2_7_sva_dfm_2_30_26,
          act_regs_data_1_8_sva_8_30_26, act_regs_data_2_7_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_7_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2604_enex5 ) begin
      act_regs_data_2_7_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_2_7_sva_dfm_2_21_0,
          act_regs_data_1_8_sva_8_21_0, act_regs_data_2_7_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_6_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2605_enex5 ) begin
      act_regs_data_2_6_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_2_6_sva_dfm_2_30_26,
          act_regs_data_1_7_sva_8_30_26, act_regs_data_2_6_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_6_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2607_enex5 ) begin
      act_regs_data_2_6_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_2_6_sva_dfm_2_21_0,
          act_regs_data_1_7_sva_8_21_0, act_regs_data_2_6_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_5_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2608_enex5 ) begin
      act_regs_data_2_5_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_2_5_sva_dfm_2_30_26,
          act_regs_data_1_6_sva_8_30_26, act_regs_data_2_5_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_5_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2610_enex5 ) begin
      act_regs_data_2_5_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_2_5_sva_dfm_2_21_0,
          act_regs_data_1_6_sva_8_21_0, act_regs_data_2_5_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_4_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2611_enex5 ) begin
      act_regs_data_2_4_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_2_4_sva_dfm_2_30_26,
          act_regs_data_1_5_sva_8_30_26, act_regs_data_2_4_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_4_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2613_enex5 ) begin
      act_regs_data_2_4_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_2_4_sva_dfm_2_21_0,
          act_regs_data_1_5_sva_8_21_0, act_regs_data_2_4_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_3_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2614_enex5 ) begin
      act_regs_data_2_3_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_2_3_sva_dfm_2_30_26,
          act_regs_data_1_4_sva_8_30_26, act_regs_data_2_3_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_3_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2616_enex5 ) begin
      act_regs_data_2_3_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_2_3_sva_dfm_2_21_0,
          act_regs_data_1_4_sva_8_21_0, act_regs_data_2_3_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_2_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2617_enex5 ) begin
      act_regs_data_2_2_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_2_2_sva_dfm_2_30_26,
          act_regs_data_1_3_sva_8_30_26, act_regs_data_2_2_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_2_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2619_enex5 ) begin
      act_regs_data_2_2_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_2_2_sva_dfm_2_21_0,
          act_regs_data_1_3_sva_8_21_0, act_regs_data_2_2_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_1_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2620_enex5 ) begin
      act_regs_data_2_1_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_2_1_sva_dfm_2_30_26,
          act_regs_data_1_10_sva_8_30_26, act_regs_data_2_1_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_1_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2622_enex5 ) begin
      act_regs_data_2_1_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_2_1_sva_dfm_2_21_0,
          act_regs_data_1_10_sva_8_21_0, act_regs_data_2_1_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_0_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2623_enex5 ) begin
      act_regs_data_2_0_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_2_0_sva_dfm_2_30_26,
          act_regs_data_1_1_sva_8_30_26, act_regs_data_2_0_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_0_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2625_enex5 ) begin
      act_regs_data_2_0_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_2_0_sva_dfm_2_21_0,
          act_regs_data_1_1_sva_8_21_0, act_regs_data_2_0_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_15_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2626_enex5 ) begin
      act_regs_data_1_15_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_1_15_sva_dfm_2_30_26,
          act_regs_data_0_2_sva_8_30_26, act_regs_data_1_15_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_15_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2628_enex5 ) begin
      act_regs_data_1_15_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_1_15_sva_dfm_2_21_0,
          act_regs_data_0_2_sva_8_21_0, act_regs_data_1_15_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_14_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2629_enex5 ) begin
      act_regs_data_1_14_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_1_14_sva_dfm_2_30_26,
          act_regs_data_0_15_sva_8_30_26, act_regs_data_1_14_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_14_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2631_enex5 ) begin
      act_regs_data_1_14_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_1_14_sva_dfm_2_21_0,
          act_regs_data_0_15_sva_8_21_0, act_regs_data_1_14_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_13_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2632_enex5 ) begin
      act_regs_data_1_13_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_1_13_sva_dfm_2_30_26,
          act_regs_data_0_14_sva_8_30_26, act_regs_data_1_13_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_13_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2634_enex5 ) begin
      act_regs_data_1_13_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_1_13_sva_dfm_2_21_0,
          act_regs_data_0_14_sva_8_21_0, act_regs_data_1_13_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_12_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2635_enex5 ) begin
      act_regs_data_1_12_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_1_12_sva_dfm_2_30_26,
          act_regs_data_0_13_sva_8_30_26, act_regs_data_1_12_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_12_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2637_enex5 ) begin
      act_regs_data_1_12_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_1_12_sva_dfm_2_21_0,
          act_regs_data_0_13_sva_8_21_0, act_regs_data_1_12_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_11_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2638_enex5 ) begin
      act_regs_data_1_11_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_1_11_sva_dfm_2_30_26,
          act_regs_data_0_12_sva_8_30_26, act_regs_data_1_11_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_11_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2640_enex5 ) begin
      act_regs_data_1_11_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_1_11_sva_dfm_2_21_0,
          act_regs_data_0_12_sva_8_21_0, act_regs_data_1_11_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_10_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2641_enex5 ) begin
      act_regs_data_1_10_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_1_10_sva_dfm_2_30_26,
          act_regs_data_0_11_sva_8_30_26, act_regs_data_1_10_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_10_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2643_enex5 ) begin
      act_regs_data_1_10_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_1_10_sva_dfm_2_21_0,
          act_regs_data_0_11_sva_8_21_0, act_regs_data_1_10_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_9_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2644_enex5 ) begin
      act_regs_data_1_9_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_1_9_sva_dfm_2_30_26,
          act_regs_data_1_0_sva_8_30_26, act_regs_data_1_9_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_9_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2646_enex5 ) begin
      act_regs_data_1_9_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_1_9_sva_dfm_2_21_0,
          act_regs_data_1_0_sva_8_21_0, act_regs_data_1_9_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_8_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2647_enex5 ) begin
      act_regs_data_1_8_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_1_8_sva_dfm_2_30_26,
          act_regs_data_0_9_sva_8_30_26, act_regs_data_1_8_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_8_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2649_enex5 ) begin
      act_regs_data_1_8_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_1_8_sva_dfm_2_21_0,
          act_regs_data_0_9_sva_8_21_0, act_regs_data_1_8_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_7_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2650_enex5 ) begin
      act_regs_data_1_7_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_1_7_sva_dfm_2_30_26,
          act_regs_data_0_8_sva_8_30_26, act_regs_data_1_7_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_7_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2652_enex5 ) begin
      act_regs_data_1_7_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_1_7_sva_dfm_2_21_0,
          act_regs_data_0_8_sva_8_21_0, act_regs_data_1_7_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_6_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2653_enex5 ) begin
      act_regs_data_1_6_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_1_6_sva_dfm_2_30_26,
          act_regs_data_0_7_sva_8_30_26, act_regs_data_1_6_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_6_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2655_enex5 ) begin
      act_regs_data_1_6_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_1_6_sva_dfm_2_21_0,
          act_regs_data_0_7_sva_8_21_0, act_regs_data_1_6_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_5_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2656_enex5 ) begin
      act_regs_data_1_5_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_1_5_sva_dfm_2_30_26,
          act_regs_data_0_6_sva_8_30_26, act_regs_data_1_5_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_5_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2658_enex5 ) begin
      act_regs_data_1_5_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_1_5_sva_dfm_2_21_0,
          act_regs_data_0_6_sva_8_21_0, act_regs_data_1_5_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_4_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2659_enex5 ) begin
      act_regs_data_1_4_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_1_4_sva_dfm_2_30_26,
          act_regs_data_0_5_sva_8_30_26, act_regs_data_1_4_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_4_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2661_enex5 ) begin
      act_regs_data_1_4_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_1_4_sva_dfm_2_21_0,
          act_regs_data_0_5_sva_8_21_0, act_regs_data_1_4_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_3_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2662_enex5 ) begin
      act_regs_data_1_3_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_1_3_sva_dfm_2_30_26,
          act_regs_data_0_4_sva_8_30_26, act_regs_data_1_3_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_3_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2664_enex5 ) begin
      act_regs_data_1_3_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_1_3_sva_dfm_2_21_0,
          act_regs_data_0_4_sva_8_21_0, act_regs_data_1_3_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_2_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2665_enex5 ) begin
      act_regs_data_1_2_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_1_2_sva_dfm_2_30_26,
          act_regs_data_0_3_sva_8_30_26, act_regs_data_1_2_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_2_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2667_enex5 ) begin
      act_regs_data_1_2_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_1_2_sva_dfm_2_21_0,
          act_regs_data_0_3_sva_8_21_0, act_regs_data_1_2_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_1_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2668_enex5 ) begin
      act_regs_data_1_1_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_1_1_sva_dfm_2_30_26,
          act_regs_data_0_10_sva_8_30_26, act_regs_data_1_1_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_1_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2670_enex5 ) begin
      act_regs_data_1_1_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_1_1_sva_dfm_2_21_0,
          act_regs_data_0_10_sva_8_21_0, act_regs_data_1_1_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_0_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2671_enex5 ) begin
      act_regs_data_1_0_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_1_0_sva_dfm_2_30_26,
          act_regs_data_0_1_sva_8_30_26, act_regs_data_1_0_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_0_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2673_enex5 ) begin
      act_regs_data_1_0_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_1_0_sva_dfm_2_21_0,
          act_regs_data_0_1_sva_8_21_0, act_regs_data_1_0_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_15_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2674_enex5 ) begin
      act_regs_data_0_15_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_0_15_sva_dfm_2_30_26,
          ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_1_30_26, act_regs_data_0_15_sva_8_30_26,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_15_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2676_enex5 ) begin
      act_regs_data_0_15_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_0_15_sva_dfm_2_21_0,
          Silu_for_3_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0,
          act_regs_data_0_15_sva_8_21_0, {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1
          , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_14_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2677_enex5 ) begin
      act_regs_data_0_14_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_0_14_sva_dfm_2_30_26,
          ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_1_30_26, act_regs_data_0_14_sva_8_30_26,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_14_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2679_enex5 ) begin
      act_regs_data_0_14_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_0_14_sva_dfm_2_21_0,
          Silu_for_2_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0,
          act_regs_data_0_14_sva_8_21_0, {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1
          , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_9_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2680_enex5 ) begin
      act_regs_data_0_9_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_0_9_sva_dfm_2_30_26,
          act_regs_data_0_0_sva_8_30_26, act_regs_data_0_9_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_9_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2682_enex5 ) begin
      act_regs_data_0_9_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_0_9_sva_dfm_2_21_0,
          act_regs_data_0_0_sva_8_21_0, act_regs_data_0_9_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_8_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2683_enex5 ) begin
      act_regs_data_0_8_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_0_8_sva_dfm_2_30_26,
          ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_1_30_26, act_regs_data_0_8_sva_8_30_26,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_8_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2685_enex5 ) begin
      act_regs_data_0_8_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_0_8_sva_dfm_2_21_0,
          Silu_for_y_8_sva_3_21_0, act_regs_data_0_8_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_7_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2686_enex5 ) begin
      act_regs_data_0_7_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_0_7_sva_dfm_2_30_26,
          ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_1_30_26, act_regs_data_0_7_sva_8_30_26,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_7_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2688_enex5 ) begin
      act_regs_data_0_7_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_0_7_sva_dfm_2_21_0,
          Silu_for_y_1_sva_3_21_0, act_regs_data_0_7_sva_8_21_0, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_6_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2689_enex5 ) begin
      act_regs_data_0_6_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_0_6_sva_dfm_2_30_26,
          ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_1_30_26, act_regs_data_0_6_sva_8_30_26,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_6_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2691_enex5 ) begin
      act_regs_data_0_6_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_0_6_sva_dfm_2_21_0,
          Silu_for_9_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0,
          act_regs_data_0_6_sva_8_21_0, {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1
          , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_5_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2692_enex5 ) begin
      act_regs_data_0_5_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_0_5_sva_dfm_2_30_26,
          ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_1_30_26, act_regs_data_0_5_sva_8_30_26,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_5_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2694_enex5 ) begin
      act_regs_data_0_5_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_0_5_sva_dfm_2_21_0,
          Silu_for_7_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0,
          act_regs_data_0_5_sva_8_21_0, {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1
          , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_4_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2695_enex5 ) begin
      act_regs_data_0_4_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_0_4_sva_dfm_2_30_26,
          ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_1_30_26, act_regs_data_0_4_sva_8_30_26,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_4_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2697_enex5 ) begin
      act_regs_data_0_4_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_0_4_sva_dfm_2_21_0,
          Silu_for_6_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0,
          act_regs_data_0_4_sva_8_21_0, {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1
          , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_3_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2698_enex5 ) begin
      act_regs_data_0_3_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_0_3_sva_dfm_2_30_26,
          ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_1_30_26, act_regs_data_0_3_sva_8_30_26,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_3_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2700_enex5 ) begin
      act_regs_data_0_3_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_0_3_sva_dfm_2_21_0,
          Silu_for_5_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0,
          act_regs_data_0_3_sva_8_21_0, {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1
          , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_2_sva_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2701_enex5 ) begin
      act_regs_data_0_2_sva_30_26 <= MUX1HOT_v_5_3_2(act_regs_data_0_2_sva_dfm_2_30_26,
          ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_1_30_26, act_regs_data_0_2_sva_8_30_26,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_2_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2703_enex5 ) begin
      act_regs_data_0_2_sva_21_0 <= MUX1HOT_v_22_3_2(act_regs_data_0_2_sva_dfm_2_21_0,
          Silu_for_4_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0,
          act_regs_data_0_2_sva_8_21_0, {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1
          , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_31_0 <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_read_read_data_and_16_enex5 ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_31_0 <= act_mem_banks_read_for_mux_15_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_63_32 <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_read_read_data_and_17_enex5 ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_63_32 <= act_mem_banks_read_for_mux_14_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_95_64 <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_read_read_data_and_18_enex5 ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_95_64 <= act_mem_banks_read_for_mux_13_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_127_96 <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_read_read_data_and_19_enex5 ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_127_96 <= act_mem_banks_read_for_mux_12_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_159_128 <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_read_read_data_and_20_enex5 ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_159_128 <= act_mem_banks_read_for_mux_11_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_191_160 <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_read_read_data_and_21_enex5 ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_191_160 <= act_mem_banks_read_for_mux_10_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_223_192 <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_read_read_data_and_22_enex5 ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_223_192 <= act_mem_banks_read_for_mux_9_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_255_224 <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_read_read_data_and_23_enex5 ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_255_224 <= act_mem_banks_read_for_mux_8_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_287_256 <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_read_read_data_and_24_enex5 ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_287_256 <= act_mem_banks_read_for_mux_7_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_319_288 <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_read_read_data_and_25_enex5 ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_319_288 <= act_mem_banks_read_for_mux_6_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_351_320 <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_read_read_data_and_26_enex5 ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_351_320 <= act_mem_banks_read_for_mux_5_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_383_352 <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_read_read_data_and_27_enex5 ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_383_352 <= act_mem_banks_read_for_mux_4_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_415_384 <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_read_read_data_and_28_enex5 ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_415_384 <= act_mem_banks_read_for_mux_3_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_447_416 <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_read_read_data_and_29_enex5 ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_447_416 <= act_mem_banks_read_for_mux_2_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_479_448 <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_read_read_data_and_30_enex5 ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_479_448 <= act_mem_banks_read_for_mux_1_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_511_480 <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_read_read_data_and_31_enex5 ) begin
      act_mem_banks_read_read_data_lpi_1_dfm_1_511_480 <= act_mem_banks_read_for_mux_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_read_out_data_0_0_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_port_read_out_data_and_16_enex5 ) begin
      act_port_read_out_data_0_0_sva_dfm <= act_mem_banks_read_read_data_lpi_1_dfm_1_31_0_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_read_out_data_0_1_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_port_read_out_data_and_17_enex5 ) begin
      act_port_read_out_data_0_1_sva_dfm <= act_mem_banks_read_read_data_lpi_1_dfm_1_63_32_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_read_out_data_0_2_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_port_read_out_data_and_18_enex5 ) begin
      act_port_read_out_data_0_2_sva_dfm <= act_mem_banks_read_read_data_lpi_1_dfm_1_95_64_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_read_out_data_0_3_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_port_read_out_data_and_19_enex5 ) begin
      act_port_read_out_data_0_3_sva_dfm <= act_mem_banks_read_read_data_lpi_1_dfm_1_127_96_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_read_out_data_0_4_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_port_read_out_data_and_20_enex5 ) begin
      act_port_read_out_data_0_4_sva_dfm <= act_mem_banks_read_read_data_lpi_1_dfm_1_159_128_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_read_out_data_0_5_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_port_read_out_data_and_21_enex5 ) begin
      act_port_read_out_data_0_5_sva_dfm <= act_mem_banks_read_read_data_lpi_1_dfm_1_191_160_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_read_out_data_0_6_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_port_read_out_data_and_22_enex5 ) begin
      act_port_read_out_data_0_6_sva_dfm <= act_mem_banks_read_read_data_lpi_1_dfm_1_223_192_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_read_out_data_0_7_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_port_read_out_data_and_23_enex5 ) begin
      act_port_read_out_data_0_7_sva_dfm <= act_mem_banks_read_read_data_lpi_1_dfm_1_255_224_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_read_out_data_0_8_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_port_read_out_data_and_24_enex5 ) begin
      act_port_read_out_data_0_8_sva_dfm <= act_mem_banks_read_read_data_lpi_1_dfm_1_287_256_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_read_out_data_0_9_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_port_read_out_data_and_25_enex5 ) begin
      act_port_read_out_data_0_9_sva_dfm <= act_mem_banks_read_read_data_lpi_1_dfm_1_319_288_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_read_out_data_0_10_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_port_read_out_data_and_26_enex5 ) begin
      act_port_read_out_data_0_10_sva_dfm <= act_mem_banks_read_read_data_lpi_1_dfm_1_351_320_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_read_out_data_0_11_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_port_read_out_data_and_27_enex5 ) begin
      act_port_read_out_data_0_11_sva_dfm <= act_mem_banks_read_read_data_lpi_1_dfm_1_383_352_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_read_out_data_0_12_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_port_read_out_data_and_28_enex5 ) begin
      act_port_read_out_data_0_12_sva_dfm <= act_mem_banks_read_read_data_lpi_1_dfm_1_415_384_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_read_out_data_0_13_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_port_read_out_data_and_29_enex5 ) begin
      act_port_read_out_data_0_13_sva_dfm <= act_mem_banks_read_read_data_lpi_1_dfm_1_447_416_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_read_out_data_0_14_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_port_read_out_data_and_30_enex5 ) begin
      act_port_read_out_data_0_14_sva_dfm <= act_mem_banks_read_read_data_lpi_1_dfm_1_479_448_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_port_read_out_data_0_15_sva_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_port_read_out_data_and_31_enex5 ) begin
      act_port_read_out_data_0_15_sva_dfm <= act_mem_banks_read_read_data_lpi_1_dfm_1_511_480_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_1_else_if_acc_itm <= 4'b0000;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_596 | or_dcpl_593 | (~ Gelu_for_1_slc_32_1_svs)))
        & and_dcpl_1112 & (~ Gelu_for_1_else_slc_32_svs) ) begin
      Gelu_for_1_else_if_acc_itm <= Gelu_for_1_else_if_acc_itm_mx1w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_2_else_if_acc_itm <= 4'b0000;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_596 | or_dcpl_593 | (~ Gelu_for_2_slc_32_1_svs)))
        & and_dcpl_1112 & (~ Gelu_for_2_else_slc_32_svs) ) begin
      Gelu_for_2_else_if_acc_itm <= Gelu_for_2_else_if_acc_itm_mx1w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_3_else_if_acc_itm <= 4'b0000;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_596 | or_dcpl_593 | (~ Gelu_for_3_slc_32_1_svs)))
        & and_dcpl_1112 & (~ Gelu_for_3_else_slc_32_svs) ) begin
      Gelu_for_3_else_if_acc_itm <= Gelu_for_3_else_if_acc_itm_mx1w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_4_else_if_acc_itm <= 4'b0000;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_596 | or_dcpl_593 | (~ Gelu_for_4_slc_32_1_svs)))
        & and_dcpl_1112 & (~ Gelu_for_4_else_slc_32_svs) ) begin
      Gelu_for_4_else_if_acc_itm <= Gelu_for_4_else_if_acc_itm_mx1w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_5_else_if_acc_itm <= 4'b0000;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_596 | or_dcpl_593 | (~ Gelu_for_5_slc_32_1_svs)))
        & and_dcpl_1112 & (~ Gelu_for_5_else_slc_32_svs) ) begin
      Gelu_for_5_else_if_acc_itm <= Gelu_for_5_else_if_acc_itm_mx1w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_6_else_if_acc_itm <= 4'b0000;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_596 | or_dcpl_593 | (~ Gelu_for_6_slc_32_1_svs)))
        & and_dcpl_1112 & (~ Gelu_for_6_else_slc_32_svs) ) begin
      Gelu_for_6_else_if_acc_itm <= Gelu_for_6_else_if_acc_itm_mx1w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_7_else_if_acc_itm <= 4'b0000;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_596 | or_dcpl_593 | (~ Gelu_for_7_slc_32_1_svs)))
        & and_dcpl_1112 & (~ Gelu_for_7_else_slc_32_svs) ) begin
      Gelu_for_7_else_if_acc_itm <= Gelu_for_7_else_if_acc_itm_mx1w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_8_else_if_acc_itm <= 4'b0000;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_596 | or_dcpl_593 | (~ Gelu_for_8_slc_32_1_svs)))
        & and_dcpl_1112 & (~ Gelu_for_8_else_slc_32_svs) ) begin
      Gelu_for_8_else_if_acc_itm <= Gelu_for_8_else_if_acc_itm_mx1w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_1_else_else_if_acc_itm <= 2'b00;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_616 | (act_config_in_InstFetch_return_sva_7_2[2])
        | (~ Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)))
        & and_dcpl_331 & and_dcpl_40 & (~ Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
        & Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
        ) begin
      Silu_for_1_else_else_if_acc_itm <= nl_Silu_for_1_else_else_if_acc_itm[1:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_623 | (~((fsm_output[0]) & operator_32_8_true_AC_TRN_AC_WRAP_less_15_tmp))
        | (fsm_output[1]) | or_dcpl_457)) ) begin
      Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_1_less_15_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_else_and_1_m1c <= 1'b0;
    end
    else if ( ActUnitRun_wen & and_dcpl_1116 & (~ (act_config_in_InstFetch_return_sva_7_2[2]))
        & Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
        & (~ (fsm_output[1])) & and_dcpl_1061 ) begin
      Silu_for_else_and_1_m1c <= Silu_for_else_and_1_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_2_else_else_if_acc_itm <= 2'b00;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_616 | (act_config_in_InstFetch_return_sva_7_2[2])
        | (~ Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)))
        & and_dcpl_331 & and_dcpl_40 & (~ Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
        & Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
        ) begin
      Silu_for_2_else_else_if_acc_itm <= nl_Silu_for_2_else_else_if_acc_itm[1:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_623 | (~((fsm_output[0]) & operator_32_8_true_AC_TRN_AC_WRAP_less_14_tmp))
        | (fsm_output[1]) | or_dcpl_457)) ) begin
      Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_1_less_14_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_else_and_3_m1c <= 1'b0;
    end
    else if ( ActUnitRun_wen & and_dcpl_1116 & and_dcpl_1118 & Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
        & and_dcpl_1061 ) begin
      Silu_for_else_and_3_m1c <= Silu_for_else_and_3_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_3_else_else_if_acc_itm <= 2'b00;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_616 | (act_config_in_InstFetch_return_sva_7_2[2])
        | (~ Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)))
        & and_dcpl_331 & and_dcpl_40 & (~ Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
        & Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
        ) begin
      Silu_for_3_else_else_if_acc_itm <= nl_Silu_for_3_else_else_if_acc_itm[1:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_623 | (~((fsm_output[0]) & operator_32_8_true_AC_TRN_AC_WRAP_less_13_tmp))
        | (fsm_output[1]) | or_dcpl_457)) ) begin
      Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_1_less_13_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_else_and_5_m1c <= 1'b0;
    end
    else if ( ActUnitRun_wen & and_dcpl_1116 & and_dcpl_1118 & Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
        & and_dcpl_1061 ) begin
      Silu_for_else_and_5_m1c <= Silu_for_else_and_5_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_4_else_else_if_acc_itm <= 2'b00;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_616 | (act_config_in_InstFetch_return_sva_7_2[2])
        | (~ Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)))
        & and_dcpl_331 & and_dcpl_40 & (~ Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
        & Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
        ) begin
      Silu_for_4_else_else_if_acc_itm <= nl_Silu_for_4_else_else_if_acc_itm[1:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_623 | (~((fsm_output[0]) & operator_32_8_true_AC_TRN_AC_WRAP_less_12_tmp))
        | (fsm_output[1]) | or_dcpl_457)) ) begin
      Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_1_less_12_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_else_and_7_m1c <= 1'b0;
    end
    else if ( ActUnitRun_wen & and_dcpl_1116 & and_dcpl_1118 & Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
        & and_dcpl_1061 ) begin
      Silu_for_else_and_7_m1c <= Silu_for_else_and_7_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_5_else_else_if_acc_itm <= 2'b00;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_616 | (act_config_in_InstFetch_return_sva_7_2[2])
        | (~ Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)))
        & and_dcpl_331 & and_dcpl_40 & (~ Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
        & Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
        ) begin
      Silu_for_5_else_else_if_acc_itm <= nl_Silu_for_5_else_else_if_acc_itm[1:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_623 | (~((fsm_output[0]) & operator_32_8_true_AC_TRN_AC_WRAP_less_11_tmp))
        | (fsm_output[1]) | or_dcpl_457)) ) begin
      Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_1_less_11_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_else_and_9_m1c <= 1'b0;
    end
    else if ( ActUnitRun_wen & and_dcpl_1116 & and_dcpl_1118 & Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
        & and_dcpl_1061 ) begin
      Silu_for_else_and_9_m1c <= Silu_for_else_and_9_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_6_else_else_if_acc_itm <= 2'b00;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_616 | (act_config_in_InstFetch_return_sva_7_2[2])
        | (~ Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)))
        & and_dcpl_331 & and_dcpl_40 & (~ Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
        & Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
        ) begin
      Silu_for_6_else_else_if_acc_itm <= nl_Silu_for_6_else_else_if_acc_itm[1:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_623 | (~((fsm_output[0]) & operator_32_8_true_AC_TRN_AC_WRAP_less_10_tmp))
        | (fsm_output[1]) | or_dcpl_457)) ) begin
      Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_1_less_10_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_else_and_11_m1c <= 1'b0;
    end
    else if ( ActUnitRun_wen & and_dcpl_1116 & and_dcpl_1118 & Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
        & and_dcpl_1061 ) begin
      Silu_for_else_and_11_m1c <= Silu_for_else_and_11_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_7_else_else_if_acc_itm <= 2'b00;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_616 | (act_config_in_InstFetch_return_sva_7_2[2])
        | (~ Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)))
        & and_dcpl_331 & and_dcpl_40 & (~ Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
        & Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
        ) begin
      Silu_for_7_else_else_if_acc_itm <= nl_Silu_for_7_else_else_if_acc_itm[1:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_623 | (~((fsm_output[0]) & operator_32_8_true_AC_TRN_AC_WRAP_less_9_tmp))
        | (fsm_output[1]) | or_dcpl_457)) ) begin
      Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_1_less_9_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_else_and_13_m1c <= 1'b0;
    end
    else if ( ActUnitRun_wen & and_dcpl_1116 & and_dcpl_1118 & Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
        & and_dcpl_1061 ) begin
      Silu_for_else_and_13_m1c <= Silu_for_else_and_13_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_8_else_else_if_acc_itm <= 2'b00;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_616 | (act_config_in_InstFetch_return_sva_7_2[2])
        | (~ Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)))
        & and_dcpl_331 & and_dcpl_40 & (~ Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
        & Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
        ) begin
      Silu_for_8_else_else_if_acc_itm <= nl_Silu_for_8_else_else_if_acc_itm[1:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_623 | (~((fsm_output[0]) & operator_32_8_true_AC_TRN_AC_WRAP_less_8_tmp))
        | (fsm_output[1]) | or_dcpl_457)) ) begin
      Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_1_less_8_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_else_and_15_m1c <= 1'b0;
    end
    else if ( ActUnitRun_wen & and_dcpl_1116 & and_dcpl_1118 & Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
        & and_dcpl_1061 ) begin
      Silu_for_else_and_15_m1c <= Silu_for_else_and_15_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_623 | (~((fsm_output[0]) & operator_32_8_true_AC_TRN_AC_WRAP_less_7_tmp))
        | (fsm_output[1]) | or_dcpl_457)) ) begin
      Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= $signed(26'b10000000000000000000000000) < $signed(({nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
          , nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
          , nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          , nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
          , nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_623 | (~((fsm_output[0]) & operator_32_8_true_AC_TRN_AC_WRAP_less_6_tmp))
        | (fsm_output[1]) | or_dcpl_457)) ) begin
      Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= $signed(26'b10000000000000000000000000) < $signed(({nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
          , nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
          , nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          , nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
          , nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_623 | (~((fsm_output[0]) & operator_32_8_true_AC_TRN_AC_WRAP_less_5_tmp))
        | (fsm_output[1]) | or_dcpl_457)) ) begin
      Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= $signed(26'b10000000000000000000000000) < $signed(({nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
          , nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
          , nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          , nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
          , nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_623 | (~((fsm_output[0]) & operator_32_8_true_AC_TRN_AC_WRAP_less_4_tmp))
        | (fsm_output[1]) | or_dcpl_457)) ) begin
      Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= $signed(26'b10000000000000000000000000) < $signed(({nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
          , nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
          , nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          , nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
          , nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_623 | (~((fsm_output[0]) & operator_32_8_true_AC_TRN_AC_WRAP_less_3_tmp))
        | (fsm_output[1]) | or_dcpl_457)) ) begin
      Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= $signed(26'b10000000000000000000000000) < $signed(({nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
          , nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
          , nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          , nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
          , nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_623 | (~((fsm_output[0]) & operator_32_8_true_AC_TRN_AC_WRAP_less_2_tmp))
        | (fsm_output[1]) | or_dcpl_457)) ) begin
      Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= $signed(26'b10000000000000000000000000) < $signed(({nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
          , nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
          , nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          , nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
          , nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_623 | (~((fsm_output[0]) & operator_32_8_true_AC_TRN_AC_WRAP_less_1_tmp))
        | (fsm_output[1]) | or_dcpl_457)) ) begin
      Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= $signed(26'b10000000000000000000000000) < $signed(({nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
          , nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
          , nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          , nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
          , nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_623 | (~((fsm_output[0]) & operator_32_8_true_AC_TRN_AC_WRAP_less_tmp))
        | (fsm_output[1]) | or_dcpl_457)) ) begin
      Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
          <= $signed(26'b10000000000000000000000000) < $signed(({nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
          , nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
          , nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          , nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
          , nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_1_else_slc_32_svs <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_717 | (~((fsm_output[0]) & Gelu_for_if_less_15_tmp))
        | (fsm_output[1]) | or_dcpl_457)) ) begin
      Gelu_for_1_else_slc_32_svs <= Gelu_for_else_if_less_15_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_2_else_slc_32_svs <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_717 | (~((fsm_output[0]) & Gelu_for_if_less_14_tmp))
        | (fsm_output[1]) | or_dcpl_457)) ) begin
      Gelu_for_2_else_slc_32_svs <= Gelu_for_else_if_less_14_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_3_else_slc_32_svs <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_717 | (~((fsm_output[0]) & Gelu_for_if_less_13_tmp))
        | (fsm_output[1]) | or_dcpl_457)) ) begin
      Gelu_for_3_else_slc_32_svs <= Gelu_for_else_if_less_13_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_4_else_slc_32_svs <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_717 | (~((fsm_output[0]) & Gelu_for_if_less_12_tmp))
        | (fsm_output[1]) | or_dcpl_457)) ) begin
      Gelu_for_4_else_slc_32_svs <= Gelu_for_else_if_less_12_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_5_else_slc_32_svs <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_717 | (~((fsm_output[0]) & Gelu_for_if_less_11_tmp))
        | (fsm_output[1]) | or_dcpl_457)) ) begin
      Gelu_for_5_else_slc_32_svs <= Gelu_for_else_if_less_11_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_6_else_slc_32_svs <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_717 | (~((fsm_output[0]) & Gelu_for_if_less_10_tmp))
        | (fsm_output[1]) | or_dcpl_457)) ) begin
      Gelu_for_6_else_slc_32_svs <= Gelu_for_else_if_less_10_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_7_else_slc_32_svs <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_717 | (~((fsm_output[0]) & Gelu_for_if_less_9_tmp))
        | (fsm_output[1]) | or_dcpl_457)) ) begin
      Gelu_for_7_else_slc_32_svs <= Gelu_for_else_if_less_9_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_8_else_slc_32_svs <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_717 | (~((fsm_output[0]) & Gelu_for_if_less_8_tmp))
        | (fsm_output[1]) | or_dcpl_457)) ) begin
      Gelu_for_8_else_slc_32_svs <= Gelu_for_else_if_less_8_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_9_else_slc_32_svs <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_717 | (~((fsm_output[0]) & Gelu_for_if_less_7_tmp))
        | (fsm_output[1]) | or_dcpl_457)) ) begin
      Gelu_for_9_else_slc_32_svs <= $signed(25'b1010000000000000000000000) < $signed(({nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
          , nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
          , nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          , nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
          , nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_10_else_slc_32_svs <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_717 | (~((fsm_output[0]) & Gelu_for_if_less_6_tmp))
        | (fsm_output[1]) | or_dcpl_457)) ) begin
      Gelu_for_10_else_slc_32_svs <= $signed(25'b1010000000000000000000000) < $signed(({nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
          , nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
          , nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          , nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
          , nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_11_else_slc_32_svs <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_717 | (~((fsm_output[0]) & Gelu_for_if_less_5_tmp))
        | (fsm_output[1]) | or_dcpl_457)) ) begin
      Gelu_for_11_else_slc_32_svs <= $signed(25'b1010000000000000000000000) < $signed(({nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
          , nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
          , nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          , nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
          , nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_12_else_slc_32_svs <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_717 | (~((fsm_output[0]) & Gelu_for_if_less_4_tmp))
        | (fsm_output[1]) | or_dcpl_457)) ) begin
      Gelu_for_12_else_slc_32_svs <= $signed(25'b1010000000000000000000000) < $signed(({nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
          , nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
          , nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          , nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
          , nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_13_else_slc_32_svs <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_717 | (~((fsm_output[0]) & Gelu_for_if_less_3_tmp))
        | (fsm_output[1]) | or_dcpl_457)) ) begin
      Gelu_for_13_else_slc_32_svs <= $signed(25'b1010000000000000000000000) < $signed(({nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
          , nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
          , nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          , nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
          , nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_14_else_slc_32_svs <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_717 | (~((fsm_output[0]) & Gelu_for_if_less_2_tmp))
        | (fsm_output[1]) | or_dcpl_457)) ) begin
      Gelu_for_14_else_slc_32_svs <= $signed(25'b1010000000000000000000000) < $signed(({nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
          , nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
          , nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          , nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
          , nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_15_else_slc_32_svs <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_717 | (~((fsm_output[0]) & Gelu_for_if_less_1_tmp))
        | (fsm_output[1]) | or_dcpl_457)) ) begin
      Gelu_for_15_else_slc_32_svs <= $signed(25'b1010000000000000000000000) < $signed(({nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
          , nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
          , nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          , nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
          , nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_16_else_slc_32_svs <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_717 | (~((fsm_output[0]) & Gelu_for_if_less_tmp))
        | (fsm_output[1]) | or_dcpl_457)) ) begin
      Gelu_for_16_else_slc_32_svs <= $signed(25'b1010000000000000000000000) < $signed(({nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
          , nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
          , nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          , nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
          , nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_9_else_else_if_acc_itm <= 2'b00;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_616 | (act_config_in_InstFetch_return_sva_7_2[2])
        | (~ Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)))
        & and_dcpl_331 & and_dcpl_40 & (~ Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
        & Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
        ) begin
      Silu_for_9_else_else_if_acc_itm <= nl_Silu_for_9_else_else_if_acc_itm[1:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_else_and_17_m1c <= 1'b0;
    end
    else if ( ActUnitRun_wen & and_dcpl_1144 & (~ (act_config_in_InstFetch_return_sva_7_2[2]))
        & Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
        & (~ (fsm_output[1])) & and_dcpl_1061 ) begin
      Silu_for_else_and_17_m1c <= Silu_for_else_and_17_m1c_mx0w1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_10_else_else_if_acc_itm <= 2'b00;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_616 | (act_config_in_InstFetch_return_sva_7_2[2])
        | (~ Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)))
        & and_dcpl_331 & and_dcpl_40 & (~ Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
        & Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
        ) begin
      Silu_for_10_else_else_if_acc_itm <= nl_Silu_for_10_else_else_if_acc_itm[1:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_else_and_19_m1c <= 1'b0;
    end
    else if ( ActUnitRun_wen & and_dcpl_1144 & (~ (act_config_in_InstFetch_return_sva_7_2[2]))
        & Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
        & (~ (fsm_output[1])) & and_dcpl_1061 ) begin
      Silu_for_else_and_19_m1c <= Silu_for_else_and_19_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_11_else_else_if_acc_itm <= 2'b00;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_616 | (act_config_in_InstFetch_return_sva_7_2[2])
        | (~ Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)))
        & and_dcpl_331 & and_dcpl_40 & Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
        & (~ Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
        ) begin
      Silu_for_11_else_else_if_acc_itm <= nl_Silu_for_11_else_else_if_acc_itm[1:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_else_and_21_m1c <= 1'b0;
    end
    else if ( ActUnitRun_wen & and_dcpl_1144 & (~ (act_config_in_InstFetch_return_sva_7_2[2]))
        & Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
        & (~ (fsm_output[1])) & and_dcpl_1061 ) begin
      Silu_for_else_and_21_m1c <= Silu_for_else_and_21_m1c_mx0w1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_12_else_else_if_acc_itm <= 2'b00;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_616 | (act_config_in_InstFetch_return_sva_7_2[2])
        | (~ Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)))
        & and_dcpl_331 & and_dcpl_40 & Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
        & (~ Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
        ) begin
      Silu_for_12_else_else_if_acc_itm <= nl_Silu_for_12_else_else_if_acc_itm[1:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_else_and_23_m1c <= 1'b0;
    end
    else if ( ActUnitRun_wen & and_dcpl_1144 & (~ (act_config_in_InstFetch_return_sva_7_2[2]))
        & Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
        & (~ (fsm_output[1])) & and_dcpl_1061 ) begin
      Silu_for_else_and_23_m1c <= Silu_for_else_and_23_m1c_mx0w1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_13_else_else_if_acc_itm <= 2'b00;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_616 | (act_config_in_InstFetch_return_sva_7_2[2])
        | (~ Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)))
        & and_dcpl_331 & and_dcpl_40 & Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
        & (~ Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
        ) begin
      Silu_for_13_else_else_if_acc_itm <= nl_Silu_for_13_else_else_if_acc_itm[1:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_else_and_25_m1c <= 1'b0;
    end
    else if ( ActUnitRun_wen & and_dcpl_1144 & (~ (act_config_in_InstFetch_return_sva_7_2[2]))
        & Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
        & (~ (fsm_output[1])) & and_dcpl_1061 ) begin
      Silu_for_else_and_25_m1c <= Silu_for_else_and_25_m1c_mx0w1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_14_else_else_if_acc_itm <= 2'b00;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_616 | (act_config_in_InstFetch_return_sva_7_2[2])
        | (~ Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)))
        & and_dcpl_331 & and_dcpl_40 & Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
        & (~ Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
        ) begin
      Silu_for_14_else_else_if_acc_itm <= nl_Silu_for_14_else_else_if_acc_itm[1:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_else_and_27_m1c <= 1'b0;
    end
    else if ( ActUnitRun_wen & and_dcpl_1144 & (~ (act_config_in_InstFetch_return_sva_7_2[2]))
        & Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
        & (~ (fsm_output[1])) & and_dcpl_1061 ) begin
      Silu_for_else_and_27_m1c <= Silu_for_else_and_27_m1c_mx0w1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_15_else_else_if_acc_itm <= 2'b00;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_616 | (act_config_in_InstFetch_return_sva_7_2[2])
        | (~ Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)))
        & and_dcpl_331 & and_dcpl_40 & Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
        & (~ Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
        ) begin
      Silu_for_15_else_else_if_acc_itm <= nl_Silu_for_15_else_else_if_acc_itm[1:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_else_and_29_m1c <= 1'b0;
    end
    else if ( ActUnitRun_wen & and_dcpl_1144 & (~ (act_config_in_InstFetch_return_sva_7_2[2]))
        & Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
        & (~ (fsm_output[1])) & and_dcpl_1061 ) begin
      Silu_for_else_and_29_m1c <= Silu_for_else_and_29_m1c_mx0w1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_16_else_else_if_acc_itm <= 2'b00;
    end
    else if ( ActUnitRun_wen & (~(or_dcpl_616 | (act_config_in_InstFetch_return_sva_7_2[2])
        | (~ Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs)))
        & and_dcpl_331 & and_dcpl_40 & (~ Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs)
        & Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
        ) begin
      Silu_for_16_else_else_if_acc_itm <= nl_Silu_for_16_else_else_if_acc_itm[1:0];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_else_and_31_m1c <= 1'b0;
    end
    else if ( ActUnitRun_wen & and_dcpl_1144 & (~ (act_config_in_InstFetch_return_sva_7_2[2]))
        & Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
        & (~ (fsm_output[1])) & and_dcpl_1061 ) begin
      Silu_for_else_and_31_m1c <= Silu_for_else_and_31_m1c_mx0w1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_else_and_1_m1c <= 1'b0;
    end
    else if ( ActUnitRun_wen & and_dcpl_1144 & and_dcpl_1174 & Gelu_for_1_slc_32_1_svs
        & and_dcpl_1061 ) begin
      Gelu_for_else_and_1_m1c <= Gelu_for_else_and_1_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_else_and_3_m1c <= 1'b0;
    end
    else if ( ActUnitRun_wen & and_dcpl_1144 & and_dcpl_1174 & Gelu_for_2_slc_32_1_svs
        & and_dcpl_1061 ) begin
      Gelu_for_else_and_3_m1c <= Gelu_for_else_and_3_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_else_and_5_m1c <= 1'b0;
    end
    else if ( ActUnitRun_wen & and_dcpl_1144 & and_dcpl_1174 & Gelu_for_3_slc_32_1_svs
        & and_dcpl_1061 ) begin
      Gelu_for_else_and_5_m1c <= Gelu_for_else_and_5_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_else_and_7_m1c <= 1'b0;
    end
    else if ( ActUnitRun_wen & and_dcpl_1144 & and_dcpl_1174 & Gelu_for_4_slc_32_1_svs
        & and_dcpl_1061 ) begin
      Gelu_for_else_and_7_m1c <= Gelu_for_else_and_7_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_else_and_9_m1c <= 1'b0;
    end
    else if ( ActUnitRun_wen & and_dcpl_1144 & and_dcpl_1174 & Gelu_for_5_slc_32_1_svs
        & and_dcpl_1061 ) begin
      Gelu_for_else_and_9_m1c <= Gelu_for_else_and_9_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_else_and_11_m1c <= 1'b0;
    end
    else if ( ActUnitRun_wen & and_dcpl_1144 & and_dcpl_1174 & Gelu_for_6_slc_32_1_svs
        & and_dcpl_1061 ) begin
      Gelu_for_else_and_11_m1c <= Gelu_for_else_and_11_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_else_and_13_m1c <= 1'b0;
    end
    else if ( ActUnitRun_wen & and_dcpl_1144 & and_dcpl_1174 & Gelu_for_7_slc_32_1_svs
        & and_dcpl_1061 ) begin
      Gelu_for_else_and_13_m1c <= Gelu_for_else_and_13_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_else_and_15_m1c <= 1'b0;
    end
    else if ( ActUnitRun_wen & and_dcpl_1144 & and_dcpl_1174 & Gelu_for_8_slc_32_1_svs
        & and_dcpl_1061 ) begin
      Gelu_for_else_and_15_m1c <= Gelu_for_else_and_15_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_else_and_17_m1c <= 1'b0;
    end
    else if ( ActUnitRun_wen & and_dcpl_1144 & and_dcpl_1174 & Gelu_for_9_slc_32_1_svs
        & and_dcpl_1061 ) begin
      Gelu_for_else_and_17_m1c <= Gelu_for_else_and_17_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_else_and_19_m1c <= 1'b0;
    end
    else if ( ActUnitRun_wen & and_dcpl_1144 & and_dcpl_1174 & Gelu_for_10_slc_32_1_svs
        & and_dcpl_1061 ) begin
      Gelu_for_else_and_19_m1c <= Gelu_for_else_and_19_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_else_and_21_m1c <= 1'b0;
    end
    else if ( ActUnitRun_wen & and_dcpl_1144 & and_dcpl_1174 & Gelu_for_11_slc_32_1_svs
        & and_dcpl_1061 ) begin
      Gelu_for_else_and_21_m1c <= Gelu_for_else_and_21_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_else_and_23_m1c <= 1'b0;
    end
    else if ( ActUnitRun_wen & and_dcpl_1144 & and_dcpl_1174 & Gelu_for_12_slc_32_1_svs
        & and_dcpl_1061 ) begin
      Gelu_for_else_and_23_m1c <= Gelu_for_else_and_23_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_else_and_25_m1c <= 1'b0;
    end
    else if ( ActUnitRun_wen & and_dcpl_1144 & and_dcpl_1174 & Gelu_for_13_slc_32_1_svs
        & and_dcpl_1061 ) begin
      Gelu_for_else_and_25_m1c <= Gelu_for_else_and_25_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_else_and_27_m1c <= 1'b0;
    end
    else if ( ActUnitRun_wen & and_dcpl_1144 & and_dcpl_1174 & Gelu_for_14_slc_32_1_svs
        & and_dcpl_1061 ) begin
      Gelu_for_else_and_27_m1c <= Gelu_for_else_and_27_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_else_and_29_m1c <= 1'b0;
    end
    else if ( ActUnitRun_wen & and_dcpl_1144 & and_dcpl_1174 & Gelu_for_15_slc_32_1_svs
        & and_dcpl_1061 ) begin
      Gelu_for_else_and_29_m1c <= Gelu_for_else_and_29_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_else_and_31_m1c <= 1'b0;
    end
    else if ( ActUnitRun_wen & and_dcpl_1144 & (act_config_in_InstFetch_return_sva_7_2[2])
        & Gelu_for_16_slc_32_1_svs & (~ (fsm_output[1])) & and_dcpl_1061 ) begin
      Gelu_for_else_and_31_m1c <= Gelu_for_else_and_31_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_write_addrs_lpi_1_dfm_5 <= 5'b00000;
    end
    else if ( mux_622_nl & nor_1441_cse & (fsm_output[0]) & ActUnitRun_wen ) begin
      act_write_addrs_lpi_1_dfm_5 <= MUX_v_5_2_2(act_read_addrs_sva_2_mx0w0, ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_2_mx0w2,
          and_1276_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_for_and_stg_2_7_sva <= 1'b0;
      Gelu_for_and_2_cse_sva <= 1'b0;
    end
    else if ( ActUnit_PushOutput_if_for_and_28_cse ) begin
      ActUnit_PushOutput_if_for_and_stg_2_7_sva <= MUX1HOT_s_1_4_2(Tanh_for_and_1_cse_sva_mx0w0,
          and_2350_cse, rva_out_reg_data_0_sva_dfm_3, (act_mem_banks_read_read_data_lpi_1_dfm_1_31_0[0]),
          {and_dcpl_331 , and_dcpl_1235 , Tanh_for_or_cse , Tanh_for_and_87_cse});
      Gelu_for_and_2_cse_sva <= MUX1HOT_s_1_3_2(Tanh_for_and_2_cse_sva_mx0w0, rva_out_reg_data_8_sva_dfm_3,
          (act_mem_banks_read_read_data_lpi_1_dfm_1_31_0[8]), {and_dcpl_331 , Tanh_for_or_cse
          , Tanh_for_and_87_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_1_30_26 <= 5'b00000;
    end
    else if ( and_1808_tmp ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_1_30_26 <= MUX1HOT_v_5_5_2(Silu_for_Silu_for_and_19_nl,
          ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_30_26_2,
          nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_121_nl, (act_mem_banks_read_read_data_lpi_1_dfm_1_63_32[20:16]),
          rva_out_reg_data_52_48_sva_dfm_3, {and_dcpl_1112 , and_dcpl_1235 , and_dcpl_1236
          , and_dcpl_1094 , and_dcpl_1096});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_159_128_sva_dfm_3 <= 32'b00000000000000000000000000000000;
      rva_out_reg_data_191_160_sva_dfm_3 <= 32'b00000000000000000000000000000000;
      rva_out_reg_data_223_192_sva_dfm_3 <= 32'b00000000000000000000000000000000;
      rva_out_reg_data_255_224_sva_dfm_3 <= 32'b00000000000000000000000000000000;
      rva_out_reg_data_287_256_sva_dfm_3 <= 32'b00000000000000000000000000000000;
      rva_out_reg_data_319_288_sva_dfm_3 <= 32'b00000000000000000000000000000000;
      rva_out_reg_data_351_320_sva_dfm_3 <= 32'b00000000000000000000000000000000;
      rva_out_reg_data_383_352_sva_dfm_3 <= 32'b00000000000000000000000000000000;
      rva_out_reg_data_415_384_sva_dfm_3 <= 32'b00000000000000000000000000000000;
      rva_out_reg_data_447_416_sva_dfm_3 <= 32'b00000000000000000000000000000000;
      rva_out_reg_data_479_448_sva_dfm_3 <= 32'b00000000000000000000000000000000;
      rva_out_reg_data_511_480_sva_dfm_3 <= 32'b00000000000000000000000000000000;
    end
    else if ( and_1809_cse ) begin
      rva_out_reg_data_159_128_sva_dfm_3 <= MUX_v_32_2_2(ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_13_nl,
          act_mem_banks_read_read_data_lpi_1_dfm_1_159_128, and_dcpl_1094);
      rva_out_reg_data_191_160_sva_dfm_3 <= MUX_v_32_2_2(ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_12_nl,
          act_mem_banks_read_read_data_lpi_1_dfm_1_191_160, and_dcpl_1094);
      rva_out_reg_data_223_192_sva_dfm_3 <= MUX_v_32_2_2(ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_11_nl,
          act_mem_banks_read_read_data_lpi_1_dfm_1_223_192, and_dcpl_1094);
      rva_out_reg_data_255_224_sva_dfm_3 <= MUX_v_32_2_2(ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_10_nl,
          act_mem_banks_read_read_data_lpi_1_dfm_1_255_224, and_dcpl_1094);
      rva_out_reg_data_287_256_sva_dfm_3 <= MUX_v_32_2_2(ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_9_nl,
          act_mem_banks_read_read_data_lpi_1_dfm_1_287_256, and_dcpl_1094);
      rva_out_reg_data_319_288_sva_dfm_3 <= MUX_v_32_2_2(ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_8_nl,
          act_mem_banks_read_read_data_lpi_1_dfm_1_319_288, and_dcpl_1094);
      rva_out_reg_data_351_320_sva_dfm_3 <= MUX_v_32_2_2(ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_7_nl,
          act_mem_banks_read_read_data_lpi_1_dfm_1_351_320, and_dcpl_1094);
      rva_out_reg_data_383_352_sva_dfm_3 <= MUX_v_32_2_2(ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_6_nl,
          act_mem_banks_read_read_data_lpi_1_dfm_1_383_352, and_dcpl_1094);
      rva_out_reg_data_415_384_sva_dfm_3 <= MUX_v_32_2_2(ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_5_nl,
          act_mem_banks_read_read_data_lpi_1_dfm_1_415_384, and_dcpl_1094);
      rva_out_reg_data_447_416_sva_dfm_3 <= MUX_v_32_2_2(ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_4_nl,
          act_mem_banks_read_read_data_lpi_1_dfm_1_447_416, and_dcpl_1094);
      rva_out_reg_data_479_448_sva_dfm_3 <= MUX_v_32_2_2(ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_3_nl,
          act_mem_banks_read_read_data_lpi_1_dfm_1_479_448, and_dcpl_1094);
      rva_out_reg_data_511_480_sva_dfm_3 <= MUX_v_32_2_2(ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_nl,
          act_mem_banks_read_read_data_lpi_1_dfm_1_511_480, and_dcpl_1094);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_31_30_sva_dfm_3 <= 2'b00;
      rva_out_reg_data_103_96_sva_dfm_3 <= 8'b00000000;
      rva_out_reg_data_111_104_sva_dfm_3 <= 8'b00000000;
      rva_out_reg_data_119_112_sva_dfm_3 <= 8'b00000000;
      rva_out_reg_data_127_120_sva_dfm_3 <= 8'b00000000;
      rva_out_reg_data_23_16_sva_dfm_3 <= 8'b00000000;
      rva_out_reg_data_47_40_sva_dfm_3 <= 8'b00000000;
      rva_out_reg_data_63_56_sva_dfm_3 <= 8'b00000000;
      rva_out_reg_data_79_72_sva_dfm_3 <= 8'b00000000;
      rva_out_reg_data_87_80_sva_dfm_3 <= 8'b00000000;
      rva_out_reg_data_95_88_sva_dfm_3 <= 8'b00000000;
      rva_out_reg_data_15_9_sva_dfm_3 <= 7'b0000000;
      rva_out_reg_data_7_1_sva_dfm_3 <= 7'b0000000;
      rva_out_reg_data_55_53_sva_dfm_3 <= 3'b000;
    end
    else if ( rva_out_reg_data_and_15_cse ) begin
      rva_out_reg_data_31_30_sva_dfm_3 <= MUX_v_2_2_2(and_1721_nl, (act_mem_banks_read_read_data_lpi_1_dfm_1_31_0[31:30]),
          and_dcpl_1094);
      rva_out_reg_data_103_96_sva_dfm_3 <= MUX_v_8_2_2(and_1723_nl, (act_mem_banks_read_read_data_lpi_1_dfm_1_127_96[7:0]),
          and_dcpl_1094);
      rva_out_reg_data_111_104_sva_dfm_3 <= MUX_v_8_2_2(and_1725_nl, (act_mem_banks_read_read_data_lpi_1_dfm_1_127_96[15:8]),
          and_dcpl_1094);
      rva_out_reg_data_119_112_sva_dfm_3 <= MUX_v_8_2_2(and_1727_nl, (act_mem_banks_read_read_data_lpi_1_dfm_1_127_96[23:16]),
          and_dcpl_1094);
      rva_out_reg_data_127_120_sva_dfm_3 <= MUX_v_8_2_2(and_1729_nl, (act_mem_banks_read_read_data_lpi_1_dfm_1_127_96[31:24]),
          and_dcpl_1094);
      rva_out_reg_data_23_16_sva_dfm_3 <= MUX_v_8_2_2(and_1731_nl, (act_mem_banks_read_read_data_lpi_1_dfm_1_31_0[23:16]),
          and_dcpl_1094);
      rva_out_reg_data_47_40_sva_dfm_3 <= MUX_v_8_2_2(and_1733_nl, (act_mem_banks_read_read_data_lpi_1_dfm_1_63_32[15:8]),
          and_dcpl_1094);
      rva_out_reg_data_63_56_sva_dfm_3 <= MUX_v_8_2_2(and_1735_nl, (act_mem_banks_read_read_data_lpi_1_dfm_1_63_32[31:24]),
          and_dcpl_1094);
      rva_out_reg_data_79_72_sva_dfm_3 <= MUX_v_8_2_2(and_1737_nl, (act_mem_banks_read_read_data_lpi_1_dfm_1_95_64[15:8]),
          and_dcpl_1094);
      rva_out_reg_data_87_80_sva_dfm_3 <= MUX_v_8_2_2(and_1739_nl, (act_mem_banks_read_read_data_lpi_1_dfm_1_95_64[23:16]),
          and_dcpl_1094);
      rva_out_reg_data_95_88_sva_dfm_3 <= MUX_v_8_2_2(and_1741_nl, (act_mem_banks_read_read_data_lpi_1_dfm_1_95_64[31:24]),
          and_dcpl_1094);
      rva_out_reg_data_15_9_sva_dfm_3 <= MUX_v_7_2_2(and_1743_nl, (act_mem_banks_read_read_data_lpi_1_dfm_1_31_0[15:9]),
          and_dcpl_1094);
      rva_out_reg_data_7_1_sva_dfm_3 <= MUX_v_7_2_2(and_1745_nl, (act_mem_banks_read_read_data_lpi_1_dfm_1_31_0[7:1]),
          and_dcpl_1094);
      rva_out_reg_data_55_53_sva_dfm_3 <= MUX_v_3_2_2(and_1747_nl, (act_mem_banks_read_read_data_lpi_1_dfm_1_63_32[23:21]),
          and_dcpl_1094);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      w_load_lpi_1_dfm_1 <= 1'b0;
    end
    else if ( w_load_and_tmp ) begin
      w_load_lpi_1_dfm_1 <= ~(ActUnit_RunInst_switch_lp_mux_3_nl | ActUnit_RunInst_switch_lp_mux_4_nl
          | ActUnit_RunInst_switch_lp_mux_6_nl | ActUnit_RunInst_switch_lp_mux_8_nl
          | ActUnit_RunInst_switch_lp_mux_10_nl | ActUnit_RunInst_switch_lp_mux_12_nl
          | ActUnit_RunInst_switch_lp_mux_14_nl | ActUnit_RunInst_switch_lp_mux_16_nl
          | ActUnit_RunInst_switch_lp_nor_tmp_mx0);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_RunInst_switch_lp_equal_tmp_2 <= 1'b0;
      ActUnit_RunInst_switch_lp_equal_tmp_4 <= 1'b0;
      ActUnit_RunInst_switch_lp_equal_tmp_5 <= 1'b0;
      ActUnit_RunInst_switch_lp_equal_tmp_6 <= 1'b0;
      ActUnit_RunInst_switch_lp_equal_tmp_7 <= 1'b0;
      ActUnit_RunInst_switch_lp_equal_tmp_8 <= 1'b0;
      Gelu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
          <= 1'b0;
      Gelu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
          <= 1'b0;
      Gelu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
          <= 1'b0;
      Gelu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
          <= 1'b0;
      Gelu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
          <= 1'b0;
      Gelu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
          <= 1'b0;
      Gelu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
          <= 1'b0;
      Gelu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
          <= 1'b0;
    end
    else if ( ActUnit_RunInst_switch_lp_and_802_cse ) begin
      ActUnit_RunInst_switch_lp_equal_tmp_2 <= ActUnit_RunInst_switch_lp_equal_tmp_2_mx0w0;
      ActUnit_RunInst_switch_lp_equal_tmp_4 <= ActUnit_RunInst_switch_lp_equal_tmp_4_mx0w0;
      ActUnit_RunInst_switch_lp_equal_tmp_5 <= ActUnit_RunInst_switch_lp_equal_tmp_5_mx0w0;
      ActUnit_RunInst_switch_lp_equal_tmp_6 <= ActUnit_RunInst_switch_lp_equal_tmp_6_mx0w0;
      ActUnit_RunInst_switch_lp_equal_tmp_7 <= ActUnit_RunInst_switch_lp_equal_tmp_7_mx0w0;
      ActUnit_RunInst_switch_lp_equal_tmp_8 <= ActUnit_RunInst_switch_lp_equal_tmp_8_mx0w0;
      Gelu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
          <= Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs_mx0w0;
      Gelu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
          <= Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs_mx0w0;
      Gelu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
          <= Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs_mx0w0;
      Gelu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
          <= Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs_mx0w0;
      Gelu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
          <= Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs_mx0w0;
      Gelu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
          <= Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs_mx0w0;
      Gelu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
          <= Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs_mx0w0;
      Gelu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
          <= Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_RunInst_switch_lp_equal_tmp_3 <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~(mux_444_nl & (~ (fsm_output[3])))) ) begin
      ActUnit_RunInst_switch_lp_equal_tmp_3 <= ActUnit_RunInst_switch_lp_equal_tmp_3_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= 1'b0;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_ssc ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= MUX_s_1_4_2(act_regs_data_0_15_sva_31, act_regs_data_1_15_sva_31, act_regs_data_2_15_sva_31,
          act_regs_data_3_15_sva_31, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= MUX_s_1_4_2(act_regs_data_0_14_sva_31, act_regs_data_1_14_sva_31, act_regs_data_2_14_sva_31,
          act_regs_data_3_14_sva_31, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= MUX_s_1_4_2(reg_act_regs_data_0_13_ftd, act_regs_data_1_13_sva_31, act_regs_data_2_13_sva_31,
          act_regs_data_3_13_sva_31, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= MUX_s_1_4_2(reg_act_regs_data_0_12_ftd, act_regs_data_1_12_sva_31, act_regs_data_2_12_sva_31,
          act_regs_data_3_12_sva_31, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= MUX_s_1_4_2(reg_act_regs_data_0_11_ftd, act_regs_data_1_11_sva_31, act_regs_data_2_11_sva_31,
          act_regs_data_3_11_sva_31, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= MUX_s_1_4_2(reg_act_regs_data_0_10_ftd, act_regs_data_1_10_sva_31, act_regs_data_2_10_sva_31,
          act_regs_data_3_10_sva_31, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= MUX_s_1_4_2(act_regs_data_0_9_sva_31, act_regs_data_1_9_sva_31, act_regs_data_2_9_sva_31,
          act_regs_data_3_9_sva_31, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= MUX_s_1_4_2(act_regs_data_0_8_sva_31, act_regs_data_1_8_sva_31, act_regs_data_2_8_sva_31,
          act_regs_data_3_8_sva_31, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= MUX_s_1_4_2(act_regs_data_0_7_sva_31, act_regs_data_1_7_sva_31, act_regs_data_2_7_sva_31,
          act_regs_data_3_7_sva_31, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= MUX_s_1_4_2(act_regs_data_0_6_sva_31, act_regs_data_1_6_sva_31, act_regs_data_2_6_sva_31,
          act_regs_data_3_6_sva_31, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= MUX_s_1_4_2(act_regs_data_0_5_sva_31, act_regs_data_1_5_sva_31, act_regs_data_2_5_sva_31,
          act_regs_data_3_5_sva_31, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= MUX_s_1_4_2(act_regs_data_0_4_sva_31, act_regs_data_1_4_sva_31, act_regs_data_2_4_sva_31,
          act_regs_data_3_4_sva_31, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= MUX_s_1_4_2(act_regs_data_0_3_sva_31, act_regs_data_1_3_sva_31, act_regs_data_2_3_sva_31,
          act_regs_data_3_3_sva_31, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= MUX_s_1_4_2(act_regs_data_0_2_sva_31, act_regs_data_1_2_sva_31, act_regs_data_2_2_sva_31,
          act_regs_data_3_2_sva_31, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= MUX_s_1_4_2(reg_act_regs_data_0_1_ftd, act_regs_data_1_1_sva_31, act_regs_data_2_1_sva_31,
          act_regs_data_3_1_sva_31, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31
          <= MUX_s_1_4_2(reg_act_regs_data_0_0_ftd, act_regs_data_1_0_sva_31, act_regs_data_2_0_sva_31,
          act_regs_data_3_0_sva_31, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26
          <= 5'b00000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_37_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26
          <= MUX_v_5_4_2(act_regs_data_0_15_sva_30_26, act_regs_data_1_15_sva_30_26,
          act_regs_data_2_15_sva_30_26, act_regs_data_3_15_sva_30_26, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0
          <= 22'b0000000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_39_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0
          <= MUX_v_22_4_2(act_regs_data_0_15_sva_21_0, act_regs_data_1_15_sva_21_0,
          act_regs_data_2_15_sva_21_0, act_regs_data_3_15_sva_21_0, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26
          <= 5'b00000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_40_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26
          <= MUX_v_5_4_2(act_regs_data_0_14_sva_30_26, act_regs_data_1_14_sva_30_26,
          act_regs_data_2_14_sva_30_26, act_regs_data_3_14_sva_30_26, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0
          <= 22'b0000000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_42_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0
          <= MUX_v_22_4_2(act_regs_data_0_14_sva_21_0, act_regs_data_1_14_sva_21_0,
          act_regs_data_2_14_sva_21_0, act_regs_data_3_14_sva_21_0, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26
          <= 5'b00000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_43_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26
          <= MUX_v_5_4_2(reg_act_regs_data_0_13_ftd_1, act_regs_data_1_13_sva_30_26,
          act_regs_data_2_13_sva_30_26, act_regs_data_3_13_sva_30_26, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0
          <= 22'b0000000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_45_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0
          <= MUX_v_22_4_2(reg_act_regs_data_0_13_ftd_3, act_regs_data_1_13_sva_21_0,
          act_regs_data_2_13_sva_21_0, act_regs_data_3_13_sva_21_0, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26
          <= 5'b00000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_46_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26
          <= MUX_v_5_4_2(reg_act_regs_data_0_12_ftd_1, act_regs_data_1_12_sva_30_26,
          act_regs_data_2_12_sva_30_26, act_regs_data_3_12_sva_30_26, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0
          <= 22'b0000000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_48_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0
          <= MUX_v_22_4_2(reg_act_regs_data_0_12_ftd_3, act_regs_data_1_12_sva_21_0,
          act_regs_data_2_12_sva_21_0, act_regs_data_3_12_sva_21_0, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26
          <= 5'b00000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_49_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26
          <= MUX_v_5_4_2(reg_act_regs_data_0_11_ftd_1, act_regs_data_1_11_sva_30_26,
          act_regs_data_2_11_sva_30_26, act_regs_data_3_11_sva_30_26, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0
          <= 22'b0000000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_51_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0
          <= MUX_v_22_4_2(reg_act_regs_data_0_11_ftd_3, act_regs_data_1_11_sva_21_0,
          act_regs_data_2_11_sva_21_0, act_regs_data_3_11_sva_21_0, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26
          <= 5'b00000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_52_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26
          <= MUX_v_5_4_2(reg_act_regs_data_0_10_ftd_1, act_regs_data_1_10_sva_30_26,
          act_regs_data_2_10_sva_30_26, act_regs_data_3_10_sva_30_26, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0
          <= 22'b0000000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_54_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0
          <= MUX_v_22_4_2(reg_act_regs_data_0_10_ftd_3, act_regs_data_1_10_sva_21_0,
          act_regs_data_2_10_sva_21_0, act_regs_data_3_10_sva_21_0, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26
          <= 5'b00000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_55_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26
          <= MUX_v_5_4_2(act_regs_data_0_9_sva_30_26, act_regs_data_1_9_sva_30_26,
          act_regs_data_2_9_sva_30_26, act_regs_data_3_9_sva_30_26, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0
          <= 22'b0000000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_57_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0
          <= MUX_v_22_4_2(act_regs_data_0_9_sva_21_0, act_regs_data_1_9_sva_21_0,
          act_regs_data_2_9_sva_21_0, act_regs_data_3_9_sva_21_0, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26
          <= 5'b00000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_58_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26
          <= MUX_v_5_4_2(act_regs_data_0_8_sva_30_26, act_regs_data_1_8_sva_30_26,
          act_regs_data_2_8_sva_30_26, act_regs_data_3_8_sva_30_26, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0
          <= 22'b0000000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_60_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0
          <= MUX_v_22_4_2(act_regs_data_0_8_sva_21_0, act_regs_data_1_8_sva_21_0,
          act_regs_data_2_8_sva_21_0, act_regs_data_3_8_sva_21_0, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26
          <= 5'b00000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_61_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26
          <= MUX_v_5_4_2(act_regs_data_0_7_sva_30_26, act_regs_data_1_7_sva_30_26,
          act_regs_data_2_7_sva_30_26, act_regs_data_3_7_sva_30_26, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0
          <= 22'b0000000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_63_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0
          <= MUX_v_22_4_2(act_regs_data_0_7_sva_21_0, act_regs_data_1_7_sva_21_0,
          act_regs_data_2_7_sva_21_0, act_regs_data_3_7_sva_21_0, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26
          <= 5'b00000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_64_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26
          <= MUX_v_5_4_2(act_regs_data_0_6_sva_30_26, act_regs_data_1_6_sva_30_26,
          act_regs_data_2_6_sva_30_26, act_regs_data_3_6_sva_30_26, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0
          <= 22'b0000000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_66_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0
          <= MUX_v_22_4_2(act_regs_data_0_6_sva_21_0, act_regs_data_1_6_sva_21_0,
          act_regs_data_2_6_sva_21_0, act_regs_data_3_6_sva_21_0, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26
          <= 5'b00000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_67_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26
          <= MUX_v_5_4_2(act_regs_data_0_5_sva_30_26, act_regs_data_1_5_sva_30_26,
          act_regs_data_2_5_sva_30_26, act_regs_data_3_5_sva_30_26, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0
          <= 22'b0000000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_69_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0
          <= MUX_v_22_4_2(act_regs_data_0_5_sva_21_0, act_regs_data_1_5_sva_21_0,
          act_regs_data_2_5_sva_21_0, act_regs_data_3_5_sva_21_0, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26
          <= 5'b00000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_70_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26
          <= MUX_v_5_4_2(act_regs_data_0_4_sva_30_26, act_regs_data_1_4_sva_30_26,
          act_regs_data_2_4_sva_30_26, act_regs_data_3_4_sva_30_26, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0
          <= 22'b0000000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_72_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0
          <= MUX_v_22_4_2(act_regs_data_0_4_sva_21_0, act_regs_data_1_4_sva_21_0,
          act_regs_data_2_4_sva_21_0, act_regs_data_3_4_sva_21_0, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26
          <= 5'b00000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_73_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26
          <= MUX_v_5_4_2(act_regs_data_0_3_sva_30_26, act_regs_data_1_3_sva_30_26,
          act_regs_data_2_3_sva_30_26, act_regs_data_3_3_sva_30_26, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0
          <= 22'b0000000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_75_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0
          <= MUX_v_22_4_2(act_regs_data_0_3_sva_21_0, act_regs_data_1_3_sva_21_0,
          act_regs_data_2_3_sva_21_0, act_regs_data_3_3_sva_21_0, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26
          <= 5'b00000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_76_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26
          <= MUX_v_5_4_2(act_regs_data_0_2_sva_30_26, act_regs_data_1_2_sva_30_26,
          act_regs_data_2_2_sva_30_26, act_regs_data_3_2_sva_30_26, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0
          <= 22'b0000000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_78_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0
          <= MUX_v_22_4_2(act_regs_data_0_2_sva_21_0, act_regs_data_1_2_sva_21_0,
          act_regs_data_2_2_sva_21_0, act_regs_data_3_2_sva_21_0, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26
          <= 5'b00000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_79_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26
          <= MUX_v_5_4_2(reg_act_regs_data_0_1_ftd_1, act_regs_data_1_1_sva_30_26,
          act_regs_data_2_1_sva_30_26, act_regs_data_3_1_sva_30_26, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0
          <= 22'b0000000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_81_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0
          <= MUX_v_22_4_2(reg_act_regs_data_0_1_ftd_3, act_regs_data_1_1_sva_21_0,
          act_regs_data_2_1_sva_21_0, act_regs_data_3_1_sva_21_0, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26
          <= 5'b00000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_82_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26
          <= MUX_v_5_4_2(reg_act_regs_data_0_0_ftd_1, act_regs_data_1_0_sva_30_26,
          act_regs_data_2_0_sva_30_26, act_regs_data_3_0_sva_30_26, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0
          <= 22'b0000000000000000000000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_84_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0
          <= MUX_v_22_4_2(reg_act_regs_data_0_0_ftd_3, act_regs_data_1_0_sva_21_0,
          act_regs_data_2_0_sva_21_0, act_regs_data_3_0_sva_21_0, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Tanh_for_y_25_0_lpi_1_dfm_1_ftd <= 1'b0;
      reg_Tanh_for_y_25_0_lpi_1_dfm_1_ftd_1 <= 3'b000;
    end
    else if ( Tanh_for_y_and_31_enex5 ) begin
      reg_Tanh_for_y_25_0_lpi_1_dfm_1_ftd <= (nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          & (~ Tanh_for_and_79_ssc)) | Tanh_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
      reg_Tanh_for_y_25_0_lpi_1_dfm_1_ftd_1 <= MUX_v_3_2_2(nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0,
          3'b100, Tanh_for_or_2_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Tanh_for_y_25_0_lpi_1_dfm_1_21_0 <= 22'b0000000000000000000000;
    end
    else if ( Tanh_for_y_and_32_enex5 ) begin
      Tanh_for_y_25_0_lpi_1_dfm_1_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm,
          Tanh_for_nor_1_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Tanh_for_y_25_0_15_lpi_1_dfm_1_ftd <= 1'b0;
      reg_Tanh_for_y_25_0_15_lpi_1_dfm_1_ftd_1 <= 3'b000;
    end
    else if ( Tanh_for_y_and_33_enex5 ) begin
      reg_Tanh_for_y_25_0_15_lpi_1_dfm_1_ftd <= (nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          & (~ Tanh_for_and_77_ssc)) | Tanh_for_15_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
      reg_Tanh_for_y_25_0_15_lpi_1_dfm_1_ftd_1 <= MUX_v_3_2_2(nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0,
          3'b100, Tanh_for_or_3_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Tanh_for_y_25_0_15_lpi_1_dfm_1_21_0 <= 22'b0000000000000000000000;
    end
    else if ( Tanh_for_y_and_34_enex5 ) begin
      Tanh_for_y_25_0_15_lpi_1_dfm_1_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm,
          Tanh_for_nor_2_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Tanh_for_y_25_0_14_lpi_1_dfm_1_ftd <= 1'b0;
      reg_Tanh_for_y_25_0_14_lpi_1_dfm_1_ftd_1 <= 3'b000;
    end
    else if ( Tanh_for_y_and_35_enex5 ) begin
      reg_Tanh_for_y_25_0_14_lpi_1_dfm_1_ftd <= (nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          & (~ Tanh_for_and_75_ssc)) | Tanh_for_14_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
      reg_Tanh_for_y_25_0_14_lpi_1_dfm_1_ftd_1 <= MUX_v_3_2_2(nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0,
          3'b100, Tanh_for_or_4_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Tanh_for_y_25_0_14_lpi_1_dfm_1_21_0 <= 22'b0000000000000000000000;
    end
    else if ( Tanh_for_y_and_36_enex5 ) begin
      Tanh_for_y_25_0_14_lpi_1_dfm_1_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm,
          Tanh_for_nor_3_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Tanh_for_y_25_0_13_lpi_1_dfm_1_ftd <= 1'b0;
      reg_Tanh_for_y_25_0_13_lpi_1_dfm_1_ftd_1 <= 3'b000;
    end
    else if ( Tanh_for_y_and_37_enex5 ) begin
      reg_Tanh_for_y_25_0_13_lpi_1_dfm_1_ftd <= (nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          & (~ Tanh_for_and_73_ssc)) | Tanh_for_13_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
      reg_Tanh_for_y_25_0_13_lpi_1_dfm_1_ftd_1 <= MUX_v_3_2_2(nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0,
          3'b100, Tanh_for_or_5_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Tanh_for_y_25_0_13_lpi_1_dfm_1_21_0 <= 22'b0000000000000000000000;
    end
    else if ( Tanh_for_y_and_38_enex5 ) begin
      Tanh_for_y_25_0_13_lpi_1_dfm_1_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm,
          Tanh_for_nor_4_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Tanh_for_y_25_0_12_lpi_1_dfm_1_ftd <= 1'b0;
      reg_Tanh_for_y_25_0_12_lpi_1_dfm_1_ftd_1 <= 3'b000;
    end
    else if ( Tanh_for_y_and_39_enex5 ) begin
      reg_Tanh_for_y_25_0_12_lpi_1_dfm_1_ftd <= (nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          & (~ Tanh_for_and_71_ssc)) | Tanh_for_12_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
      reg_Tanh_for_y_25_0_12_lpi_1_dfm_1_ftd_1 <= MUX_v_3_2_2(nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0,
          3'b100, Tanh_for_or_6_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Tanh_for_y_25_0_12_lpi_1_dfm_1_21_0 <= 22'b0000000000000000000000;
    end
    else if ( Tanh_for_y_and_40_enex5 ) begin
      Tanh_for_y_25_0_12_lpi_1_dfm_1_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm,
          Tanh_for_nor_5_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Tanh_for_y_25_0_11_lpi_1_dfm_1_ftd <= 1'b0;
      reg_Tanh_for_y_25_0_11_lpi_1_dfm_1_ftd_1 <= 3'b000;
    end
    else if ( Tanh_for_y_and_41_enex5 ) begin
      reg_Tanh_for_y_25_0_11_lpi_1_dfm_1_ftd <= (nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          & (~ Tanh_for_and_69_ssc)) | Tanh_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
      reg_Tanh_for_y_25_0_11_lpi_1_dfm_1_ftd_1 <= MUX_v_3_2_2(nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0,
          3'b100, Tanh_for_or_7_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Tanh_for_y_25_0_11_lpi_1_dfm_1_21_0 <= 22'b0000000000000000000000;
    end
    else if ( Tanh_for_y_and_42_enex5 ) begin
      Tanh_for_y_25_0_11_lpi_1_dfm_1_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm,
          Tanh_for_nor_6_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Tanh_for_y_25_0_10_lpi_1_dfm_1_ftd <= 1'b0;
      reg_Tanh_for_y_25_0_10_lpi_1_dfm_1_ftd_1 <= 3'b000;
    end
    else if ( Tanh_for_y_and_43_enex5 ) begin
      reg_Tanh_for_y_25_0_10_lpi_1_dfm_1_ftd <= (nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          & (~ Tanh_for_and_67_ssc)) | Tanh_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
      reg_Tanh_for_y_25_0_10_lpi_1_dfm_1_ftd_1 <= MUX_v_3_2_2(nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0,
          3'b100, Tanh_for_or_8_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Tanh_for_y_25_0_10_lpi_1_dfm_1_21_0 <= 22'b0000000000000000000000;
    end
    else if ( Tanh_for_y_and_44_enex5 ) begin
      Tanh_for_y_25_0_10_lpi_1_dfm_1_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm,
          Tanh_for_nor_7_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Tanh_for_y_25_0_9_lpi_1_dfm_1_ftd <= 1'b0;
      reg_Tanh_for_y_25_0_9_lpi_1_dfm_1_ftd_1 <= 3'b000;
    end
    else if ( Tanh_for_y_and_45_enex5 ) begin
      reg_Tanh_for_y_25_0_9_lpi_1_dfm_1_ftd <= (nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          & (~ Tanh_for_and_65_ssc)) | Tanh_for_9_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
      reg_Tanh_for_y_25_0_9_lpi_1_dfm_1_ftd_1 <= MUX_v_3_2_2(nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0,
          3'b100, Tanh_for_or_9_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Tanh_for_y_25_0_9_lpi_1_dfm_1_21_0 <= 22'b0000000000000000000000;
    end
    else if ( Tanh_for_y_and_46_enex5 ) begin
      Tanh_for_y_25_0_9_lpi_1_dfm_1_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm,
          Tanh_for_nor_8_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Tanh_for_y_25_0_8_lpi_1_dfm_1_ftd <= 1'b0;
      reg_Tanh_for_y_25_0_8_lpi_1_dfm_1_ftd_1 <= 3'b000;
    end
    else if ( Tanh_for_y_and_47_enex5 ) begin
      reg_Tanh_for_y_25_0_8_lpi_1_dfm_1_ftd <= (nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          & (~ Tanh_for_and_63_ssc)) | Tanh_for_8_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
      reg_Tanh_for_y_25_0_8_lpi_1_dfm_1_ftd_1 <= MUX_v_3_2_2(nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0,
          3'b100, Tanh_for_or_10_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Tanh_for_y_25_0_8_lpi_1_dfm_1_21_0 <= 22'b0000000000000000000000;
    end
    else if ( Tanh_for_y_and_48_enex5 ) begin
      Tanh_for_y_25_0_8_lpi_1_dfm_1_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm,
          Tanh_for_nor_9_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Tanh_for_y_25_0_7_lpi_1_dfm_1_ftd <= 1'b0;
      reg_Tanh_for_y_25_0_7_lpi_1_dfm_1_ftd_1 <= 3'b000;
    end
    else if ( Tanh_for_y_and_49_enex5 ) begin
      reg_Tanh_for_y_25_0_7_lpi_1_dfm_1_ftd <= (nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          & (~ Tanh_for_and_61_ssc)) | Tanh_for_7_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
      reg_Tanh_for_y_25_0_7_lpi_1_dfm_1_ftd_1 <= MUX_v_3_2_2(nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0,
          3'b100, Tanh_for_or_11_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Tanh_for_y_25_0_7_lpi_1_dfm_1_21_0 <= 22'b0000000000000000000000;
    end
    else if ( Tanh_for_y_and_50_enex5 ) begin
      Tanh_for_y_25_0_7_lpi_1_dfm_1_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm,
          Tanh_for_nor_10_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Tanh_for_y_25_0_6_lpi_1_dfm_1_ftd <= 1'b0;
      reg_Tanh_for_y_25_0_6_lpi_1_dfm_1_ftd_1 <= 3'b000;
    end
    else if ( Tanh_for_y_and_51_enex5 ) begin
      reg_Tanh_for_y_25_0_6_lpi_1_dfm_1_ftd <= (nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          & (~ Tanh_for_and_59_ssc)) | Tanh_for_6_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
      reg_Tanh_for_y_25_0_6_lpi_1_dfm_1_ftd_1 <= MUX_v_3_2_2(nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0,
          3'b100, Tanh_for_or_12_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Tanh_for_y_25_0_6_lpi_1_dfm_1_21_0 <= 22'b0000000000000000000000;
    end
    else if ( Tanh_for_y_and_52_enex5 ) begin
      Tanh_for_y_25_0_6_lpi_1_dfm_1_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm,
          Tanh_for_nor_11_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Tanh_for_y_25_0_5_lpi_1_dfm_1_ftd <= 1'b0;
      reg_Tanh_for_y_25_0_5_lpi_1_dfm_1_ftd_1 <= 3'b000;
    end
    else if ( Tanh_for_y_and_53_enex5 ) begin
      reg_Tanh_for_y_25_0_5_lpi_1_dfm_1_ftd <= (nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          & (~ Tanh_for_and_57_ssc)) | Tanh_for_5_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
      reg_Tanh_for_y_25_0_5_lpi_1_dfm_1_ftd_1 <= MUX_v_3_2_2(nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0,
          3'b100, Tanh_for_or_13_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Tanh_for_y_25_0_5_lpi_1_dfm_1_21_0 <= 22'b0000000000000000000000;
    end
    else if ( Tanh_for_y_and_54_enex5 ) begin
      Tanh_for_y_25_0_5_lpi_1_dfm_1_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm,
          Tanh_for_nor_12_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Tanh_for_y_25_0_4_lpi_1_dfm_1_ftd <= 1'b0;
      reg_Tanh_for_y_25_0_4_lpi_1_dfm_1_ftd_1 <= 3'b000;
    end
    else if ( Tanh_for_y_and_55_enex5 ) begin
      reg_Tanh_for_y_25_0_4_lpi_1_dfm_1_ftd <= (nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          & (~ Tanh_for_and_55_ssc)) | Tanh_for_4_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
      reg_Tanh_for_y_25_0_4_lpi_1_dfm_1_ftd_1 <= MUX_v_3_2_2(nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0,
          3'b100, Tanh_for_or_14_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Tanh_for_y_25_0_4_lpi_1_dfm_1_21_0 <= 22'b0000000000000000000000;
    end
    else if ( Tanh_for_y_and_56_enex5 ) begin
      Tanh_for_y_25_0_4_lpi_1_dfm_1_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm,
          Tanh_for_nor_13_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Tanh_for_y_25_0_3_lpi_1_dfm_1_ftd <= 1'b0;
      reg_Tanh_for_y_25_0_3_lpi_1_dfm_1_ftd_1 <= 3'b000;
    end
    else if ( Tanh_for_y_and_57_enex5 ) begin
      reg_Tanh_for_y_25_0_3_lpi_1_dfm_1_ftd <= (nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          & (~ Tanh_for_and_53_ssc)) | Tanh_for_3_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
      reg_Tanh_for_y_25_0_3_lpi_1_dfm_1_ftd_1 <= MUX_v_3_2_2(nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0,
          3'b100, Tanh_for_or_15_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Tanh_for_y_25_0_3_lpi_1_dfm_1_21_0 <= 22'b0000000000000000000000;
    end
    else if ( Tanh_for_y_and_58_enex5 ) begin
      Tanh_for_y_25_0_3_lpi_1_dfm_1_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm,
          Tanh_for_nor_14_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Tanh_for_y_25_0_2_lpi_1_dfm_1_ftd <= 1'b0;
      reg_Tanh_for_y_25_0_2_lpi_1_dfm_1_ftd_1 <= 3'b000;
    end
    else if ( Tanh_for_y_and_59_enex5 ) begin
      reg_Tanh_for_y_25_0_2_lpi_1_dfm_1_ftd <= (nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          & (~ Tanh_for_and_51_ssc)) | Tanh_for_2_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
      reg_Tanh_for_y_25_0_2_lpi_1_dfm_1_ftd_1 <= MUX_v_3_2_2(nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0,
          3'b100, Tanh_for_or_16_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Tanh_for_y_25_0_2_lpi_1_dfm_1_21_0 <= 22'b0000000000000000000000;
    end
    else if ( Tanh_for_y_and_60_enex5 ) begin
      Tanh_for_y_25_0_2_lpi_1_dfm_1_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm,
          Tanh_for_nor_15_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Tanh_for_y_25_0_1_lpi_1_dfm_1_ftd <= 1'b0;
      reg_Tanh_for_y_25_0_1_lpi_1_dfm_1_ftd_1 <= 3'b000;
    end
    else if ( Tanh_for_y_and_61_enex5 ) begin
      reg_Tanh_for_y_25_0_1_lpi_1_dfm_1_ftd <= (nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          & (~ Tanh_for_and_49_ssc)) | Tanh_for_1_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
      reg_Tanh_for_y_25_0_1_lpi_1_dfm_1_ftd_1 <= MUX_v_3_2_2(nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0,
          3'b100, Tanh_for_or_17_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Tanh_for_y_25_0_1_lpi_1_dfm_1_21_0 <= 22'b0000000000000000000000;
    end
    else if ( Tanh_for_y_and_62_enex5 ) begin
      Tanh_for_y_25_0_1_lpi_1_dfm_1_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm,
          Tanh_for_nor_16_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_lpi_1_dfm_30_26 <= 5'b00000;
    end
    else if ( Relu_for_y_qelse_and_31_enex5 ) begin
      Relu_for_y_qr_30_0_lpi_1_dfm_30_26 <= MUX_v_5_2_2(5'b00000, nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm,
          nv_scvector_cctor_nv_scvector_4_for_not_43_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_lpi_1_dfm_25 <= 1'b0;
      Relu_for_y_qr_30_0_lpi_1_dfm_24_22 <= 3'b000;
    end
    else if ( Relu_for_y_qelse_and_32_enex5 ) begin
      Relu_for_y_qr_30_0_lpi_1_dfm_25 <= nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          & (~ nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm);
      Relu_for_y_qr_30_0_lpi_1_dfm_24_22 <= MUX_v_3_2_2(3'b000, nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0,
          nv_scvector_cctor_nv_scvector_4_for_not_59_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_lpi_1_dfm_21_0 <= 22'b0000000000000000000000;
    end
    else if ( Relu_for_y_qelse_and_33_enex5 ) begin
      Relu_for_y_qr_30_0_lpi_1_dfm_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm,
          nv_scvector_cctor_nv_scvector_4_for_not_14_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_15_lpi_1_dfm_30_26 <= 5'b00000;
    end
    else if ( Relu_for_y_qelse_and_34_enex5 ) begin
      Relu_for_y_qr_30_0_15_lpi_1_dfm_30_26 <= MUX_v_5_2_2(5'b00000, nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm,
          nv_scvector_cctor_nv_scvector_4_for_not_41_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_15_lpi_1_dfm_25 <= 1'b0;
      Relu_for_y_qr_30_0_15_lpi_1_dfm_24_22 <= 3'b000;
    end
    else if ( Relu_for_y_qelse_and_35_enex5 ) begin
      Relu_for_y_qr_30_0_15_lpi_1_dfm_25 <= nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          & (~ nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm);
      Relu_for_y_qr_30_0_15_lpi_1_dfm_24_22 <= MUX_v_3_2_2(3'b000, nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0,
          nv_scvector_cctor_nv_scvector_4_for_not_58_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_15_lpi_1_dfm_21_0 <= 22'b0000000000000000000000;
    end
    else if ( Relu_for_y_qelse_and_36_enex5 ) begin
      Relu_for_y_qr_30_0_15_lpi_1_dfm_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm,
          nv_scvector_cctor_nv_scvector_4_for_not_13_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_14_lpi_1_dfm_30_26 <= 5'b00000;
    end
    else if ( Relu_for_y_qelse_and_37_enex5 ) begin
      Relu_for_y_qr_30_0_14_lpi_1_dfm_30_26 <= MUX_v_5_2_2(5'b00000, nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm,
          nv_scvector_cctor_nv_scvector_4_for_not_39_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_14_lpi_1_dfm_25 <= 1'b0;
      Relu_for_y_qr_30_0_14_lpi_1_dfm_24_22 <= 3'b000;
    end
    else if ( Relu_for_y_qelse_and_38_enex5 ) begin
      Relu_for_y_qr_30_0_14_lpi_1_dfm_25 <= nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          & (~ nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm);
      Relu_for_y_qr_30_0_14_lpi_1_dfm_24_22 <= MUX_v_3_2_2(3'b000, nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0,
          nv_scvector_cctor_nv_scvector_4_for_not_57_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_14_lpi_1_dfm_21_0 <= 22'b0000000000000000000000;
    end
    else if ( Relu_for_y_qelse_and_39_enex5 ) begin
      Relu_for_y_qr_30_0_14_lpi_1_dfm_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm,
          nv_scvector_cctor_nv_scvector_4_for_not_12_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_13_lpi_1_dfm_30_26 <= 5'b00000;
    end
    else if ( Relu_for_y_qelse_and_40_enex5 ) begin
      Relu_for_y_qr_30_0_13_lpi_1_dfm_30_26 <= MUX_v_5_2_2(5'b00000, nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm,
          nv_scvector_cctor_nv_scvector_4_for_not_37_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_13_lpi_1_dfm_25 <= 1'b0;
      Relu_for_y_qr_30_0_13_lpi_1_dfm_24_22 <= 3'b000;
    end
    else if ( Relu_for_y_qelse_and_41_enex5 ) begin
      Relu_for_y_qr_30_0_13_lpi_1_dfm_25 <= nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          & (~ nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm);
      Relu_for_y_qr_30_0_13_lpi_1_dfm_24_22 <= MUX_v_3_2_2(3'b000, nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0,
          nv_scvector_cctor_nv_scvector_4_for_not_56_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_13_lpi_1_dfm_21_0 <= 22'b0000000000000000000000;
    end
    else if ( Relu_for_y_qelse_and_42_enex5 ) begin
      Relu_for_y_qr_30_0_13_lpi_1_dfm_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm,
          nv_scvector_cctor_nv_scvector_4_for_not_11_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_12_lpi_1_dfm_30_26 <= 5'b00000;
    end
    else if ( Relu_for_y_qelse_and_43_enex5 ) begin
      Relu_for_y_qr_30_0_12_lpi_1_dfm_30_26 <= MUX_v_5_2_2(5'b00000, nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm,
          nv_scvector_cctor_nv_scvector_4_for_not_35_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_12_lpi_1_dfm_25 <= 1'b0;
      Relu_for_y_qr_30_0_12_lpi_1_dfm_24_22 <= 3'b000;
    end
    else if ( Relu_for_y_qelse_and_44_enex5 ) begin
      Relu_for_y_qr_30_0_12_lpi_1_dfm_25 <= nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          & (~ nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm);
      Relu_for_y_qr_30_0_12_lpi_1_dfm_24_22 <= MUX_v_3_2_2(3'b000, nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0,
          nv_scvector_cctor_nv_scvector_4_for_not_55_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_12_lpi_1_dfm_21_0 <= 22'b0000000000000000000000;
    end
    else if ( Relu_for_y_qelse_and_45_enex5 ) begin
      Relu_for_y_qr_30_0_12_lpi_1_dfm_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm,
          nv_scvector_cctor_nv_scvector_4_for_not_10_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_11_lpi_1_dfm_30_26 <= 5'b00000;
    end
    else if ( Relu_for_y_qelse_and_46_enex5 ) begin
      Relu_for_y_qr_30_0_11_lpi_1_dfm_30_26 <= MUX_v_5_2_2(5'b00000, nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm,
          nv_scvector_cctor_nv_scvector_4_for_not_33_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_11_lpi_1_dfm_25 <= 1'b0;
      Relu_for_y_qr_30_0_11_lpi_1_dfm_24_22 <= 3'b000;
    end
    else if ( Relu_for_y_qelse_and_47_enex5 ) begin
      Relu_for_y_qr_30_0_11_lpi_1_dfm_25 <= nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          & (~ nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm);
      Relu_for_y_qr_30_0_11_lpi_1_dfm_24_22 <= MUX_v_3_2_2(3'b000, nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0,
          nv_scvector_cctor_nv_scvector_4_for_not_54_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_11_lpi_1_dfm_21_0 <= 22'b0000000000000000000000;
    end
    else if ( Relu_for_y_qelse_and_48_enex5 ) begin
      Relu_for_y_qr_30_0_11_lpi_1_dfm_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm,
          nv_scvector_cctor_nv_scvector_4_for_not_9_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_10_lpi_1_dfm_30_26 <= 5'b00000;
    end
    else if ( Relu_for_y_qelse_and_49_enex5 ) begin
      Relu_for_y_qr_30_0_10_lpi_1_dfm_30_26 <= MUX_v_5_2_2(5'b00000, nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm,
          nv_scvector_cctor_nv_scvector_4_for_not_31_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_10_lpi_1_dfm_25 <= 1'b0;
      Relu_for_y_qr_30_0_10_lpi_1_dfm_24_22 <= 3'b000;
    end
    else if ( Relu_for_y_qelse_and_50_enex5 ) begin
      Relu_for_y_qr_30_0_10_lpi_1_dfm_25 <= nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          & (~ nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm);
      Relu_for_y_qr_30_0_10_lpi_1_dfm_24_22 <= MUX_v_3_2_2(3'b000, nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0,
          nv_scvector_cctor_nv_scvector_4_for_not_53_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_10_lpi_1_dfm_21_0 <= 22'b0000000000000000000000;
    end
    else if ( Relu_for_y_qelse_and_51_enex5 ) begin
      Relu_for_y_qr_30_0_10_lpi_1_dfm_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm,
          nv_scvector_cctor_nv_scvector_4_for_not_8_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_9_lpi_1_dfm_30_26 <= 5'b00000;
    end
    else if ( Relu_for_y_qelse_and_52_enex5 ) begin
      Relu_for_y_qr_30_0_9_lpi_1_dfm_30_26 <= MUX_v_5_2_2(5'b00000, nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm,
          nv_scvector_cctor_nv_scvector_4_for_not_29_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_9_lpi_1_dfm_25 <= 1'b0;
      Relu_for_y_qr_30_0_9_lpi_1_dfm_24_22 <= 3'b000;
    end
    else if ( Relu_for_y_qelse_and_53_enex5 ) begin
      Relu_for_y_qr_30_0_9_lpi_1_dfm_25 <= nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          & (~ nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm);
      Relu_for_y_qr_30_0_9_lpi_1_dfm_24_22 <= MUX_v_3_2_2(3'b000, nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0,
          nv_scvector_cctor_nv_scvector_4_for_not_52_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_9_lpi_1_dfm_21_0 <= 22'b0000000000000000000000;
    end
    else if ( Relu_for_y_qelse_and_54_enex5 ) begin
      Relu_for_y_qr_30_0_9_lpi_1_dfm_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm,
          nv_scvector_cctor_nv_scvector_4_for_not_7_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_8_lpi_1_dfm_30_26 <= 5'b00000;
    end
    else if ( Relu_for_y_qelse_and_55_enex5 ) begin
      Relu_for_y_qr_30_0_8_lpi_1_dfm_30_26 <= MUX_v_5_2_2(5'b00000, nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm,
          nv_scvector_cctor_nv_scvector_4_for_not_27_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_8_lpi_1_dfm_25 <= 1'b0;
      Relu_for_y_qr_30_0_8_lpi_1_dfm_24_22 <= 3'b000;
    end
    else if ( Relu_for_y_qelse_and_56_enex5 ) begin
      Relu_for_y_qr_30_0_8_lpi_1_dfm_25 <= nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          & (~ nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm);
      Relu_for_y_qr_30_0_8_lpi_1_dfm_24_22 <= MUX_v_3_2_2(3'b000, nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0,
          nv_scvector_cctor_nv_scvector_4_for_not_51_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_8_lpi_1_dfm_21_0 <= 22'b0000000000000000000000;
    end
    else if ( Relu_for_y_qelse_and_57_enex5 ) begin
      Relu_for_y_qr_30_0_8_lpi_1_dfm_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm,
          nv_scvector_cctor_nv_scvector_4_for_not_6_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_7_lpi_1_dfm_30_26 <= 5'b00000;
    end
    else if ( Relu_for_y_qelse_and_58_enex5 ) begin
      Relu_for_y_qr_30_0_7_lpi_1_dfm_30_26 <= MUX_v_5_2_2(5'b00000, nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm,
          nv_scvector_cctor_nv_scvector_4_for_not_25_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_7_lpi_1_dfm_25 <= 1'b0;
      Relu_for_y_qr_30_0_7_lpi_1_dfm_24_22 <= 3'b000;
    end
    else if ( Relu_for_y_qelse_and_59_enex5 ) begin
      Relu_for_y_qr_30_0_7_lpi_1_dfm_25 <= nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          & (~ nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm);
      Relu_for_y_qr_30_0_7_lpi_1_dfm_24_22 <= MUX_v_3_2_2(3'b000, nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0,
          nv_scvector_cctor_nv_scvector_4_for_not_50_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_7_lpi_1_dfm_21_0 <= 22'b0000000000000000000000;
    end
    else if ( Relu_for_y_qelse_and_60_enex5 ) begin
      Relu_for_y_qr_30_0_7_lpi_1_dfm_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm,
          nv_scvector_cctor_nv_scvector_4_for_not_5_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_6_lpi_1_dfm_30_26 <= 5'b00000;
    end
    else if ( Relu_for_y_qelse_and_61_enex5 ) begin
      Relu_for_y_qr_30_0_6_lpi_1_dfm_30_26 <= MUX_v_5_2_2(5'b00000, nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm,
          nv_scvector_cctor_nv_scvector_4_for_not_23_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_6_lpi_1_dfm_25 <= 1'b0;
      Relu_for_y_qr_30_0_6_lpi_1_dfm_24_22 <= 3'b000;
    end
    else if ( Relu_for_y_qelse_and_62_enex5 ) begin
      Relu_for_y_qr_30_0_6_lpi_1_dfm_25 <= nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          & (~ nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm);
      Relu_for_y_qr_30_0_6_lpi_1_dfm_24_22 <= MUX_v_3_2_2(3'b000, nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0,
          nv_scvector_cctor_nv_scvector_4_for_not_49_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_6_lpi_1_dfm_21_0 <= 22'b0000000000000000000000;
    end
    else if ( Relu_for_y_qelse_and_63_enex5 ) begin
      Relu_for_y_qr_30_0_6_lpi_1_dfm_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm,
          nv_scvector_cctor_nv_scvector_4_for_not_4_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_5_lpi_1_dfm_30_26 <= 5'b00000;
    end
    else if ( Relu_for_y_qelse_and_64_enex5 ) begin
      Relu_for_y_qr_30_0_5_lpi_1_dfm_30_26 <= MUX_v_5_2_2(5'b00000, nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm,
          nv_scvector_cctor_nv_scvector_4_for_not_21_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_5_lpi_1_dfm_25 <= 1'b0;
      Relu_for_y_qr_30_0_5_lpi_1_dfm_24_22 <= 3'b000;
    end
    else if ( Relu_for_y_qelse_and_65_enex5 ) begin
      Relu_for_y_qr_30_0_5_lpi_1_dfm_25 <= nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          & (~ nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm);
      Relu_for_y_qr_30_0_5_lpi_1_dfm_24_22 <= MUX_v_3_2_2(3'b000, nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0,
          nv_scvector_cctor_nv_scvector_4_for_not_48_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_5_lpi_1_dfm_21_0 <= 22'b0000000000000000000000;
    end
    else if ( Relu_for_y_qelse_and_66_enex5 ) begin
      Relu_for_y_qr_30_0_5_lpi_1_dfm_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm,
          nv_scvector_cctor_nv_scvector_4_for_not_3_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_4_lpi_1_dfm_30_26 <= 5'b00000;
    end
    else if ( Relu_for_y_qelse_and_67_enex5 ) begin
      Relu_for_y_qr_30_0_4_lpi_1_dfm_30_26 <= MUX_v_5_2_2(5'b00000, nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm,
          nv_scvector_cctor_nv_scvector_4_for_not_19_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_4_lpi_1_dfm_25 <= 1'b0;
      Relu_for_y_qr_30_0_4_lpi_1_dfm_24_22 <= 3'b000;
    end
    else if ( Relu_for_y_qelse_and_68_enex5 ) begin
      Relu_for_y_qr_30_0_4_lpi_1_dfm_25 <= nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          & (~ nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm);
      Relu_for_y_qr_30_0_4_lpi_1_dfm_24_22 <= MUX_v_3_2_2(3'b000, nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0,
          nv_scvector_cctor_nv_scvector_4_for_not_47_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_4_lpi_1_dfm_21_0 <= 22'b0000000000000000000000;
    end
    else if ( Relu_for_y_qelse_and_69_enex5 ) begin
      Relu_for_y_qr_30_0_4_lpi_1_dfm_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm,
          nv_scvector_cctor_nv_scvector_4_for_not_2_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_3_lpi_1_dfm_30_26 <= 5'b00000;
    end
    else if ( Relu_for_y_qelse_and_70_enex5 ) begin
      Relu_for_y_qr_30_0_3_lpi_1_dfm_30_26 <= MUX_v_5_2_2(5'b00000, nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm,
          nv_scvector_cctor_nv_scvector_4_for_not_17_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_3_lpi_1_dfm_25 <= 1'b0;
      Relu_for_y_qr_30_0_3_lpi_1_dfm_24_22 <= 3'b000;
    end
    else if ( Relu_for_y_qelse_and_71_enex5 ) begin
      Relu_for_y_qr_30_0_3_lpi_1_dfm_25 <= nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          & (~ nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm);
      Relu_for_y_qr_30_0_3_lpi_1_dfm_24_22 <= MUX_v_3_2_2(3'b000, nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0,
          nv_scvector_cctor_nv_scvector_4_for_not_46_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_3_lpi_1_dfm_21_0 <= 22'b0000000000000000000000;
    end
    else if ( Relu_for_y_qelse_and_72_enex5 ) begin
      Relu_for_y_qr_30_0_3_lpi_1_dfm_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm,
          nv_scvector_cctor_nv_scvector_4_for_not_1_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_2_lpi_1_dfm_30_26 <= 5'b00000;
    end
    else if ( Relu_for_y_qelse_and_73_enex5 ) begin
      Relu_for_y_qr_30_0_2_lpi_1_dfm_30_26 <= MUX_v_5_2_2(5'b00000, nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm,
          nv_scvector_cctor_nv_scvector_4_for_not_15_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_2_lpi_1_dfm_25 <= 1'b0;
      Relu_for_y_qr_30_0_2_lpi_1_dfm_24_22 <= 3'b000;
    end
    else if ( Relu_for_y_qelse_and_74_enex5 ) begin
      Relu_for_y_qr_30_0_2_lpi_1_dfm_25 <= nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          & (~ nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm);
      Relu_for_y_qr_30_0_2_lpi_1_dfm_24_22 <= MUX_v_3_2_2(3'b000, nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0,
          nv_scvector_cctor_nv_scvector_4_for_not_45_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_2_lpi_1_dfm_21_0 <= 22'b0000000000000000000000;
    end
    else if ( Relu_for_y_qelse_and_75_enex5 ) begin
      Relu_for_y_qr_30_0_2_lpi_1_dfm_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm,
          nv_scvector_cctor_nv_scvector_4_for_not_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_1_lpi_1_dfm_30_26 <= 5'b00000;
    end
    else if ( Relu_for_y_qelse_and_76_enex5 ) begin
      Relu_for_y_qr_30_0_1_lpi_1_dfm_30_26 <= MUX_v_5_2_2(5'b00000, nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm,
          ActUnit_RunInst_switch_lp_not_10_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_1_lpi_1_dfm_25 <= 1'b0;
      Relu_for_y_qr_30_0_1_lpi_1_dfm_24_22 <= 3'b000;
    end
    else if ( Relu_for_y_qelse_and_77_enex5 ) begin
      Relu_for_y_qr_30_0_1_lpi_1_dfm_25 <= nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          & (~ nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm);
      Relu_for_y_qr_30_0_1_lpi_1_dfm_24_22 <= MUX_v_3_2_2(3'b000, nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0,
          ActUnit_RunInst_switch_lp_not_12_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Relu_for_y_qr_30_0_1_lpi_1_dfm_21_0 <= 22'b0000000000000000000000;
    end
    else if ( Relu_for_y_qelse_and_78_enex5 ) begin
      Relu_for_y_qr_30_0_1_lpi_1_dfm_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm,
          ActUnit_RunInst_switch_lp_not_1_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= 1'b0;
      Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= 1'b0;
      Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= 1'b0;
      Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= 1'b0;
      Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= 1'b0;
      Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= 1'b0;
      Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= 1'b0;
      Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= 1'b0;
    end
    else if ( operator_32_8_true_AC_TRN_AC_WRAP_2_and_cse ) begin
      Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs_mx0w0;
      Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs_mx0w0;
      Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs_mx0w0;
      Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs_mx0w0;
      Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs_mx0w0;
      Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs_mx0w0;
      Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs_mx0w0;
      Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs_mx0w0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= 1'b0;
      Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= 1'b0;
      Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= 1'b0;
      Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= 1'b0;
      Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= 1'b0;
      Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= 1'b0;
      Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= 1'b0;
      Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= 1'b0;
    end
    else if ( operator_32_8_true_AC_TRN_AC_WRAP_2_and_16_cse ) begin
      Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= $signed(1'b0) < $signed(({nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
          , nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
          , nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          , nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
          , nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
      Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= $signed(1'b0) < $signed(({nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
          , nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
          , nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          , nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
          , nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
      Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= $signed(1'b0) < $signed(({nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
          , nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
          , nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          , nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
          , nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
      Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= $signed(1'b0) < $signed(({nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
          , nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
          , nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          , nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
          , nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
      Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= $signed(1'b0) < $signed(({nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
          , nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
          , nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          , nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
          , nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
      Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= $signed(1'b0) < $signed(({nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
          , nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
          , nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          , nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
          , nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
      Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= $signed(1'b0) < $signed(({nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
          , nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
          , nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          , nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
          , nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
      Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
          <= $signed(1'b0) < $signed(({nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm
          , nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm
          , nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3
          , nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0
          , nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm}));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_config_in_InstFetch_return_sva_7_2 <= 6'b000000;
    end
    else if ( ActUnit_RunInst_curr_inst_and_enex5 ) begin
      act_config_in_InstFetch_return_sva_7_2 <= act_config_in_InstFetch_mux_tmp[7:2];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= 1'b0;
      Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= 1'b0;
      Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= 1'b0;
      Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= 1'b0;
      Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= 1'b0;
      Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= 1'b0;
      Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= 1'b0;
      Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= 1'b0;
    end
    else if ( operator_32_8_true_AC_TRN_AC_WRAP_and_cse ) begin
      Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_less_tmp;
      Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_less_1_tmp;
      Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_less_2_tmp;
      Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_less_3_tmp;
      Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_less_4_tmp;
      Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_less_5_tmp;
      Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_less_6_tmp;
      Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_less_7_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= 1'b0;
      Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= 1'b0;
      Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= 1'b0;
      Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= 1'b0;
      Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= 1'b0;
      Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= 1'b0;
      Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= 1'b0;
      Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= 1'b0;
    end
    else if ( operator_32_8_true_AC_TRN_AC_WRAP_and_23_cse ) begin
      Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_less_8_tmp;
      Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_less_9_tmp;
      Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_less_10_tmp;
      Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_less_11_tmp;
      Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_less_12_tmp;
      Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_less_13_tmp;
      Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_less_14_tmp;
      Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
          <= operator_32_8_true_AC_TRN_AC_WRAP_less_15_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_RunInst_case_15_nv_scvector_cctor_data_0_ftd_1 <= 22'b0000000000000000000000;
    end
    else if ( ActUnit_RunInst_switch_lp_and_814_enex5 ) begin
      reg_ActUnit_RunInst_case_15_nv_scvector_cctor_data_0_ftd_1 <= nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_RunInst_case_15_nv_scvector_cctor_data_0_sva_30_26 <= 5'b00000;
    end
    else if ( ActUnit_RunInst_switch_lp_and_815_enex5 ) begin
      ActUnit_RunInst_case_15_nv_scvector_cctor_data_0_sva_30_26 <= nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_2_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1
          <= 22'b0000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_15_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_2_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1
          <= nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_6_for_2_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
          <= 5'b00000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_16_enex5 ) begin
      nv_scvector_cctor_nv_scvector_6_for_2_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
          <= nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_3_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1
          <= 22'b0000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_18_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_3_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1
          <= nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_6_for_3_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
          <= 5'b00000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_19_enex5 ) begin
      nv_scvector_cctor_nv_scvector_6_for_3_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
          <= nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_4_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1
          <= 22'b0000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_21_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_4_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1
          <= nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_6_for_4_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
          <= 5'b00000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_22_enex5 ) begin
      nv_scvector_cctor_nv_scvector_6_for_4_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
          <= nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_5_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1
          <= 22'b0000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_24_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_5_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1
          <= nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_6_for_5_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
          <= 5'b00000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_25_enex5 ) begin
      nv_scvector_cctor_nv_scvector_6_for_5_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
          <= nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_6_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1
          <= 22'b0000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_27_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_6_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1
          <= nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_6_for_6_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
          <= 5'b00000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_28_enex5 ) begin
      nv_scvector_cctor_nv_scvector_6_for_6_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
          <= nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_7_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1
          <= 22'b0000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_30_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_7_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1
          <= nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_6_for_7_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
          <= 5'b00000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_31_enex5 ) begin
      nv_scvector_cctor_nv_scvector_6_for_7_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
          <= nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_8_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1
          <= 22'b0000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_33_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_8_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1
          <= nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_6_for_8_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
          <= 5'b00000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_34_enex5 ) begin
      nv_scvector_cctor_nv_scvector_6_for_8_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
          <= nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_9_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1
          <= 22'b0000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_36_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_9_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1
          <= nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_6_for_9_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
          <= 5'b00000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_37_enex5 ) begin
      nv_scvector_cctor_nv_scvector_6_for_9_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
          <= nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_10_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1
          <= 22'b0000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_39_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_10_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1
          <= nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_6_for_10_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
          <= 5'b00000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_40_enex5 ) begin
      nv_scvector_cctor_nv_scvector_6_for_10_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
          <= nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_11_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1
          <= 22'b0000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_42_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_11_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1
          <= nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_6_for_11_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
          <= 5'b00000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_43_enex5 ) begin
      nv_scvector_cctor_nv_scvector_6_for_11_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
          <= nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_12_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1
          <= 22'b0000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_45_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_12_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1
          <= nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_6_for_12_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
          <= 5'b00000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_46_enex5 ) begin
      nv_scvector_cctor_nv_scvector_6_for_12_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
          <= nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_13_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1
          <= 22'b0000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_48_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_13_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1
          <= nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_6_for_13_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
          <= 5'b00000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_49_enex5 ) begin
      nv_scvector_cctor_nv_scvector_6_for_13_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
          <= nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_14_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1
          <= 22'b0000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_51_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_14_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1
          <= nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_6_for_14_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
          <= 5'b00000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_52_enex5 ) begin
      nv_scvector_cctor_nv_scvector_6_for_14_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
          <= nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_15_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1
          <= 22'b0000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_54_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_15_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1
          <= nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_6_for_15_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
          <= 5'b00000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_55_enex5 ) begin
      nv_scvector_cctor_nv_scvector_6_for_15_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
          <= nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_16_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1
          <= 22'b0000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_57_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_16_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1
          <= nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nv_scvector_cctor_nv_scvector_6_for_16_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
          <= 5'b00000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_58_enex5 ) begin
      nv_scvector_cctor_nv_scvector_6_for_16_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26
          <= nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_16_slc_32_1_svs <= 1'b0;
      Gelu_for_15_slc_32_1_svs <= 1'b0;
      Gelu_for_14_slc_32_1_svs <= 1'b0;
      Gelu_for_13_slc_32_1_svs <= 1'b0;
      Gelu_for_12_slc_32_1_svs <= 1'b0;
      Gelu_for_11_slc_32_1_svs <= 1'b0;
      Gelu_for_10_slc_32_1_svs <= 1'b0;
      Gelu_for_9_slc_32_1_svs <= 1'b0;
      Gelu_for_8_slc_32_1_svs <= 1'b0;
      Gelu_for_7_slc_32_1_svs <= 1'b0;
      Gelu_for_6_slc_32_1_svs <= 1'b0;
      Gelu_for_5_slc_32_1_svs <= 1'b0;
      Gelu_for_4_slc_32_1_svs <= 1'b0;
      Gelu_for_3_slc_32_1_svs <= 1'b0;
      Gelu_for_2_slc_32_1_svs <= 1'b0;
      Gelu_for_1_slc_32_1_svs <= 1'b0;
    end
    else if ( Gelu_for_if_and_cse ) begin
      Gelu_for_16_slc_32_1_svs <= Gelu_for_if_less_tmp;
      Gelu_for_15_slc_32_1_svs <= Gelu_for_if_less_1_tmp;
      Gelu_for_14_slc_32_1_svs <= Gelu_for_if_less_2_tmp;
      Gelu_for_13_slc_32_1_svs <= Gelu_for_if_less_3_tmp;
      Gelu_for_12_slc_32_1_svs <= Gelu_for_if_less_4_tmp;
      Gelu_for_11_slc_32_1_svs <= Gelu_for_if_less_5_tmp;
      Gelu_for_10_slc_32_1_svs <= Gelu_for_if_less_6_tmp;
      Gelu_for_9_slc_32_1_svs <= Gelu_for_if_less_7_tmp;
      Gelu_for_8_slc_32_1_svs <= Gelu_for_if_less_8_tmp;
      Gelu_for_7_slc_32_1_svs <= Gelu_for_if_less_9_tmp;
      Gelu_for_6_slc_32_1_svs <= Gelu_for_if_less_10_tmp;
      Gelu_for_5_slc_32_1_svs <= Gelu_for_if_less_11_tmp;
      Gelu_for_4_slc_32_1_svs <= Gelu_for_if_less_12_tmp;
      Gelu_for_3_slc_32_1_svs <= Gelu_for_if_less_13_tmp;
      Gelu_for_2_slc_32_1_svs <= Gelu_for_if_less_14_tmp;
      Gelu_for_1_slc_32_1_svs <= Gelu_for_if_less_15_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_asn_262_itm <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~ or_dcpl_822) & or_243_cse ) begin
      while_asn_262_itm <= is_start_sva;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_write_data_data_0_15_sva_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & while_and_1_tmp & (z_out[4]) ) begin
      act_write_data_data_0_15_sva_2_31 <= ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_31
          & ActUnit_RunInst_case_2_for_and_27_seb;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_write_data_data_0_15_sva_2_30_26 <= 5'b00000;
      reg_act_write_data_data_0_15_2_ftd <= 1'b0;
      reg_act_write_data_data_0_15_2_ftd_1 <= 3'b000;
      act_write_data_data_0_15_sva_2_21_0 <= 22'b0000000000000000000000;
      reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_nor_cse <= 1'b0;
      reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_2_cse <= 1'b0;
      reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_1_cse <= 1'b0;
      reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_cse <= 1'b0;
      ActUnit_RunInst_switch_lp_and_tmp <= 1'b0;
      while_nor_48_itm <= 1'b0;
      while_nor_32_itm <= 1'b0;
      while_nor_16_itm <= 1'b0;
      while_nor_itm <= 1'b0;
    end
    else if ( act_write_data_data_and_15_cse ) begin
      act_write_data_data_0_15_sva_2_30_26 <= MUX_v_5_2_2(ActUnit_RunInst_case_2_for_ActUnit_RunInst_case_2_for_and_1_nl,
          nv_scvector_cctor_nv_scvector_6_for_16_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26,
          and_dcpl_1240);
      reg_act_write_data_data_0_15_2_ftd <= MUX_s_1_2_2(ActUnit_RunInst_case_2_for_ActUnit_RunInst_case_2_for_and_2_nl,
          reg_nv_scvector_cctor_nv_scvector_6_for_16_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0,
          and_dcpl_1240);
      reg_act_write_data_data_0_15_2_ftd_1 <= MUX_v_3_2_2(ActUnit_RunInst_case_2_for_ActUnit_RunInst_case_2_for_and_4_nl,
          reg_nv_scvector_cctor_nv_scvector_6_for_16_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1,
          and_dcpl_1240);
      act_write_data_data_0_15_sva_2_21_0 <= MUX_v_22_2_2(ActUnit_RunInst_case_2_for_ActUnit_RunInst_case_2_for_and_3_nl,
          reg_nv_scvector_cctor_nv_scvector_6_for_16_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1,
          and_dcpl_1240);
      reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_nor_cse <= Tanh_for_nor_cse_sva_mx0w0;
      reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_2_cse <= Tanh_for_and_2_cse_sva_mx0w0;
      reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_1_cse <= Tanh_for_and_1_cse_sva_mx0w0;
      reg_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_cse <= Tanh_for_and_cse_sva_mx0w0;
      ActUnit_RunInst_switch_lp_and_tmp <= ActUnit_RunInst_switch_lp_and_tmp_mx0w0;
      while_nor_48_itm <= ~(ActUnit_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva
          | ActUnit_RunInst_switch_lp_and_32_tmp | ActUnit_RunInst_switch_lp_equal_tmp_3
          | ActUnit_RunInst_switch_lp_nor_tmp | ((~ Tanh_for_and_2_cse_sva_mx0w0)
          & ActUnit_RunInst_switch_lp_equal_tmp_4) | ((~ Tanh_for_and_2_cse_sva_mx0w0)
          & ActUnit_RunInst_switch_lp_equal_tmp_5) | ((~ Tanh_for_and_2_cse_sva_mx0w0)
          & ActUnit_RunInst_switch_lp_equal_tmp_6) | ((~ Tanh_for_and_2_cse_sva_mx0w0)
          & ActUnit_RunInst_switch_lp_equal_tmp_7) | ((~ Tanh_for_and_2_cse_sva_mx0w0)
          & ActUnit_RunInst_switch_lp_equal_tmp_8) | ((~ ActUnit_RunInst_switch_lp_and_48_tmp_1)
          & ActUnit_RunInst_switch_lp_equal_tmp_2));
      while_nor_32_itm <= ~(ActUnit_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva
          | ActUnit_RunInst_switch_lp_and_32_tmp | ActUnit_RunInst_switch_lp_equal_tmp_3
          | ActUnit_RunInst_switch_lp_nor_tmp | ((~ Tanh_for_and_cse_sva_mx0w0) &
          ActUnit_RunInst_switch_lp_equal_tmp_4) | ((~ Tanh_for_and_cse_sva_mx0w0)
          & ActUnit_RunInst_switch_lp_equal_tmp_5) | ((~ Tanh_for_and_cse_sva_mx0w0)
          & ActUnit_RunInst_switch_lp_equal_tmp_6) | ((~ Tanh_for_and_cse_sva_mx0w0)
          & ActUnit_RunInst_switch_lp_equal_tmp_7) | ((~ Tanh_for_and_cse_sva_mx0w0)
          & ActUnit_RunInst_switch_lp_equal_tmp_8) | ((~ ActUnit_RunInst_switch_lp_and_32_tmp_mx0w1)
          & ActUnit_RunInst_switch_lp_equal_tmp_2));
      while_nor_16_itm <= ~(ActUnit_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva
          | ActUnit_RunInst_switch_lp_and_32_tmp | ActUnit_RunInst_switch_lp_equal_tmp_3
          | ActUnit_RunInst_switch_lp_nor_tmp | ((~ Tanh_for_and_1_cse_sva_mx0w0)
          & ActUnit_RunInst_switch_lp_equal_tmp_4) | ((~ Tanh_for_and_1_cse_sva_mx0w0)
          & ActUnit_RunInst_switch_lp_equal_tmp_5) | ((~ Tanh_for_and_1_cse_sva_mx0w0)
          & ActUnit_RunInst_switch_lp_equal_tmp_6) | ((~ Tanh_for_and_1_cse_sva_mx0w0)
          & ActUnit_RunInst_switch_lp_equal_tmp_7) | ((~ Tanh_for_and_1_cse_sva_mx0w0)
          & ActUnit_RunInst_switch_lp_equal_tmp_8) | ((~ ActUnit_RunInst_switch_lp_and_16_tmp_mx0w1)
          & ActUnit_RunInst_switch_lp_equal_tmp_2));
      while_nor_itm <= ~(ActUnit_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva
          | ActUnit_RunInst_switch_lp_and_32_tmp | ActUnit_RunInst_switch_lp_equal_tmp_3
          | ActUnit_RunInst_switch_lp_nor_tmp | ((~ Tanh_for_nor_cse_sva_mx0w0) &
          ActUnit_RunInst_switch_lp_equal_tmp_4) | ((~ Tanh_for_nor_cse_sva_mx0w0)
          & ActUnit_RunInst_switch_lp_equal_tmp_5) | ((~ Tanh_for_nor_cse_sva_mx0w0)
          & ActUnit_RunInst_switch_lp_equal_tmp_6) | ((~ Tanh_for_nor_cse_sva_mx0w0)
          & ActUnit_RunInst_switch_lp_equal_tmp_7) | ((~ Tanh_for_nor_cse_sva_mx0w0)
          & ActUnit_RunInst_switch_lp_equal_tmp_8) | ((~ ActUnit_RunInst_switch_lp_and_tmp_mx0w0)
          & ActUnit_RunInst_switch_lp_equal_tmp_2));
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_write_data_data_0_0_sva_31 <= 1'b0;
    end
    else if ( act_write_data_data_and_ssc ) begin
      act_write_data_data_0_0_sva_31 <= ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_31;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_write_data_data_0_0_sva_30_26 <= 5'b00000;
      reg_act_write_data_data_0_0_2_ftd <= 1'b0;
      reg_act_write_data_data_0_0_2_ftd_1 <= 3'b000;
      act_write_data_data_0_0_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_write_data_data_and_16_ssc ) begin
      act_write_data_data_0_0_sva_30_26 <= MUX_v_5_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_30_26,
          ActUnit_RunInst_case_15_nv_scvector_cctor_data_0_sva_30_26, and_dcpl_1240);
      reg_act_write_data_data_0_0_2_ftd <= MUX_s_1_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_25,
          reg_ActUnit_RunInst_case_15_nv_scvector_cctor_data_0_ftd_rsp_0, and_dcpl_1240);
      reg_act_write_data_data_0_0_2_ftd_1 <= MUX_v_3_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_24_22,
          reg_ActUnit_RunInst_case_15_nv_scvector_cctor_data_0_ftd_rsp_1, and_dcpl_1240);
      act_write_data_data_0_0_sva_21_0 <= MUX_v_22_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_21_0,
          reg_ActUnit_RunInst_case_15_nv_scvector_cctor_data_0_ftd_1, and_dcpl_1240);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_write_data_data_0_14_sva_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~ or_dcpl_826) | and_dcpl_847 | and_dcpl_1240) )
        begin
      act_write_data_data_0_14_sva_31 <= act_write_data_data_act_write_data_data_and_26_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_write_data_data_0_14_sva_30_26 <= 5'b00000;
      act_write_data_data_0_14_sva_25 <= 1'b0;
      act_write_data_data_0_14_sva_24_22 <= 3'b000;
      act_write_data_data_0_14_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( and_1821_cse ) begin
      act_write_data_data_0_14_sva_30_26 <= MUX_v_5_2_2(5'b00000, act_write_data_data_act_write_data_data_act_write_data_data_mux_nl,
          not_3249_nl);
      act_write_data_data_0_14_sva_25 <= act_write_data_data_act_write_data_data_act_write_data_data_mux_1_nl
          & (~ and_dcpl_847);
      act_write_data_data_0_14_sva_24_22 <= MUX_v_3_2_2(3'b000, act_write_data_data_act_write_data_data_act_write_data_data_mux_42_nl,
          not_8967_nl);
      act_write_data_data_0_14_sva_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          act_write_data_data_act_write_data_data_act_write_data_data_mux_2_nl, not_2573_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_write_data_data_0_1_sva_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~ or_dcpl_828) | and_dcpl_847 | and_dcpl_1240) )
        begin
      act_write_data_data_0_1_sva_31 <= act_write_data_data_act_write_data_data_and_26_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_write_data_data_0_1_sva_30_26 <= 5'b00000;
      act_write_data_data_0_1_sva_25 <= 1'b0;
      act_write_data_data_0_1_sva_24_22 <= 3'b000;
      act_write_data_data_0_1_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( and_1824_cse ) begin
      act_write_data_data_0_1_sva_30_26 <= MUX_v_5_2_2(5'b00000, act_write_data_data_act_write_data_data_act_write_data_data_mux_3_nl,
          not_3247_nl);
      act_write_data_data_0_1_sva_25 <= act_write_data_data_act_write_data_data_act_write_data_data_mux_4_nl
          & (~ and_dcpl_847);
      act_write_data_data_0_1_sva_24_22 <= MUX_v_3_2_2(3'b000, act_write_data_data_act_write_data_data_act_write_data_data_mux_43_nl,
          not_8966_nl);
      act_write_data_data_0_1_sva_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          act_write_data_data_act_write_data_data_act_write_data_data_mux_5_nl, not_2571_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_write_data_data_0_13_sva_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~ or_dcpl_829) | and_dcpl_847 | and_dcpl_1240) )
        begin
      act_write_data_data_0_13_sva_31 <= act_write_data_data_act_write_data_data_and_26_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_write_data_data_0_13_sva_30_26 <= 5'b00000;
      act_write_data_data_0_13_sva_25 <= 1'b0;
      act_write_data_data_0_13_sva_24_22 <= 3'b000;
      act_write_data_data_0_13_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( and_1827_cse ) begin
      act_write_data_data_0_13_sva_30_26 <= MUX_v_5_2_2(5'b00000, act_write_data_data_act_write_data_data_act_write_data_data_mux_6_nl,
          not_3245_nl);
      act_write_data_data_0_13_sva_25 <= act_write_data_data_act_write_data_data_act_write_data_data_mux_7_nl
          & (~ and_dcpl_847);
      act_write_data_data_0_13_sva_24_22 <= MUX_v_3_2_2(3'b000, act_write_data_data_act_write_data_data_act_write_data_data_mux_44_nl,
          not_8965_nl);
      act_write_data_data_0_13_sva_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          act_write_data_data_act_write_data_data_act_write_data_data_mux_8_nl, not_2569_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_write_data_data_0_2_sva_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~ or_dcpl_830) | and_dcpl_847 | and_dcpl_1240) )
        begin
      act_write_data_data_0_2_sva_31 <= act_write_data_data_act_write_data_data_and_26_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_write_data_data_0_2_sva_30_26 <= 5'b00000;
      act_write_data_data_0_2_sva_25 <= 1'b0;
      act_write_data_data_0_2_sva_24_22 <= 3'b000;
      act_write_data_data_0_2_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( and_1830_cse ) begin
      act_write_data_data_0_2_sva_30_26 <= MUX_v_5_2_2(5'b00000, act_write_data_data_act_write_data_data_act_write_data_data_mux_9_nl,
          not_3243_nl);
      act_write_data_data_0_2_sva_25 <= act_write_data_data_act_write_data_data_act_write_data_data_mux_10_nl
          & (~ and_dcpl_847);
      act_write_data_data_0_2_sva_24_22 <= MUX_v_3_2_2(3'b000, act_write_data_data_act_write_data_data_act_write_data_data_mux_45_nl,
          not_8964_nl);
      act_write_data_data_0_2_sva_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          act_write_data_data_act_write_data_data_act_write_data_data_mux_11_nl,
          not_2567_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_write_data_data_0_12_sva_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~ or_dcpl_831) | and_dcpl_847 | and_dcpl_1240) )
        begin
      act_write_data_data_0_12_sva_31 <= act_write_data_data_act_write_data_data_and_26_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_write_data_data_0_12_sva_30_26 <= 5'b00000;
      act_write_data_data_0_12_sva_25 <= 1'b0;
      act_write_data_data_0_12_sva_24_22 <= 3'b000;
      act_write_data_data_0_12_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( and_1833_cse ) begin
      act_write_data_data_0_12_sva_30_26 <= MUX_v_5_2_2(5'b00000, act_write_data_data_act_write_data_data_act_write_data_data_mux_12_nl,
          not_3241_nl);
      act_write_data_data_0_12_sva_25 <= act_write_data_data_act_write_data_data_act_write_data_data_mux_13_nl
          & (~ and_dcpl_847);
      act_write_data_data_0_12_sva_24_22 <= MUX_v_3_2_2(3'b000, act_write_data_data_act_write_data_data_act_write_data_data_mux_46_nl,
          not_8963_nl);
      act_write_data_data_0_12_sva_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          act_write_data_data_act_write_data_data_act_write_data_data_mux_14_nl,
          not_2565_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_write_data_data_0_3_sva_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~ or_dcpl_833) | and_dcpl_847 | and_dcpl_1240) )
        begin
      act_write_data_data_0_3_sva_31 <= act_write_data_data_act_write_data_data_and_26_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_write_data_data_0_3_sva_30_26 <= 5'b00000;
      act_write_data_data_0_3_sva_25 <= 1'b0;
      act_write_data_data_0_3_sva_24_22 <= 3'b000;
      act_write_data_data_0_3_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( and_1836_cse ) begin
      act_write_data_data_0_3_sva_30_26 <= MUX_v_5_2_2(5'b00000, act_write_data_data_act_write_data_data_act_write_data_data_mux_15_nl,
          not_3239_nl);
      act_write_data_data_0_3_sva_25 <= act_write_data_data_act_write_data_data_act_write_data_data_mux_16_nl
          & (~ and_dcpl_847);
      act_write_data_data_0_3_sva_24_22 <= MUX_v_3_2_2(3'b000, act_write_data_data_act_write_data_data_act_write_data_data_mux_47_nl,
          not_8962_nl);
      act_write_data_data_0_3_sva_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          act_write_data_data_act_write_data_data_act_write_data_data_mux_17_nl,
          not_2563_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_write_data_data_0_11_sva_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~ or_dcpl_835) | and_dcpl_847 | and_dcpl_1240) )
        begin
      act_write_data_data_0_11_sva_31 <= act_write_data_data_act_write_data_data_and_26_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_write_data_data_0_11_sva_30_26 <= 5'b00000;
      act_write_data_data_0_11_sva_25 <= 1'b0;
      act_write_data_data_0_11_sva_24_22 <= 3'b000;
      act_write_data_data_0_11_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( and_1839_cse ) begin
      act_write_data_data_0_11_sva_30_26 <= MUX_v_5_2_2(5'b00000, act_write_data_data_act_write_data_data_act_write_data_data_mux_18_nl,
          not_3237_nl);
      act_write_data_data_0_11_sva_25 <= act_write_data_data_act_write_data_data_act_write_data_data_mux_19_nl
          & (~ and_dcpl_847);
      act_write_data_data_0_11_sva_24_22 <= MUX_v_3_2_2(3'b000, act_write_data_data_act_write_data_data_act_write_data_data_mux_48_nl,
          not_8961_nl);
      act_write_data_data_0_11_sva_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          act_write_data_data_act_write_data_data_act_write_data_data_mux_20_nl,
          not_2561_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_write_data_data_0_4_sva_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~ or_dcpl_837) | and_dcpl_847 | and_dcpl_1240) )
        begin
      act_write_data_data_0_4_sva_31 <= act_write_data_data_act_write_data_data_and_26_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_write_data_data_0_4_sva_30_26 <= 5'b00000;
      act_write_data_data_0_4_sva_25 <= 1'b0;
      act_write_data_data_0_4_sva_24_22 <= 3'b000;
      act_write_data_data_0_4_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( and_1842_cse ) begin
      act_write_data_data_0_4_sva_30_26 <= MUX_v_5_2_2(5'b00000, act_write_data_data_act_write_data_data_act_write_data_data_mux_21_nl,
          not_3235_nl);
      act_write_data_data_0_4_sva_25 <= act_write_data_data_act_write_data_data_act_write_data_data_mux_22_nl
          & (~ and_dcpl_847);
      act_write_data_data_0_4_sva_24_22 <= MUX_v_3_2_2(3'b000, act_write_data_data_act_write_data_data_act_write_data_data_mux_49_nl,
          not_8960_nl);
      act_write_data_data_0_4_sva_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          act_write_data_data_act_write_data_data_act_write_data_data_mux_23_nl,
          not_2559_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_write_data_data_0_10_sva_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~ or_dcpl_838) | and_dcpl_847 | and_dcpl_1240) )
        begin
      act_write_data_data_0_10_sva_31 <= act_write_data_data_act_write_data_data_and_26_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_write_data_data_0_10_sva_30_26 <= 5'b00000;
      act_write_data_data_0_10_sva_25 <= 1'b0;
      act_write_data_data_0_10_sva_24_22 <= 3'b000;
      act_write_data_data_0_10_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( and_1845_cse ) begin
      act_write_data_data_0_10_sva_30_26 <= MUX_v_5_2_2(5'b00000, act_write_data_data_act_write_data_data_act_write_data_data_mux_24_nl,
          not_3233_nl);
      act_write_data_data_0_10_sva_25 <= act_write_data_data_act_write_data_data_act_write_data_data_mux_25_nl
          & (~ and_dcpl_847);
      act_write_data_data_0_10_sva_24_22 <= MUX_v_3_2_2(3'b000, act_write_data_data_act_write_data_data_act_write_data_data_mux_50_nl,
          not_8959_nl);
      act_write_data_data_0_10_sva_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          act_write_data_data_act_write_data_data_act_write_data_data_mux_26_nl,
          not_2557_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_write_data_data_0_5_sva_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~ or_dcpl_839) | and_dcpl_847 | and_dcpl_1240) )
        begin
      act_write_data_data_0_5_sva_31 <= act_write_data_data_act_write_data_data_and_26_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_write_data_data_0_5_sva_30_26 <= 5'b00000;
      act_write_data_data_0_5_sva_25 <= 1'b0;
      act_write_data_data_0_5_sva_24_22 <= 3'b000;
      act_write_data_data_0_5_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( and_1848_cse ) begin
      act_write_data_data_0_5_sva_30_26 <= MUX_v_5_2_2(5'b00000, act_write_data_data_act_write_data_data_act_write_data_data_mux_27_nl,
          not_3231_nl);
      act_write_data_data_0_5_sva_25 <= act_write_data_data_act_write_data_data_act_write_data_data_mux_28_nl
          & (~ and_dcpl_847);
      act_write_data_data_0_5_sva_24_22 <= MUX_v_3_2_2(3'b000, act_write_data_data_act_write_data_data_act_write_data_data_mux_51_nl,
          not_8958_nl);
      act_write_data_data_0_5_sva_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          act_write_data_data_act_write_data_data_act_write_data_data_mux_29_nl,
          not_2555_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_write_data_data_0_9_sva_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~ or_dcpl_840) | and_dcpl_847 | and_dcpl_1240) )
        begin
      act_write_data_data_0_9_sva_31 <= act_write_data_data_act_write_data_data_and_26_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_write_data_data_0_9_sva_30_26 <= 5'b00000;
      act_write_data_data_0_9_sva_25 <= 1'b0;
      act_write_data_data_0_9_sva_24_22 <= 3'b000;
      act_write_data_data_0_9_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( and_1851_cse ) begin
      act_write_data_data_0_9_sva_30_26 <= MUX_v_5_2_2(5'b00000, act_write_data_data_act_write_data_data_act_write_data_data_mux_30_nl,
          not_3229_nl);
      act_write_data_data_0_9_sva_25 <= act_write_data_data_act_write_data_data_act_write_data_data_mux_31_nl
          & (~ and_dcpl_847);
      act_write_data_data_0_9_sva_24_22 <= MUX_v_3_2_2(3'b000, act_write_data_data_act_write_data_data_act_write_data_data_mux_52_nl,
          not_8957_nl);
      act_write_data_data_0_9_sva_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          act_write_data_data_act_write_data_data_act_write_data_data_mux_32_nl,
          not_2553_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_write_data_data_0_6_sva_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~ or_dcpl_841) | and_dcpl_847 | and_dcpl_1240) )
        begin
      act_write_data_data_0_6_sva_31 <= act_write_data_data_act_write_data_data_and_26_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_write_data_data_0_6_sva_30_26 <= 5'b00000;
      act_write_data_data_0_6_sva_25 <= 1'b0;
      act_write_data_data_0_6_sva_24_22 <= 3'b000;
      act_write_data_data_0_6_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( and_1854_cse ) begin
      act_write_data_data_0_6_sva_30_26 <= MUX_v_5_2_2(5'b00000, act_write_data_data_act_write_data_data_act_write_data_data_mux_33_nl,
          not_3227_nl);
      act_write_data_data_0_6_sva_25 <= act_write_data_data_act_write_data_data_act_write_data_data_mux_34_nl
          & (~ and_dcpl_847);
      act_write_data_data_0_6_sva_24_22 <= MUX_v_3_2_2(3'b000, act_write_data_data_act_write_data_data_act_write_data_data_mux_53_nl,
          not_8956_nl);
      act_write_data_data_0_6_sva_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          act_write_data_data_act_write_data_data_act_write_data_data_mux_35_nl,
          not_2551_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_write_data_data_0_8_sva_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~ or_dcpl_842) | and_dcpl_847 | and_dcpl_1240) )
        begin
      act_write_data_data_0_8_sva_31 <= act_write_data_data_act_write_data_data_and_26_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_write_data_data_0_8_sva_30_26 <= 5'b00000;
      act_write_data_data_0_8_sva_25 <= 1'b0;
      act_write_data_data_0_8_sva_24_22 <= 3'b000;
      act_write_data_data_0_8_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( and_1857_cse ) begin
      act_write_data_data_0_8_sva_30_26 <= MUX_v_5_2_2(5'b00000, act_write_data_data_act_write_data_data_act_write_data_data_mux_36_nl,
          not_3225_nl);
      act_write_data_data_0_8_sva_25 <= act_write_data_data_act_write_data_data_act_write_data_data_mux_37_nl
          & (~ and_dcpl_847);
      act_write_data_data_0_8_sva_24_22 <= MUX_v_3_2_2(3'b000, act_write_data_data_act_write_data_data_act_write_data_data_mux_54_nl,
          not_8955_nl);
      act_write_data_data_0_8_sva_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          act_write_data_data_act_write_data_data_act_write_data_data_mux_38_nl,
          not_2549_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_write_data_data_0_7_sva_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~ or_dcpl_843) | and_dcpl_847 | and_dcpl_1240) )
        begin
      act_write_data_data_0_7_sva_31 <= act_write_data_data_act_write_data_data_and_26_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_write_data_data_0_7_sva_30_26 <= 5'b00000;
      act_write_data_data_0_7_sva_25 <= 1'b0;
      act_write_data_data_0_7_sva_24_22 <= 3'b000;
      act_write_data_data_0_7_sva_21_0 <= 22'b0000000000000000000000;
    end
    else if ( and_1860_cse ) begin
      act_write_data_data_0_7_sva_30_26 <= MUX_v_5_2_2(5'b00000, act_write_data_data_act_write_data_data_act_write_data_data_mux_39_nl,
          not_3223_nl);
      act_write_data_data_0_7_sva_25 <= act_write_data_data_act_write_data_data_act_write_data_data_mux_40_nl
          & (~ and_dcpl_847);
      act_write_data_data_0_7_sva_24_22 <= MUX_v_3_2_2(3'b000, act_write_data_data_act_write_data_data_act_write_data_data_mux_55_nl,
          not_8954_nl);
      act_write_data_data_0_7_sva_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000,
          act_write_data_data_act_write_data_data_act_write_data_data_mux_41_nl,
          not_2547_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_RunInst_switch_lp_and_32_tmp <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~(((fsm_output[1]) ^ (fsm_output[2])) & (~((fsm_output[0])
        | (fsm_output[3]))))) ) begin
      ActUnit_RunInst_switch_lp_and_32_tmp <= MUX_s_1_2_2(ActUnit_RunInst_switch_lp_equal_tmp_1_mx0w0,
          ActUnit_RunInst_switch_lp_and_32_tmp_mx0w1, and_dcpl_331);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva
          <= 1'b0;
    end
    else if ( ActUnitRun_wen & (((z_out[4]) & (~(mux_445_nl & (~ (fsm_output[3])))))
        | and_dcpl_847 | and_dcpl_331 | and_dcpl_1244 | ActUnit_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva_mx0c4
        | and_dcpl_1104) ) begin
      ActUnit_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva
          <= MUX1HOT_s_1_5_2(ActUnit_RunInst_switch_lp_equal_tmp_9, ActUnit_RunInst_switch_lp_and_16_tmp_mx0w1,
          start_PopNB_mioi_return_rsc_z_mxwt, ActUnit_CheckStart_if_ActUnit_CheckStart_if_and_nl,
          act_config_InstIncr_act_config_InstIncr_if_and_svs_1, {and_dcpl_847 , and_dcpl_331
          , and_dcpl_1244 , ActUnit_RunInst_switch_lp_or_1_nl , and_dcpl_1104});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_for_i_4_0_sva_3_0 <= 4'b0000;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp ) begin
      ActUnit_PushOutput_if_for_i_4_0_sva_3_0 <= MUX_v_4_2_2(4'b0000, (z_out[3:0]),
          ActUnit_PushOutput_if_for_i_not_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_30_26 <= 5'b00000;
    end
    else if ( ActUnit_RunInst_switch_lp_and_811_cse ) begin
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_30_26 <= MUX1HOT_v_5_3_2(act_read_addrs_sva_2_mx0w0,
          Silu_for_Silu_for_and_16_nl, ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_30_26_2,
          {and_dcpl_847 , and_dcpl_1112 , and_dcpl_1235});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_read_req_valid_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((and_dcpl_1143 & (fsm_output[1]) & nor_1441_cse)
        | and_dcpl_1233) ) begin
      act_read_req_valid_lpi_1_dfm_6 <= MUX_s_1_2_2(ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_ActUnit_RunInst_switch_lp_nor_2_tmp,
          ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_5_nl, and_dcpl_1233);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_mem_banks_read_for_mux_15_itm <= 32'b00000000000000000000000000000000;
      act_mem_banks_read_for_mux_14_itm <= 32'b00000000000000000000000000000000;
      act_mem_banks_read_for_mux_13_itm <= 32'b00000000000000000000000000000000;
      act_mem_banks_read_for_mux_12_itm <= 32'b00000000000000000000000000000000;
      act_mem_banks_read_for_mux_11_itm <= 32'b00000000000000000000000000000000;
      act_mem_banks_read_for_mux_10_itm <= 32'b00000000000000000000000000000000;
      act_mem_banks_read_for_mux_9_itm <= 32'b00000000000000000000000000000000;
      act_mem_banks_read_for_mux_8_itm <= 32'b00000000000000000000000000000000;
      act_mem_banks_read_for_mux_7_itm <= 32'b00000000000000000000000000000000;
      act_mem_banks_read_for_mux_6_itm <= 32'b00000000000000000000000000000000;
      act_mem_banks_read_for_mux_5_itm <= 32'b00000000000000000000000000000000;
      act_mem_banks_read_for_mux_4_itm <= 32'b00000000000000000000000000000000;
      act_mem_banks_read_for_mux_3_itm <= 32'b00000000000000000000000000000000;
      act_mem_banks_read_for_mux_2_itm <= 32'b00000000000000000000000000000000;
      act_mem_banks_read_for_mux_1_itm <= 32'b00000000000000000000000000000000;
      act_mem_banks_read_for_mux_itm <= 32'b00000000000000000000000000000000;
    end
    else if ( act_mem_banks_read_for_and_cse ) begin
      act_mem_banks_read_for_mux_15_itm <= MUX_v_32_32_2(act_mem_banks_bank_a_0_31_0_sva_dfm,
          act_mem_banks_bank_a_1_31_0_sva_dfm, act_mem_banks_bank_a_2_31_0_sva_dfm,
          act_mem_banks_bank_a_3_31_0_sva_dfm, act_mem_banks_bank_a_4_31_0_sva_dfm,
          act_mem_banks_bank_a_5_31_0_sva_dfm, act_mem_banks_bank_a_6_31_0_sva_dfm,
          act_mem_banks_bank_a_7_31_0_sva_dfm, act_mem_banks_bank_a_8_31_0_sva_dfm,
          act_mem_banks_bank_a_9_31_0_sva_dfm, act_mem_banks_bank_a_10_31_0_sva_dfm,
          act_mem_banks_bank_a_11_31_0_sva_dfm, act_mem_banks_bank_a_12_31_0_sva_dfm,
          act_mem_banks_bank_a_13_31_0_sva_dfm, act_mem_banks_bank_a_14_31_0_sva_dfm,
          act_mem_banks_bank_a_15_31_0_sva_dfm, act_mem_banks_bank_a_16_31_0_sva_dfm,
          act_mem_banks_bank_a_17_31_0_sva_dfm, act_mem_banks_bank_a_18_31_0_sva_dfm,
          act_mem_banks_bank_a_19_31_0_sva_dfm, act_mem_banks_bank_a_20_31_0_sva_dfm,
          act_mem_banks_bank_a_21_31_0_sva_dfm, act_mem_banks_bank_a_22_31_0_sva_dfm,
          act_mem_banks_bank_a_23_31_0_sva_dfm, act_mem_banks_bank_a_24_31_0_sva_dfm,
          act_mem_banks_bank_a_25_31_0_sva_dfm, act_mem_banks_bank_a_26_31_0_sva_dfm,
          act_mem_banks_bank_a_27_31_0_sva_dfm, act_mem_banks_bank_a_28_31_0_sva_dfm,
          act_mem_banks_bank_a_29_31_0_sva_dfm, act_mem_banks_bank_a_30_31_0_sva_dfm,
          act_mem_banks_bank_a_31_31_0_sva_dfm, while_mux_53_ssc_mx0);
      act_mem_banks_read_for_mux_14_itm <= MUX_v_32_32_2(act_mem_banks_bank_a_0_63_32_sva_dfm,
          act_mem_banks_bank_a_1_63_32_sva_dfm, act_mem_banks_bank_a_2_63_32_sva_dfm,
          act_mem_banks_bank_a_3_63_32_sva_dfm, act_mem_banks_bank_a_4_63_32_sva_dfm,
          act_mem_banks_bank_a_5_63_32_sva_dfm, act_mem_banks_bank_a_6_63_32_sva_dfm,
          act_mem_banks_bank_a_7_63_32_sva_dfm, act_mem_banks_bank_a_8_63_32_sva_dfm,
          act_mem_banks_bank_a_9_63_32_sva_dfm, act_mem_banks_bank_a_10_63_32_sva_dfm,
          act_mem_banks_bank_a_11_63_32_sva_dfm, act_mem_banks_bank_a_12_63_32_sva_dfm,
          act_mem_banks_bank_a_13_63_32_sva_dfm, act_mem_banks_bank_a_14_63_32_sva_dfm,
          act_mem_banks_bank_a_15_63_32_sva_dfm, act_mem_banks_bank_a_16_63_32_sva_dfm,
          act_mem_banks_bank_a_17_63_32_sva_dfm, act_mem_banks_bank_a_18_63_32_sva_dfm,
          act_mem_banks_bank_a_19_63_32_sva_dfm, act_mem_banks_bank_a_20_63_32_sva_dfm,
          act_mem_banks_bank_a_21_63_32_sva_dfm, act_mem_banks_bank_a_22_63_32_sva_dfm,
          act_mem_banks_bank_a_23_63_32_sva_dfm, act_mem_banks_bank_a_24_63_32_sva_dfm,
          act_mem_banks_bank_a_25_63_32_sva_dfm, act_mem_banks_bank_a_26_63_32_sva_dfm,
          act_mem_banks_bank_a_27_63_32_sva_dfm, act_mem_banks_bank_a_28_63_32_sva_dfm,
          act_mem_banks_bank_a_29_63_32_sva_dfm, act_mem_banks_bank_a_30_63_32_sva_dfm,
          act_mem_banks_bank_a_31_63_32_sva_dfm, while_mux_53_ssc_mx0);
      act_mem_banks_read_for_mux_13_itm <= MUX_v_32_32_2(act_mem_banks_bank_a_0_95_64_sva_dfm,
          act_mem_banks_bank_a_1_95_64_sva_dfm, act_mem_banks_bank_a_2_95_64_sva_dfm,
          act_mem_banks_bank_a_3_95_64_sva_dfm, act_mem_banks_bank_a_4_95_64_sva_dfm,
          act_mem_banks_bank_a_5_95_64_sva_dfm, act_mem_banks_bank_a_6_95_64_sva_dfm,
          act_mem_banks_bank_a_7_95_64_sva_dfm, act_mem_banks_bank_a_8_95_64_sva_dfm,
          act_mem_banks_bank_a_9_95_64_sva_dfm, act_mem_banks_bank_a_10_95_64_sva_dfm,
          act_mem_banks_bank_a_11_95_64_sva_dfm, act_mem_banks_bank_a_12_95_64_sva_dfm,
          act_mem_banks_bank_a_13_95_64_sva_dfm, act_mem_banks_bank_a_14_95_64_sva_dfm,
          act_mem_banks_bank_a_15_95_64_sva_dfm, act_mem_banks_bank_a_16_95_64_sva_dfm,
          act_mem_banks_bank_a_17_95_64_sva_dfm, act_mem_banks_bank_a_18_95_64_sva_dfm,
          act_mem_banks_bank_a_19_95_64_sva_dfm, act_mem_banks_bank_a_20_95_64_sva_dfm,
          act_mem_banks_bank_a_21_95_64_sva_dfm, act_mem_banks_bank_a_22_95_64_sva_dfm,
          act_mem_banks_bank_a_23_95_64_sva_dfm, act_mem_banks_bank_a_24_95_64_sva_dfm,
          act_mem_banks_bank_a_25_95_64_sva_dfm, act_mem_banks_bank_a_26_95_64_sva_dfm,
          act_mem_banks_bank_a_27_95_64_sva_dfm, act_mem_banks_bank_a_28_95_64_sva_dfm,
          act_mem_banks_bank_a_29_95_64_sva_dfm, act_mem_banks_bank_a_30_95_64_sva_dfm,
          act_mem_banks_bank_a_31_95_64_sva_dfm, while_mux_53_ssc_mx0);
      act_mem_banks_read_for_mux_12_itm <= MUX_v_32_32_2(act_mem_banks_bank_a_0_127_96_sva_dfm,
          act_mem_banks_bank_a_1_127_96_sva_dfm, act_mem_banks_bank_a_2_127_96_sva_dfm,
          act_mem_banks_bank_a_3_127_96_sva_dfm, act_mem_banks_bank_a_4_127_96_sva_dfm,
          act_mem_banks_bank_a_5_127_96_sva_dfm, act_mem_banks_bank_a_6_127_96_sva_dfm,
          act_mem_banks_bank_a_7_127_96_sva_dfm, act_mem_banks_bank_a_8_127_96_sva_dfm,
          act_mem_banks_bank_a_9_127_96_sva_dfm, act_mem_banks_bank_a_10_127_96_sva_dfm,
          act_mem_banks_bank_a_11_127_96_sva_dfm, act_mem_banks_bank_a_12_127_96_sva_dfm,
          act_mem_banks_bank_a_13_127_96_sva_dfm, act_mem_banks_bank_a_14_127_96_sva_dfm,
          act_mem_banks_bank_a_15_127_96_sva_dfm, act_mem_banks_bank_a_16_127_96_sva_dfm,
          act_mem_banks_bank_a_17_127_96_sva_dfm, act_mem_banks_bank_a_18_127_96_sva_dfm,
          act_mem_banks_bank_a_19_127_96_sva_dfm, act_mem_banks_bank_a_20_127_96_sva_dfm,
          act_mem_banks_bank_a_21_127_96_sva_dfm, act_mem_banks_bank_a_22_127_96_sva_dfm,
          act_mem_banks_bank_a_23_127_96_sva_dfm, act_mem_banks_bank_a_24_127_96_sva_dfm,
          act_mem_banks_bank_a_25_127_96_sva_dfm, act_mem_banks_bank_a_26_127_96_sva_dfm,
          act_mem_banks_bank_a_27_127_96_sva_dfm, act_mem_banks_bank_a_28_127_96_sva_dfm,
          act_mem_banks_bank_a_29_127_96_sva_dfm, act_mem_banks_bank_a_30_127_96_sva_dfm,
          act_mem_banks_bank_a_31_127_96_sva_dfm, while_mux_53_ssc_mx0);
      act_mem_banks_read_for_mux_11_itm <= MUX_v_32_32_2(act_mem_banks_bank_a_0_159_128_sva_dfm,
          act_mem_banks_bank_a_1_159_128_sva_dfm, act_mem_banks_bank_a_2_159_128_sva_dfm,
          act_mem_banks_bank_a_3_159_128_sva_dfm, act_mem_banks_bank_a_4_159_128_sva_dfm,
          act_mem_banks_bank_a_5_159_128_sva_dfm, act_mem_banks_bank_a_6_159_128_sva_dfm,
          act_mem_banks_bank_a_7_159_128_sva_dfm, act_mem_banks_bank_a_8_159_128_sva_dfm,
          act_mem_banks_bank_a_9_159_128_sva_dfm, act_mem_banks_bank_a_10_159_128_sva_dfm,
          act_mem_banks_bank_a_11_159_128_sva_dfm, act_mem_banks_bank_a_12_159_128_sva_dfm,
          act_mem_banks_bank_a_13_159_128_sva_dfm, act_mem_banks_bank_a_14_159_128_sva_dfm,
          act_mem_banks_bank_a_15_159_128_sva_dfm, act_mem_banks_bank_a_16_159_128_sva_dfm,
          act_mem_banks_bank_a_17_159_128_sva_dfm, act_mem_banks_bank_a_18_159_128_sva_dfm,
          act_mem_banks_bank_a_19_159_128_sva_dfm, act_mem_banks_bank_a_20_159_128_sva_dfm,
          act_mem_banks_bank_a_21_159_128_sva_dfm, act_mem_banks_bank_a_22_159_128_sva_dfm,
          act_mem_banks_bank_a_23_159_128_sva_dfm, act_mem_banks_bank_a_24_159_128_sva_dfm,
          act_mem_banks_bank_a_25_159_128_sva_dfm, act_mem_banks_bank_a_26_159_128_sva_dfm,
          act_mem_banks_bank_a_27_159_128_sva_dfm, act_mem_banks_bank_a_28_159_128_sva_dfm,
          act_mem_banks_bank_a_29_159_128_sva_dfm, act_mem_banks_bank_a_30_159_128_sva_dfm,
          act_mem_banks_bank_a_31_159_128_sva_dfm, while_mux_53_ssc_mx0);
      act_mem_banks_read_for_mux_10_itm <= MUX_v_32_32_2(act_mem_banks_bank_a_0_191_160_sva_dfm,
          act_mem_banks_bank_a_1_191_160_sva_dfm, act_mem_banks_bank_a_2_191_160_sva_dfm,
          act_mem_banks_bank_a_3_191_160_sva_dfm, act_mem_banks_bank_a_4_191_160_sva_dfm,
          act_mem_banks_bank_a_5_191_160_sva_dfm, act_mem_banks_bank_a_6_191_160_sva_dfm,
          act_mem_banks_bank_a_7_191_160_sva_dfm, act_mem_banks_bank_a_8_191_160_sva_dfm,
          act_mem_banks_bank_a_9_191_160_sva_dfm, act_mem_banks_bank_a_10_191_160_sva_dfm,
          act_mem_banks_bank_a_11_191_160_sva_dfm, act_mem_banks_bank_a_12_191_160_sva_dfm,
          act_mem_banks_bank_a_13_191_160_sva_dfm, act_mem_banks_bank_a_14_191_160_sva_dfm,
          act_mem_banks_bank_a_15_191_160_sva_dfm, act_mem_banks_bank_a_16_191_160_sva_dfm,
          act_mem_banks_bank_a_17_191_160_sva_dfm, act_mem_banks_bank_a_18_191_160_sva_dfm,
          act_mem_banks_bank_a_19_191_160_sva_dfm, act_mem_banks_bank_a_20_191_160_sva_dfm,
          act_mem_banks_bank_a_21_191_160_sva_dfm, act_mem_banks_bank_a_22_191_160_sva_dfm,
          act_mem_banks_bank_a_23_191_160_sva_dfm, act_mem_banks_bank_a_24_191_160_sva_dfm,
          act_mem_banks_bank_a_25_191_160_sva_dfm, act_mem_banks_bank_a_26_191_160_sva_dfm,
          act_mem_banks_bank_a_27_191_160_sva_dfm, act_mem_banks_bank_a_28_191_160_sva_dfm,
          act_mem_banks_bank_a_29_191_160_sva_dfm, act_mem_banks_bank_a_30_191_160_sva_dfm,
          act_mem_banks_bank_a_31_191_160_sva_dfm, while_mux_53_ssc_mx0);
      act_mem_banks_read_for_mux_9_itm <= MUX_v_32_32_2(act_mem_banks_bank_a_0_223_192_sva_dfm,
          act_mem_banks_bank_a_1_223_192_sva_dfm, act_mem_banks_bank_a_2_223_192_sva_dfm,
          act_mem_banks_bank_a_3_223_192_sva_dfm, act_mem_banks_bank_a_4_223_192_sva_dfm,
          act_mem_banks_bank_a_5_223_192_sva_dfm, act_mem_banks_bank_a_6_223_192_sva_dfm,
          act_mem_banks_bank_a_7_223_192_sva_dfm, act_mem_banks_bank_a_8_223_192_sva_dfm,
          act_mem_banks_bank_a_9_223_192_sva_dfm, act_mem_banks_bank_a_10_223_192_sva_dfm,
          act_mem_banks_bank_a_11_223_192_sva_dfm, act_mem_banks_bank_a_12_223_192_sva_dfm,
          act_mem_banks_bank_a_13_223_192_sva_dfm, act_mem_banks_bank_a_14_223_192_sva_dfm,
          act_mem_banks_bank_a_15_223_192_sva_dfm, act_mem_banks_bank_a_16_223_192_sva_dfm,
          act_mem_banks_bank_a_17_223_192_sva_dfm, act_mem_banks_bank_a_18_223_192_sva_dfm,
          act_mem_banks_bank_a_19_223_192_sva_dfm, act_mem_banks_bank_a_20_223_192_sva_dfm,
          act_mem_banks_bank_a_21_223_192_sva_dfm, act_mem_banks_bank_a_22_223_192_sva_dfm,
          act_mem_banks_bank_a_23_223_192_sva_dfm, act_mem_banks_bank_a_24_223_192_sva_dfm,
          act_mem_banks_bank_a_25_223_192_sva_dfm, act_mem_banks_bank_a_26_223_192_sva_dfm,
          act_mem_banks_bank_a_27_223_192_sva_dfm, act_mem_banks_bank_a_28_223_192_sva_dfm,
          act_mem_banks_bank_a_29_223_192_sva_dfm, act_mem_banks_bank_a_30_223_192_sva_dfm,
          act_mem_banks_bank_a_31_223_192_sva_dfm, while_mux_53_ssc_mx0);
      act_mem_banks_read_for_mux_8_itm <= MUX_v_32_32_2(act_mem_banks_bank_a_0_255_224_sva_dfm,
          act_mem_banks_bank_a_1_255_224_sva_dfm, act_mem_banks_bank_a_2_255_224_sva_dfm,
          act_mem_banks_bank_a_3_255_224_sva_dfm, act_mem_banks_bank_a_4_255_224_sva_dfm,
          act_mem_banks_bank_a_5_255_224_sva_dfm, act_mem_banks_bank_a_6_255_224_sva_dfm,
          act_mem_banks_bank_a_7_255_224_sva_dfm, act_mem_banks_bank_a_8_255_224_sva_dfm,
          act_mem_banks_bank_a_9_255_224_sva_dfm, act_mem_banks_bank_a_10_255_224_sva_dfm,
          act_mem_banks_bank_a_11_255_224_sva_dfm, act_mem_banks_bank_a_12_255_224_sva_dfm,
          act_mem_banks_bank_a_13_255_224_sva_dfm, act_mem_banks_bank_a_14_255_224_sva_dfm,
          act_mem_banks_bank_a_15_255_224_sva_dfm, act_mem_banks_bank_a_16_255_224_sva_dfm,
          act_mem_banks_bank_a_17_255_224_sva_dfm, act_mem_banks_bank_a_18_255_224_sva_dfm,
          act_mem_banks_bank_a_19_255_224_sva_dfm, act_mem_banks_bank_a_20_255_224_sva_dfm,
          act_mem_banks_bank_a_21_255_224_sva_dfm, act_mem_banks_bank_a_22_255_224_sva_dfm,
          act_mem_banks_bank_a_23_255_224_sva_dfm, act_mem_banks_bank_a_24_255_224_sva_dfm,
          act_mem_banks_bank_a_25_255_224_sva_dfm, act_mem_banks_bank_a_26_255_224_sva_dfm,
          act_mem_banks_bank_a_27_255_224_sva_dfm, act_mem_banks_bank_a_28_255_224_sva_dfm,
          act_mem_banks_bank_a_29_255_224_sva_dfm, act_mem_banks_bank_a_30_255_224_sva_dfm,
          act_mem_banks_bank_a_31_255_224_sva_dfm, while_mux_53_ssc_mx0);
      act_mem_banks_read_for_mux_7_itm <= MUX_v_32_32_2(act_mem_banks_bank_a_0_287_256_sva_dfm,
          act_mem_banks_bank_a_1_287_256_sva_dfm, act_mem_banks_bank_a_2_287_256_sva_dfm,
          act_mem_banks_bank_a_3_287_256_sva_dfm, act_mem_banks_bank_a_4_287_256_sva_dfm,
          act_mem_banks_bank_a_5_287_256_sva_dfm, act_mem_banks_bank_a_6_287_256_sva_dfm,
          act_mem_banks_bank_a_7_287_256_sva_dfm, act_mem_banks_bank_a_8_287_256_sva_dfm,
          act_mem_banks_bank_a_9_287_256_sva_dfm, act_mem_banks_bank_a_10_287_256_sva_dfm,
          act_mem_banks_bank_a_11_287_256_sva_dfm, act_mem_banks_bank_a_12_287_256_sva_dfm,
          act_mem_banks_bank_a_13_287_256_sva_dfm, act_mem_banks_bank_a_14_287_256_sva_dfm,
          act_mem_banks_bank_a_15_287_256_sva_dfm, act_mem_banks_bank_a_16_287_256_sva_dfm,
          act_mem_banks_bank_a_17_287_256_sva_dfm, act_mem_banks_bank_a_18_287_256_sva_dfm,
          act_mem_banks_bank_a_19_287_256_sva_dfm, act_mem_banks_bank_a_20_287_256_sva_dfm,
          act_mem_banks_bank_a_21_287_256_sva_dfm, act_mem_banks_bank_a_22_287_256_sva_dfm,
          act_mem_banks_bank_a_23_287_256_sva_dfm, act_mem_banks_bank_a_24_287_256_sva_dfm,
          act_mem_banks_bank_a_25_287_256_sva_dfm, act_mem_banks_bank_a_26_287_256_sva_dfm,
          act_mem_banks_bank_a_27_287_256_sva_dfm, act_mem_banks_bank_a_28_287_256_sva_dfm,
          act_mem_banks_bank_a_29_287_256_sva_dfm, act_mem_banks_bank_a_30_287_256_sva_dfm,
          act_mem_banks_bank_a_31_287_256_sva_dfm, while_mux_53_ssc_mx0);
      act_mem_banks_read_for_mux_6_itm <= MUX_v_32_32_2(act_mem_banks_bank_a_0_319_288_sva_dfm,
          act_mem_banks_bank_a_1_319_288_sva_dfm, act_mem_banks_bank_a_2_319_288_sva_dfm,
          act_mem_banks_bank_a_3_319_288_sva_dfm, act_mem_banks_bank_a_4_319_288_sva_dfm,
          act_mem_banks_bank_a_5_319_288_sva_dfm, act_mem_banks_bank_a_6_319_288_sva_dfm,
          act_mem_banks_bank_a_7_319_288_sva_dfm, act_mem_banks_bank_a_8_319_288_sva_dfm,
          act_mem_banks_bank_a_9_319_288_sva_dfm, act_mem_banks_bank_a_10_319_288_sva_dfm,
          act_mem_banks_bank_a_11_319_288_sva_dfm, act_mem_banks_bank_a_12_319_288_sva_dfm,
          act_mem_banks_bank_a_13_319_288_sva_dfm, act_mem_banks_bank_a_14_319_288_sva_dfm,
          act_mem_banks_bank_a_15_319_288_sva_dfm, act_mem_banks_bank_a_16_319_288_sva_dfm,
          act_mem_banks_bank_a_17_319_288_sva_dfm, act_mem_banks_bank_a_18_319_288_sva_dfm,
          act_mem_banks_bank_a_19_319_288_sva_dfm, act_mem_banks_bank_a_20_319_288_sva_dfm,
          act_mem_banks_bank_a_21_319_288_sva_dfm, act_mem_banks_bank_a_22_319_288_sva_dfm,
          act_mem_banks_bank_a_23_319_288_sva_dfm, act_mem_banks_bank_a_24_319_288_sva_dfm,
          act_mem_banks_bank_a_25_319_288_sva_dfm, act_mem_banks_bank_a_26_319_288_sva_dfm,
          act_mem_banks_bank_a_27_319_288_sva_dfm, act_mem_banks_bank_a_28_319_288_sva_dfm,
          act_mem_banks_bank_a_29_319_288_sva_dfm, act_mem_banks_bank_a_30_319_288_sva_dfm,
          act_mem_banks_bank_a_31_319_288_sva_dfm, while_mux_53_ssc_mx0);
      act_mem_banks_read_for_mux_5_itm <= MUX_v_32_32_2(act_mem_banks_bank_a_0_351_320_sva_dfm,
          act_mem_banks_bank_a_1_351_320_sva_dfm, act_mem_banks_bank_a_2_351_320_sva_dfm,
          act_mem_banks_bank_a_3_351_320_sva_dfm, act_mem_banks_bank_a_4_351_320_sva_dfm,
          act_mem_banks_bank_a_5_351_320_sva_dfm, act_mem_banks_bank_a_6_351_320_sva_dfm,
          act_mem_banks_bank_a_7_351_320_sva_dfm, act_mem_banks_bank_a_8_351_320_sva_dfm,
          act_mem_banks_bank_a_9_351_320_sva_dfm, act_mem_banks_bank_a_10_351_320_sva_dfm,
          act_mem_banks_bank_a_11_351_320_sva_dfm, act_mem_banks_bank_a_12_351_320_sva_dfm,
          act_mem_banks_bank_a_13_351_320_sva_dfm, act_mem_banks_bank_a_14_351_320_sva_dfm,
          act_mem_banks_bank_a_15_351_320_sva_dfm, act_mem_banks_bank_a_16_351_320_sva_dfm,
          act_mem_banks_bank_a_17_351_320_sva_dfm, act_mem_banks_bank_a_18_351_320_sva_dfm,
          act_mem_banks_bank_a_19_351_320_sva_dfm, act_mem_banks_bank_a_20_351_320_sva_dfm,
          act_mem_banks_bank_a_21_351_320_sva_dfm, act_mem_banks_bank_a_22_351_320_sva_dfm,
          act_mem_banks_bank_a_23_351_320_sva_dfm, act_mem_banks_bank_a_24_351_320_sva_dfm,
          act_mem_banks_bank_a_25_351_320_sva_dfm, act_mem_banks_bank_a_26_351_320_sva_dfm,
          act_mem_banks_bank_a_27_351_320_sva_dfm, act_mem_banks_bank_a_28_351_320_sva_dfm,
          act_mem_banks_bank_a_29_351_320_sva_dfm, act_mem_banks_bank_a_30_351_320_sva_dfm,
          act_mem_banks_bank_a_31_351_320_sva_dfm, while_mux_53_ssc_mx0);
      act_mem_banks_read_for_mux_4_itm <= MUX_v_32_32_2(act_mem_banks_bank_a_0_383_352_sva_dfm,
          act_mem_banks_bank_a_1_383_352_sva_dfm, act_mem_banks_bank_a_2_383_352_sva_dfm,
          act_mem_banks_bank_a_3_383_352_sva_dfm, act_mem_banks_bank_a_4_383_352_sva_dfm,
          act_mem_banks_bank_a_5_383_352_sva_dfm, act_mem_banks_bank_a_6_383_352_sva_dfm,
          act_mem_banks_bank_a_7_383_352_sva_dfm, act_mem_banks_bank_a_8_383_352_sva_dfm,
          act_mem_banks_bank_a_9_383_352_sva_dfm, act_mem_banks_bank_a_10_383_352_sva_dfm,
          act_mem_banks_bank_a_11_383_352_sva_dfm, act_mem_banks_bank_a_12_383_352_sva_dfm,
          act_mem_banks_bank_a_13_383_352_sva_dfm, act_mem_banks_bank_a_14_383_352_sva_dfm,
          act_mem_banks_bank_a_15_383_352_sva_dfm, act_mem_banks_bank_a_16_383_352_sva_dfm,
          act_mem_banks_bank_a_17_383_352_sva_dfm, act_mem_banks_bank_a_18_383_352_sva_dfm,
          act_mem_banks_bank_a_19_383_352_sva_dfm, act_mem_banks_bank_a_20_383_352_sva_dfm,
          act_mem_banks_bank_a_21_383_352_sva_dfm, act_mem_banks_bank_a_22_383_352_sva_dfm,
          act_mem_banks_bank_a_23_383_352_sva_dfm, act_mem_banks_bank_a_24_383_352_sva_dfm,
          act_mem_banks_bank_a_25_383_352_sva_dfm, act_mem_banks_bank_a_26_383_352_sva_dfm,
          act_mem_banks_bank_a_27_383_352_sva_dfm, act_mem_banks_bank_a_28_383_352_sva_dfm,
          act_mem_banks_bank_a_29_383_352_sva_dfm, act_mem_banks_bank_a_30_383_352_sva_dfm,
          act_mem_banks_bank_a_31_383_352_sva_dfm, while_mux_53_ssc_mx0);
      act_mem_banks_read_for_mux_3_itm <= MUX_v_32_32_2(act_mem_banks_bank_a_0_415_384_sva_dfm,
          act_mem_banks_bank_a_1_415_384_sva_dfm, act_mem_banks_bank_a_2_415_384_sva_dfm,
          act_mem_banks_bank_a_3_415_384_sva_dfm, act_mem_banks_bank_a_4_415_384_sva_dfm,
          act_mem_banks_bank_a_5_415_384_sva_dfm, act_mem_banks_bank_a_6_415_384_sva_dfm,
          act_mem_banks_bank_a_7_415_384_sva_dfm, act_mem_banks_bank_a_8_415_384_sva_dfm,
          act_mem_banks_bank_a_9_415_384_sva_dfm, act_mem_banks_bank_a_10_415_384_sva_dfm,
          act_mem_banks_bank_a_11_415_384_sva_dfm, act_mem_banks_bank_a_12_415_384_sva_dfm,
          act_mem_banks_bank_a_13_415_384_sva_dfm, act_mem_banks_bank_a_14_415_384_sva_dfm,
          act_mem_banks_bank_a_15_415_384_sva_dfm, act_mem_banks_bank_a_16_415_384_sva_dfm,
          act_mem_banks_bank_a_17_415_384_sva_dfm, act_mem_banks_bank_a_18_415_384_sva_dfm,
          act_mem_banks_bank_a_19_415_384_sva_dfm, act_mem_banks_bank_a_20_415_384_sva_dfm,
          act_mem_banks_bank_a_21_415_384_sva_dfm, act_mem_banks_bank_a_22_415_384_sva_dfm,
          act_mem_banks_bank_a_23_415_384_sva_dfm, act_mem_banks_bank_a_24_415_384_sva_dfm,
          act_mem_banks_bank_a_25_415_384_sva_dfm, act_mem_banks_bank_a_26_415_384_sva_dfm,
          act_mem_banks_bank_a_27_415_384_sva_dfm, act_mem_banks_bank_a_28_415_384_sva_dfm,
          act_mem_banks_bank_a_29_415_384_sva_dfm, act_mem_banks_bank_a_30_415_384_sva_dfm,
          act_mem_banks_bank_a_31_415_384_sva_dfm, while_mux_53_ssc_mx0);
      act_mem_banks_read_for_mux_2_itm <= MUX_v_32_32_2(act_mem_banks_bank_a_0_447_416_sva_dfm,
          act_mem_banks_bank_a_1_447_416_sva_dfm, act_mem_banks_bank_a_2_447_416_sva_dfm,
          act_mem_banks_bank_a_3_447_416_sva_dfm, act_mem_banks_bank_a_4_447_416_sva_dfm,
          act_mem_banks_bank_a_5_447_416_sva_dfm, act_mem_banks_bank_a_6_447_416_sva_dfm,
          act_mem_banks_bank_a_7_447_416_sva_dfm, act_mem_banks_bank_a_8_447_416_sva_dfm,
          act_mem_banks_bank_a_9_447_416_sva_dfm, act_mem_banks_bank_a_10_447_416_sva_dfm,
          act_mem_banks_bank_a_11_447_416_sva_dfm, act_mem_banks_bank_a_12_447_416_sva_dfm,
          act_mem_banks_bank_a_13_447_416_sva_dfm, act_mem_banks_bank_a_14_447_416_sva_dfm,
          act_mem_banks_bank_a_15_447_416_sva_dfm, act_mem_banks_bank_a_16_447_416_sva_dfm,
          act_mem_banks_bank_a_17_447_416_sva_dfm, act_mem_banks_bank_a_18_447_416_sva_dfm,
          act_mem_banks_bank_a_19_447_416_sva_dfm, act_mem_banks_bank_a_20_447_416_sva_dfm,
          act_mem_banks_bank_a_21_447_416_sva_dfm, act_mem_banks_bank_a_22_447_416_sva_dfm,
          act_mem_banks_bank_a_23_447_416_sva_dfm, act_mem_banks_bank_a_24_447_416_sva_dfm,
          act_mem_banks_bank_a_25_447_416_sva_dfm, act_mem_banks_bank_a_26_447_416_sva_dfm,
          act_mem_banks_bank_a_27_447_416_sva_dfm, act_mem_banks_bank_a_28_447_416_sva_dfm,
          act_mem_banks_bank_a_29_447_416_sva_dfm, act_mem_banks_bank_a_30_447_416_sva_dfm,
          act_mem_banks_bank_a_31_447_416_sva_dfm, while_mux_53_ssc_mx0);
      act_mem_banks_read_for_mux_1_itm <= MUX_v_32_32_2(act_mem_banks_bank_a_0_479_448_sva_dfm,
          act_mem_banks_bank_a_1_479_448_sva_dfm, act_mem_banks_bank_a_2_479_448_sva_dfm,
          act_mem_banks_bank_a_3_479_448_sva_dfm, act_mem_banks_bank_a_4_479_448_sva_dfm,
          act_mem_banks_bank_a_5_479_448_sva_dfm, act_mem_banks_bank_a_6_479_448_sva_dfm,
          act_mem_banks_bank_a_7_479_448_sva_dfm, act_mem_banks_bank_a_8_479_448_sva_dfm,
          act_mem_banks_bank_a_9_479_448_sva_dfm, act_mem_banks_bank_a_10_479_448_sva_dfm,
          act_mem_banks_bank_a_11_479_448_sva_dfm, act_mem_banks_bank_a_12_479_448_sva_dfm,
          act_mem_banks_bank_a_13_479_448_sva_dfm, act_mem_banks_bank_a_14_479_448_sva_dfm,
          act_mem_banks_bank_a_15_479_448_sva_dfm, act_mem_banks_bank_a_16_479_448_sva_dfm,
          act_mem_banks_bank_a_17_479_448_sva_dfm, act_mem_banks_bank_a_18_479_448_sva_dfm,
          act_mem_banks_bank_a_19_479_448_sva_dfm, act_mem_banks_bank_a_20_479_448_sva_dfm,
          act_mem_banks_bank_a_21_479_448_sva_dfm, act_mem_banks_bank_a_22_479_448_sva_dfm,
          act_mem_banks_bank_a_23_479_448_sva_dfm, act_mem_banks_bank_a_24_479_448_sva_dfm,
          act_mem_banks_bank_a_25_479_448_sva_dfm, act_mem_banks_bank_a_26_479_448_sva_dfm,
          act_mem_banks_bank_a_27_479_448_sva_dfm, act_mem_banks_bank_a_28_479_448_sva_dfm,
          act_mem_banks_bank_a_29_479_448_sva_dfm, act_mem_banks_bank_a_30_479_448_sva_dfm,
          act_mem_banks_bank_a_31_479_448_sva_dfm, while_mux_53_ssc_mx0);
      act_mem_banks_read_for_mux_itm <= MUX_v_32_32_2(act_mem_banks_bank_a_0_511_480_sva_dfm,
          act_mem_banks_bank_a_1_511_480_sva_dfm, act_mem_banks_bank_a_2_511_480_sva_dfm,
          act_mem_banks_bank_a_3_511_480_sva_dfm, act_mem_banks_bank_a_4_511_480_sva_dfm,
          act_mem_banks_bank_a_5_511_480_sva_dfm, act_mem_banks_bank_a_6_511_480_sva_dfm,
          act_mem_banks_bank_a_7_511_480_sva_dfm, act_mem_banks_bank_a_8_511_480_sva_dfm,
          act_mem_banks_bank_a_9_511_480_sva_dfm, act_mem_banks_bank_a_10_511_480_sva_dfm,
          act_mem_banks_bank_a_11_511_480_sva_dfm, act_mem_banks_bank_a_12_511_480_sva_dfm,
          act_mem_banks_bank_a_13_511_480_sva_dfm, act_mem_banks_bank_a_14_511_480_sva_dfm,
          act_mem_banks_bank_a_15_511_480_sva_dfm, act_mem_banks_bank_a_16_511_480_sva_dfm,
          act_mem_banks_bank_a_17_511_480_sva_dfm, act_mem_banks_bank_a_18_511_480_sva_dfm,
          act_mem_banks_bank_a_19_511_480_sva_dfm, act_mem_banks_bank_a_20_511_480_sva_dfm,
          act_mem_banks_bank_a_21_511_480_sva_dfm, act_mem_banks_bank_a_22_511_480_sva_dfm,
          act_mem_banks_bank_a_23_511_480_sva_dfm, act_mem_banks_bank_a_24_511_480_sva_dfm,
          act_mem_banks_bank_a_25_511_480_sva_dfm, act_mem_banks_bank_a_26_511_480_sva_dfm,
          act_mem_banks_bank_a_27_511_480_sva_dfm, act_mem_banks_bank_a_28_511_480_sva_dfm,
          act_mem_banks_bank_a_29_511_480_sva_dfm, act_mem_banks_bank_a_30_511_480_sva_dfm,
          act_mem_banks_bank_a_31_511_480_sva_dfm, while_mux_53_ssc_mx0);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_0_sva_dfm_3 <= 1'b0;
      rva_out_reg_data_8_sva_dfm_3 <= 1'b0;
      rva_out_reg_data_29_24_sva_dfm_3_5_4 <= 2'b00;
      rva_out_reg_data_39_32_sva_dfm_3_7_4 <= 4'b0000;
      rva_out_reg_data_52_48_sva_dfm_3 <= 5'b00000;
      rva_out_reg_data_71_64_sva_dfm_3_7_5 <= 3'b000;
      rva_out_reg_data_71_64_sva_dfm_3_4_0 <= 5'b00000;
      rva_out_reg_data_29_24_sva_dfm_3_3 <= 1'b0;
      rva_out_reg_data_29_24_sva_dfm_3_2_0 <= 3'b000;
      rva_out_reg_data_39_32_sva_dfm_3_3 <= 1'b0;
      rva_out_reg_data_39_32_sva_dfm_3_2_0 <= 3'b000;
    end
    else if ( rva_out_reg_data_and_62_cse ) begin
      rva_out_reg_data_0_sva_dfm_3 <= MUX_s_1_2_2(ActUnit_DecodeAxi_mux_93_nl, ActUnit_PushOutput_if_for_and_stg_2_7_sva,
          is_start_sva);
      rva_out_reg_data_8_sva_dfm_3 <= MUX_s_1_2_2(ActUnit_DecodeAxi_mux_94_nl, Gelu_for_and_2_cse_sva,
          is_start_sva);
      rva_out_reg_data_29_24_sva_dfm_3_5_4 <= MUX1HOT_v_2_4_2(rva_out_reg_data_29_24_sva_dfm_6_5_4,
          (act_config_num_inst_sva[5:4]), (act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_20_itm[5:4]),
          (act_config_inst_regs_3_sva_dfm_5[5:4]), {while_asn_2035 , while_asn_2037
          , while_and_282_cse , while_and_283_cse});
      rva_out_reg_data_39_32_sva_dfm_3_7_4 <= MUX1HOT_v_4_4_2(rva_out_reg_data_39_32_sva_dfm_6_7_4,
          (act_config_num_output_sva[7:4]), (act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_21_itm[7:4]),
          (act_config_inst_regs_4_sva_dfm_5[7:4]), {while_asn_2035 , while_asn_2037
          , while_and_282_cse , while_and_283_cse});
      rva_out_reg_data_52_48_sva_dfm_3 <= MUX1HOT_v_5_4_2(ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_1_30_26,
          act_config_buffer_addr_base_sva, act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_22_nl,
          (act_config_inst_regs_6_sva_dfm_5[4:0]), {while_asn_2035 , while_asn_2037
          , while_and_282_cse , while_and_283_cse});
      rva_out_reg_data_71_64_sva_dfm_3_7_5 <= MUX1HOT_v_3_4_2(rva_out_reg_data_71_64_sva_dfm_6_7_5,
          (act_config_output_addr_base_sva[7:5]), (act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_23_itm[7:5]),
          (act_config_inst_regs_8_sva_dfm_5[7:5]), {while_asn_2035 , while_asn_2037
          , while_and_282_cse , while_and_283_cse});
      rva_out_reg_data_71_64_sva_dfm_3_4_0 <= MUX1HOT_v_5_4_2(rva_out_reg_data_71_64_sva_dfm_6_4_0,
          (act_config_output_addr_base_sva[4:0]), (act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_23_itm[4:0]),
          (act_config_inst_regs_8_sva_dfm_5[4:0]), {while_asn_2035 , while_asn_2037
          , while_and_282_cse , while_and_283_cse});
      rva_out_reg_data_29_24_sva_dfm_3_3 <= MUX1HOT_s_1_4_2(rva_out_reg_data_29_24_sva_dfm_6_3,
          (act_config_num_inst_sva[3]), (act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_20_itm[3]),
          (act_config_inst_regs_3_sva_dfm_5[3]), {while_asn_2035 , while_asn_2037
          , while_and_282_cse , while_and_283_cse});
      rva_out_reg_data_29_24_sva_dfm_3_2_0 <= MUX1HOT_v_3_4_2(rva_out_reg_data_29_24_sva_dfm_6_2_0,
          (act_config_num_inst_sva[2:0]), (act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_20_itm[2:0]),
          (act_config_inst_regs_3_sva_dfm_5[2:0]), {while_asn_2035 , while_asn_2037
          , while_and_282_cse , while_and_283_cse});
      rva_out_reg_data_39_32_sva_dfm_3_3 <= MUX1HOT_s_1_4_2(rva_out_reg_data_39_32_sva_dfm_6_3,
          (act_config_num_output_sva[3]), (act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_21_itm[3]),
          (act_config_inst_regs_4_sva_dfm_5[3]), {while_asn_2035 , while_asn_2037
          , while_and_282_cse , while_and_283_cse});
      rva_out_reg_data_39_32_sva_dfm_3_2_0 <= MUX1HOT_v_3_4_2(rva_out_reg_data_39_32_sva_dfm_6_2_0,
          (act_config_num_output_sva[2:0]), (act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_21_itm[2:0]),
          (act_config_inst_regs_4_sva_dfm_5[2:0]), {while_asn_2035 , while_asn_2037
          , while_and_282_cse , while_and_283_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      w_axi_rsp_lpi_1_dfm_1 <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~((~ and_2371_cse) | or_dcpl_457)) ) begin
      w_axi_rsp_lpi_1_dfm_1 <= ~(ActUnit_DecodeAxi_rva_in_reg_rw_sva_mx1 | (~ ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_return_sva_mx1)
          | is_start_sva);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_RunInst_case_3_act_port_reg_data_sva <= 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( act_write_data_data_and_15_cse & (~((~ (act_config_in_InstFetch_return_sva_7_2[2]))
        | (act_config_in_InstFetch_return_sva_7_2[5]) | (~ act_port_PopNB_mioi_return_rsc_z_mxwt)
        | (act_config_in_InstFetch_return_sva_7_2[4:3]!=2'b01))) & is_start_sva &
        ActUnit_RunInst_switch_lp_equal_tmp_2 ) begin
      ActUnit_RunInst_case_3_act_port_reg_data_sva <= act_port_PopNB_mioi_data_data_rsc_z_mxwt;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_config_inst_counter_sva_dfm_3 <= 5'b00000;
    end
    else if ( ActUnitRun_wen & ((rva_in_PopNB_mioi_return_rsc_z_mxwt & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
        & and_dcpl_1072 & and_dcpl_1228) | and_dcpl_1262) ) begin
      act_config_inst_counter_sva_dfm_3 <= MUX_v_5_2_2(({{4{ActUnit_DecodeAxiRead_unequal_tmp_1}},
          ActUnit_DecodeAxiRead_unequal_tmp_1}), act_config_inst_counter_sva, or_dcpl_1014);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_output_counter_sva_dfm_3_ftd <= 4'b0000;
      reg_act_config_output_counter_sva_dfm_3_ftd_1_3 <= 1'b0;
      reg_act_config_output_counter_sva_dfm_3_ftd_1_2_0 <= 3'b000;
      is_incr_lpi_1_dfm_1 <= 1'b0;
      act_config_is_zero_first_sva_dfm_4 <= 1'b0;
    end
    else if ( act_config_output_counter_and_1_cse ) begin
      reg_act_config_output_counter_sva_dfm_3_ftd <= MUX_v_4_2_2(({{3{ActUnit_DecodeAxiRead_unequal_tmp_1}},
          ActUnit_DecodeAxiRead_unequal_tmp_1}), act_config_output_counter_sva_7_4,
          or_dcpl_1014);
      reg_act_config_output_counter_sva_dfm_3_ftd_1_3 <= MUX_s_1_2_2(ActUnit_DecodeAxiRead_unequal_tmp_1,
          act_config_output_counter_sva_3, or_dcpl_1014);
      reg_act_config_output_counter_sva_dfm_3_ftd_1_2_0 <= MUX_v_3_2_2(({{2{ActUnit_DecodeAxiRead_unequal_tmp_1}},
          ActUnit_DecodeAxiRead_unequal_tmp_1}), act_config_output_counter_sva_2_0,
          or_dcpl_1014);
      is_incr_lpi_1_dfm_1 <= act_port_PopNB_mioi_return_rsc_z_mxwt | (~ ActUnit_RunInst_switch_lp_equal_tmp_2)
          | (~ is_start_sva);
      act_config_is_zero_first_sva_dfm_4 <= MUX_s_1_2_2(ActUnit_DecodeAxiWrite_mux_4_nl,
          act_config_is_zero_first_sva, and_dcpl_1262);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_y_1_sva_3_24_22 <= 3'b000;
    end
    else if ( ActUnitRun_wen & and_dcpl_9 & (~ (act_config_in_InstFetch_return_sva_7_2[2]))
        & Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
        & Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
        & Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
        & (~ operator_32_8_true_AC_TRN_AC_WRAP_3_less_15_tmp) ) begin
      Silu_for_y_1_sva_3_24_22 <= Silu_for_1_else_else_else_if_acc_itm_25_1_1[24:22];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_y_1_sva_3_21_0 <= 22'b0000000000000000000000;
    end
    else if ( and_1864_tmp ) begin
      Silu_for_y_1_sva_3_21_0 <= MUX_v_22_2_2(and_1749_nl, (Silu_for_1_else_else_else_if_acc_itm_25_1_1[21:0]),
          mux_448_itm);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_2_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_24_22
          <= 3'b000;
    end
    else if ( ActUnitRun_wen & and_dcpl_9 & (~ (act_config_in_InstFetch_return_sva_7_2[2]))
        & Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
        & Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
        & Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
        & (~ operator_32_8_true_AC_TRN_AC_WRAP_3_less_14_tmp) ) begin
      Silu_for_2_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_24_22
          <= Silu_for_2_else_else_else_if_acc_itm_25_1_1[24:22];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_2_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0
          <= 22'b0000000000000000000000;
    end
    else if ( and_1865_tmp ) begin
      Silu_for_2_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0
          <= MUX_v_22_2_2((Silu_for_2_else_else_else_if_acc_itm_25_1_1[21:0]), and_1752_nl,
          not_tmp_495);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_3_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_24_22
          <= 3'b000;
    end
    else if ( ActUnitRun_wen & and_dcpl_9 & (~ (act_config_in_InstFetch_return_sva_7_2[2]))
        & Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
        & Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
        & Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
        & (~ operator_32_8_true_AC_TRN_AC_WRAP_3_less_13_tmp) ) begin
      Silu_for_3_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_24_22
          <= Silu_for_3_else_else_else_if_acc_itm_25_1_1[24:22];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_3_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0
          <= 22'b0000000000000000000000;
    end
    else if ( and_1867_tmp ) begin
      Silu_for_3_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0
          <= MUX_v_22_2_2(and_1756_nl, (Silu_for_3_else_else_else_if_acc_itm_25_1_1[21:0]),
          mux_448_itm);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_4_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_24_22
          <= 3'b000;
    end
    else if ( ActUnitRun_wen & and_dcpl_9 & (~ (act_config_in_InstFetch_return_sva_7_2[2]))
        & Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
        & Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
        & Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
        & (~ operator_32_8_true_AC_TRN_AC_WRAP_3_less_12_tmp) ) begin
      Silu_for_4_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_24_22
          <= Silu_for_4_else_else_else_if_acc_itm_25_1_1[24:22];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_4_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0
          <= 22'b0000000000000000000000;
    end
    else if ( and_1869_tmp ) begin
      Silu_for_4_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0
          <= MUX_v_22_2_2(and_1759_nl, (Silu_for_4_else_else_else_if_acc_itm_25_1_1[21:0]),
          mux_448_itm);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_5_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_24_22
          <= 3'b000;
    end
    else if ( ActUnitRun_wen & and_dcpl_9 & (~ (act_config_in_InstFetch_return_sva_7_2[2]))
        & Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
        & Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
        & Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
        & (~ operator_32_8_true_AC_TRN_AC_WRAP_3_less_11_tmp) ) begin
      Silu_for_5_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_24_22
          <= Silu_for_5_else_else_else_if_acc_itm_25_1_1[24:22];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_5_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0
          <= 22'b0000000000000000000000;
    end
    else if ( and_1871_tmp ) begin
      Silu_for_5_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0
          <= MUX_v_22_2_2(and_1762_nl, (Silu_for_5_else_else_else_if_acc_itm_25_1_1[21:0]),
          mux_448_itm);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_6_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_24_22
          <= 3'b000;
    end
    else if ( ActUnitRun_wen & and_dcpl_9 & (~ (act_config_in_InstFetch_return_sva_7_2[2]))
        & Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
        & Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
        & Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
        & (~ operator_32_8_true_AC_TRN_AC_WRAP_3_less_10_tmp) ) begin
      Silu_for_6_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_24_22
          <= Silu_for_6_else_else_else_if_acc_itm_25_1_1[24:22];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_6_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0
          <= 22'b0000000000000000000000;
    end
    else if ( and_1873_tmp ) begin
      Silu_for_6_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0
          <= MUX_v_22_2_2(and_1765_nl, (Silu_for_6_else_else_else_if_acc_itm_25_1_1[21:0]),
          mux_448_itm);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_7_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_24_22
          <= 3'b000;
    end
    else if ( ActUnitRun_wen & and_dcpl_9 & (~ (act_config_in_InstFetch_return_sva_7_2[2]))
        & Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
        & Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
        & Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
        & (~ operator_32_8_true_AC_TRN_AC_WRAP_3_less_9_tmp) ) begin
      Silu_for_7_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_24_22
          <= Silu_for_7_else_else_else_if_acc_itm_25_1_1[24:22];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_7_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0
          <= 22'b0000000000000000000000;
    end
    else if ( and_1875_tmp ) begin
      Silu_for_7_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0
          <= MUX_v_22_2_2(and_1768_nl, (Silu_for_7_else_else_else_if_acc_itm_25_1_1[21:0]),
          mux_448_itm);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_y_8_sva_3_24_22 <= 3'b000;
    end
    else if ( ActUnitRun_wen & and_dcpl_9 & (~ (act_config_in_InstFetch_return_sva_7_2[2]))
        & Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
        & Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
        & Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
        & (~ operator_32_8_true_AC_TRN_AC_WRAP_3_less_8_tmp) ) begin
      Silu_for_y_8_sva_3_24_22 <= Silu_for_8_else_else_else_if_acc_itm_25_1_1[24:22];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_y_8_sva_3_21_0 <= 22'b0000000000000000000000;
    end
    else if ( and_1877_tmp ) begin
      Silu_for_y_8_sva_3_21_0 <= MUX_v_22_2_2(and_1771_nl, (Silu_for_8_else_else_else_if_acc_itm_25_1_1[21:0]),
          mux_448_itm);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_9_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_24_22
          <= 3'b000;
    end
    else if ( act_write_data_data_and_15_cse & and_dcpl_9 & (~ (act_config_in_InstFetch_return_sva_7_2[2]))
        & Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
        & Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
        & Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
        & (~ operator_32_8_true_AC_TRN_AC_WRAP_3_less_7_tmp) ) begin
      Silu_for_9_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_24_22
          <= Silu_for_9_else_else_else_if_acc_itm_25_1_1[24:22];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_9_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0
          <= 22'b0000000000000000000000;
    end
    else if ( and_1879_tmp ) begin
      Silu_for_9_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0
          <= MUX_v_22_2_2(and_1774_nl, (Silu_for_9_else_else_else_if_acc_itm_25_1_1[21:0]),
          mux_448_itm);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
          <= 1'b0;
    end
    else if ( act_write_data_data_and_15_cse & mux_125_nl & and_dcpl_43 ) begin
      Gelu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
          <= MUX_s_1_2_2((27'b100000000000000000000000000 < ({reg_ActUnit_RunInst_case_14_nv_scvector_cctor_data_0_ftd_1_30_26
          , reg_ActUnit_RunInst_case_14_nv_scvector_cctor_data_0_1_ftd_rsp_0 , reg_ActUnit_RunInst_case_14_nv_scvector_cctor_data_0_1_ftd_rsp_1
          , reg_ActUnit_RunInst_case_14_nv_scvector_cctor_data_0_1_ftd_1})), operator_32_8_true_AC_TRN_AC_WRAP_7_less_15_tmp,
          act_config_in_InstFetch_return_sva_7_2[2]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
          <= 1'b0;
    end
    else if ( act_write_data_data_and_15_cse & mux_126_nl & and_dcpl_43 ) begin
      Gelu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
          <= MUX_s_1_2_2(operator_32_8_true_AC_TRN_AC_WRAP_3_less_15_tmp, operator_32_8_true_AC_TRN_AC_WRAP_6_less_15_tmp,
          act_config_in_InstFetch_return_sva_7_2[2]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
          <= 1'b0;
    end
    else if ( act_write_data_data_and_15_cse & mux_127_nl & and_dcpl_43 ) begin
      Gelu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
          <= MUX_s_1_2_2((27'b100000000000000000000000000 < ({reg_nv_scvector_cctor_nv_scvector_5_for_2_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          , reg_nv_scvector_cctor_nv_scvector_5_for_2_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          , reg_nv_scvector_cctor_nv_scvector_5_for_2_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          , reg_nv_scvector_cctor_nv_scvector_5_for_2_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1})),
          operator_32_8_true_AC_TRN_AC_WRAP_7_less_14_tmp, act_config_in_InstFetch_return_sva_7_2[2]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
          <= 1'b0;
    end
    else if ( act_write_data_data_and_15_cse & mux_128_nl & and_dcpl_43 ) begin
      Gelu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
          <= MUX_s_1_2_2(operator_32_8_true_AC_TRN_AC_WRAP_3_less_14_tmp, operator_32_8_true_AC_TRN_AC_WRAP_6_less_14_tmp,
          act_config_in_InstFetch_return_sva_7_2[2]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
          <= 1'b0;
    end
    else if ( act_write_data_data_and_15_cse & mux_129_nl & and_dcpl_43 ) begin
      Gelu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
          <= MUX_s_1_2_2((27'b100000000000000000000000000 < ({reg_nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          , reg_nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          , reg_nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          , reg_nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1})),
          operator_32_8_true_AC_TRN_AC_WRAP_7_less_13_tmp, act_config_in_InstFetch_return_sva_7_2[2]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
          <= 1'b0;
    end
    else if ( act_write_data_data_and_15_cse & mux_130_nl & and_dcpl_43 ) begin
      Gelu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
          <= MUX_s_1_2_2(operator_32_8_true_AC_TRN_AC_WRAP_3_less_13_tmp, operator_32_8_true_AC_TRN_AC_WRAP_6_less_13_tmp,
          act_config_in_InstFetch_return_sva_7_2[2]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
          <= 1'b0;
    end
    else if ( act_write_data_data_and_15_cse & mux_131_nl & and_dcpl_43 ) begin
      Gelu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
          <= MUX_s_1_2_2((27'b100000000000000000000000000 < ({reg_nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          , reg_nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          , reg_nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          , reg_nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1})),
          operator_32_8_true_AC_TRN_AC_WRAP_7_less_12_tmp, act_config_in_InstFetch_return_sva_7_2[2]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
          <= 1'b0;
    end
    else if ( act_write_data_data_and_15_cse & mux_132_nl & and_dcpl_43 ) begin
      Gelu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
          <= MUX_s_1_2_2(operator_32_8_true_AC_TRN_AC_WRAP_3_less_12_tmp, operator_32_8_true_AC_TRN_AC_WRAP_6_less_12_tmp,
          act_config_in_InstFetch_return_sva_7_2[2]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
          <= 1'b0;
    end
    else if ( act_write_data_data_and_15_cse & mux_133_nl & and_dcpl_43 ) begin
      Gelu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
          <= MUX_s_1_2_2((27'b100000000000000000000000000 < ({reg_nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          , reg_nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          , reg_nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          , reg_nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1})),
          operator_32_8_true_AC_TRN_AC_WRAP_7_less_11_tmp, act_config_in_InstFetch_return_sva_7_2[2]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
          <= 1'b0;
    end
    else if ( act_write_data_data_and_15_cse & mux_134_nl & and_dcpl_43 ) begin
      Gelu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
          <= MUX_s_1_2_2(operator_32_8_true_AC_TRN_AC_WRAP_3_less_11_tmp, operator_32_8_true_AC_TRN_AC_WRAP_6_less_11_tmp,
          act_config_in_InstFetch_return_sva_7_2[2]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
          <= 1'b0;
    end
    else if ( act_write_data_data_and_15_cse & mux_135_nl & and_dcpl_43 ) begin
      Gelu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
          <= MUX_s_1_2_2((27'b100000000000000000000000000 < ({reg_nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          , reg_nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          , reg_nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          , reg_nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1})),
          operator_32_8_true_AC_TRN_AC_WRAP_7_less_10_tmp, act_config_in_InstFetch_return_sva_7_2[2]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
          <= 1'b0;
    end
    else if ( act_write_data_data_and_15_cse & mux_136_nl & and_dcpl_43 ) begin
      Gelu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
          <= MUX_s_1_2_2(operator_32_8_true_AC_TRN_AC_WRAP_3_less_10_tmp, operator_32_8_true_AC_TRN_AC_WRAP_6_less_10_tmp,
          act_config_in_InstFetch_return_sva_7_2[2]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
          <= 1'b0;
    end
    else if ( act_write_data_data_and_15_cse & mux_137_nl & and_dcpl_43 ) begin
      Gelu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
          <= MUX_s_1_2_2((27'b100000000000000000000000000 < ({reg_nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          , reg_nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          , reg_nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          , reg_nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1})),
          operator_32_8_true_AC_TRN_AC_WRAP_7_less_9_tmp, act_config_in_InstFetch_return_sva_7_2[2]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
          <= 1'b0;
    end
    else if ( act_write_data_data_and_15_cse & mux_138_nl & and_dcpl_43 ) begin
      Gelu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
          <= MUX_s_1_2_2(operator_32_8_true_AC_TRN_AC_WRAP_3_less_9_tmp, operator_32_8_true_AC_TRN_AC_WRAP_6_less_9_tmp,
          act_config_in_InstFetch_return_sva_7_2[2]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
          <= 1'b0;
    end
    else if ( act_write_data_data_and_15_cse & mux_139_nl & and_dcpl_43 ) begin
      Gelu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
          <= MUX_s_1_2_2((27'b100000000000000000000000000 < ({reg_nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          , reg_nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          , reg_nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          , reg_nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1})),
          operator_32_8_true_AC_TRN_AC_WRAP_7_less_8_tmp, act_config_in_InstFetch_return_sva_7_2[2]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
          <= 1'b0;
    end
    else if ( act_write_data_data_and_15_cse & mux_140_nl & and_dcpl_43 ) begin
      Gelu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
          <= MUX_s_1_2_2(operator_32_8_true_AC_TRN_AC_WRAP_3_less_8_tmp, operator_32_8_true_AC_TRN_AC_WRAP_6_less_8_tmp,
          act_config_in_InstFetch_return_sva_7_2[2]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
          <= 1'b0;
    end
    else if ( act_write_data_data_and_15_cse & mux_141_nl & and_dcpl_43 ) begin
      Gelu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
          <= MUX_s_1_2_2((27'b100000000000000000000000000 < ({reg_nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          , reg_nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          , reg_nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          , reg_nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1})),
          operator_32_8_true_AC_TRN_AC_WRAP_7_less_7_tmp, act_config_in_InstFetch_return_sva_7_2[2]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
          <= 1'b0;
    end
    else if ( act_write_data_data_and_15_cse & mux_142_nl & and_dcpl_43 ) begin
      Gelu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
          <= MUX_s_1_2_2(operator_32_8_true_AC_TRN_AC_WRAP_3_less_7_tmp, operator_32_8_true_AC_TRN_AC_WRAP_6_less_7_tmp,
          act_config_in_InstFetch_return_sva_7_2[2]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
          <= 1'b0;
    end
    else if ( act_write_data_data_and_15_cse & mux_143_nl & and_dcpl_43 ) begin
      Gelu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
          <= MUX_s_1_2_2((27'b100000000000000000000000000 < ({reg_nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          , reg_nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          , reg_nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          , reg_nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1})),
          operator_32_8_true_AC_TRN_AC_WRAP_7_less_6_tmp, act_config_in_InstFetch_return_sva_7_2[2]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
          <= 1'b0;
    end
    else if ( act_write_data_data_and_15_cse & mux_144_nl & and_dcpl_43 ) begin
      Gelu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
          <= MUX_s_1_2_2(operator_32_8_true_AC_TRN_AC_WRAP_3_less_6_tmp, operator_32_8_true_AC_TRN_AC_WRAP_6_less_6_tmp,
          act_config_in_InstFetch_return_sva_7_2[2]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
          <= 1'b0;
    end
    else if ( act_write_data_data_and_15_cse & mux_145_nl & and_dcpl_43 ) begin
      Gelu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
          <= MUX_s_1_2_2((27'b100000000000000000000000000 < ({reg_nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          , reg_nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          , reg_nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          , reg_nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1})),
          operator_32_8_true_AC_TRN_AC_WRAP_7_less_5_tmp, act_config_in_InstFetch_return_sva_7_2[2]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
          <= 1'b0;
    end
    else if ( act_write_data_data_and_15_cse & mux_146_nl & and_dcpl_43 ) begin
      Gelu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
          <= MUX_s_1_2_2(operator_32_8_true_AC_TRN_AC_WRAP_3_less_5_tmp, operator_32_8_true_AC_TRN_AC_WRAP_6_less_5_tmp,
          act_config_in_InstFetch_return_sva_7_2[2]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
          <= 1'b0;
    end
    else if ( act_write_data_data_and_15_cse & mux_147_nl & and_dcpl_43 ) begin
      Gelu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
          <= MUX_s_1_2_2((27'b100000000000000000000000000 < ({reg_nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          , reg_nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          , reg_nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          , reg_nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1})),
          operator_32_8_true_AC_TRN_AC_WRAP_7_less_4_tmp, act_config_in_InstFetch_return_sva_7_2[2]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
          <= 1'b0;
    end
    else if ( act_write_data_data_and_15_cse & mux_148_nl & and_dcpl_43 ) begin
      Gelu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
          <= MUX_s_1_2_2(operator_32_8_true_AC_TRN_AC_WRAP_3_less_4_tmp, operator_32_8_true_AC_TRN_AC_WRAP_6_less_4_tmp,
          act_config_in_InstFetch_return_sva_7_2[2]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
          <= 1'b0;
    end
    else if ( act_write_data_data_and_15_cse & mux_149_nl & and_dcpl_43 ) begin
      Gelu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
          <= MUX_s_1_2_2((27'b100000000000000000000000000 < ({reg_nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          , reg_nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          , reg_nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          , reg_nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1})),
          operator_32_8_true_AC_TRN_AC_WRAP_7_less_3_tmp, act_config_in_InstFetch_return_sva_7_2[2]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
          <= 1'b0;
    end
    else if ( act_write_data_data_and_15_cse & mux_150_nl & and_dcpl_43 ) begin
      Gelu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
          <= MUX_s_1_2_2(operator_32_8_true_AC_TRN_AC_WRAP_3_less_3_tmp, operator_32_8_true_AC_TRN_AC_WRAP_6_less_3_tmp,
          act_config_in_InstFetch_return_sva_7_2[2]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
          <= 1'b0;
    end
    else if ( act_write_data_data_and_15_cse & mux_151_nl & and_dcpl_43 ) begin
      Gelu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
          <= MUX_s_1_2_2((27'b100000000000000000000000000 < ({reg_nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          , reg_nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          , reg_nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          , reg_nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1})),
          operator_32_8_true_AC_TRN_AC_WRAP_7_less_2_tmp, act_config_in_InstFetch_return_sva_7_2[2]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
          <= 1'b0;
    end
    else if ( act_write_data_data_and_15_cse & mux_152_nl & and_dcpl_43 ) begin
      Gelu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
          <= MUX_s_1_2_2(operator_32_8_true_AC_TRN_AC_WRAP_3_less_2_tmp, operator_32_8_true_AC_TRN_AC_WRAP_6_less_2_tmp,
          act_config_in_InstFetch_return_sva_7_2[2]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
          <= 1'b0;
    end
    else if ( act_write_data_data_and_15_cse & mux_153_nl & and_dcpl_43 ) begin
      Gelu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
          <= MUX_s_1_2_2((27'b100000000000000000000000000 < ({reg_nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          , reg_nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          , reg_nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          , reg_nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1})),
          operator_32_8_true_AC_TRN_AC_WRAP_7_less_1_tmp, act_config_in_InstFetch_return_sva_7_2[2]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
          <= 1'b0;
    end
    else if ( act_write_data_data_and_15_cse & mux_154_nl & and_dcpl_43 ) begin
      Gelu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
          <= MUX_s_1_2_2(operator_32_8_true_AC_TRN_AC_WRAP_3_less_1_tmp, operator_32_8_true_AC_TRN_AC_WRAP_6_less_1_tmp,
          act_config_in_InstFetch_return_sva_7_2[2]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
          <= 1'b0;
    end
    else if ( act_write_data_data_and_15_cse & mux_155_nl & and_dcpl_43 ) begin
      Gelu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_7_slc_operator_32_8_true_AC_TRN_AC_WRAP_7_acc_31_svs
          <= MUX_s_1_2_2((27'b100000000000000000000000000 < ({reg_nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          , reg_nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          , reg_nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          , reg_nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1})),
          operator_32_8_true_AC_TRN_AC_WRAP_7_less_tmp, act_config_in_InstFetch_return_sva_7_2[2]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Gelu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
          <= 1'b0;
    end
    else if ( act_write_data_data_and_15_cse & mux_156_nl & and_dcpl_43 ) begin
      Gelu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_6_slc_operator_32_8_true_AC_TRN_AC_WRAP_6_acc_31_svs
          <= MUX_s_1_2_2(operator_32_8_true_AC_TRN_AC_WRAP_3_less_tmp, operator_32_8_true_AC_TRN_AC_WRAP_6_less_tmp,
          act_config_in_InstFetch_return_sva_7_2[2]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_get_slc_2U_NVUINT8_return_2_sva <= 2'b00;
    end
    else if ( ActUnitRun_wen & (~((~ and_2371_cse) & and_dcpl_1061)) & and_dcpl_469
        ) begin
      nvhls_get_slc_2U_NVUINT8_return_2_sva <= MUX_v_2_32_2((act_config_inst_regs_0_sva_dfm_5[3:2]),
          (act_config_inst_regs_1_sva_dfm_5[3:2]), (act_config_inst_regs_2_sva_dfm_5[3:2]),
          (act_config_inst_regs_3_sva_dfm_5[3:2]), (act_config_inst_regs_4_sva_dfm_5[3:2]),
          (act_config_inst_regs_5_sva_dfm_5[3:2]), (act_config_inst_regs_6_sva_dfm_5[3:2]),
          (act_config_inst_regs_7_sva_dfm_5[3:2]), (act_config_inst_regs_8_sva_dfm_5[3:2]),
          (act_config_inst_regs_9_sva_dfm_5[3:2]), (act_config_inst_regs_10_sva_dfm_5[3:2]),
          (act_config_inst_regs_11_sva_dfm_5[3:2]), (act_config_inst_regs_12_sva_dfm_5[3:2]),
          (act_config_inst_regs_13_sva_dfm_5[3:2]), (act_config_inst_regs_14_sva_dfm_5[3:2]),
          (act_config_inst_regs_15_sva_dfm_5[3:2]), ActUnit_DecodeAxiWrite_if_mux_5_nl,
          ActUnit_DecodeAxiWrite_if_mux_7_nl, ActUnit_DecodeAxiWrite_if_mux_9_nl,
          ActUnit_DecodeAxiWrite_if_mux_11_nl, ActUnit_DecodeAxiWrite_if_mux_13_nl,
          ActUnit_DecodeAxiWrite_if_mux_15_nl, ActUnit_DecodeAxiWrite_if_mux_17_nl,
          ActUnit_DecodeAxiWrite_if_mux_19_nl, ActUnit_DecodeAxiWrite_if_mux_21_nl,
          ActUnit_DecodeAxiWrite_if_mux_23_nl, ActUnit_DecodeAxiWrite_if_mux_25_nl,
          ActUnit_DecodeAxiWrite_if_mux_27_nl, ActUnit_DecodeAxiWrite_if_mux_29_nl,
          ActUnit_DecodeAxiWrite_if_mux_31_nl, ActUnit_DecodeAxiWrite_if_mux_33_nl,
          ActUnit_DecodeAxiWrite_if_mux_35_nl, act_config_inst_counter_sva);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_15_sva_8_31 <= 1'b0;
      act_regs_data_3_14_sva_8_31 <= 1'b0;
      act_regs_data_3_13_sva_8_31 <= 1'b0;
      act_regs_data_3_12_sva_8_31 <= 1'b0;
      act_regs_data_3_11_sva_8_31 <= 1'b0;
      act_regs_data_3_10_sva_8_31 <= 1'b0;
      act_regs_data_3_9_sva_8_31 <= 1'b0;
      act_regs_data_3_8_sva_8_31 <= 1'b0;
      act_regs_data_3_7_sva_8_31 <= 1'b0;
      act_regs_data_3_6_sva_8_31 <= 1'b0;
      act_regs_data_3_5_sva_8_31 <= 1'b0;
      act_regs_data_3_4_sva_8_31 <= 1'b0;
      act_regs_data_3_3_sva_8_31 <= 1'b0;
      act_regs_data_3_2_sva_8_31 <= 1'b0;
      act_regs_data_3_1_sva_8_31 <= 1'b0;
    end
    else if ( act_regs_data_and_832_cse ) begin
      act_regs_data_3_15_sva_8_31 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_3_15_sva_dfm_2_31, or_dcpl_850);
      act_regs_data_3_14_sva_8_31 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_3_14_sva_dfm_2_31, or_dcpl_852);
      act_regs_data_3_13_sva_8_31 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_3_13_sva_dfm_2_31, or_dcpl_855);
      act_regs_data_3_12_sva_8_31 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_3_12_sva_dfm_2_31, or_dcpl_857);
      act_regs_data_3_11_sva_8_31 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_3_11_sva_dfm_2_31, or_dcpl_860);
      act_regs_data_3_10_sva_8_31 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_3_10_sva_dfm_2_31, or_dcpl_862);
      act_regs_data_3_9_sva_8_31 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_3_9_sva_dfm_2_31, or_dcpl_865);
      act_regs_data_3_8_sva_8_31 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_3_8_sva_dfm_2_31, or_dcpl_867);
      act_regs_data_3_7_sva_8_31 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_3_7_sva_dfm_2_31, or_dcpl_869);
      act_regs_data_3_6_sva_8_31 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_3_6_sva_dfm_2_31, or_dcpl_870);
      act_regs_data_3_5_sva_8_31 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_3_5_sva_dfm_2_31, or_dcpl_871);
      act_regs_data_3_4_sva_8_31 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_3_4_sva_dfm_2_31, or_dcpl_872);
      act_regs_data_3_3_sva_8_31 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_3_3_sva_dfm_2_31, or_dcpl_873);
      act_regs_data_3_2_sva_8_31 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_3_2_sva_dfm_2_31, or_dcpl_874);
      act_regs_data_3_1_sva_8_31 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          act_regs_data_3_1_sva_dfm_2_31, or_dcpl_875);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_15_sva_8_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2704_enex5 ) begin
      act_regs_data_3_15_sva_8_30_26 <= MUX_v_5_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_3_15_sva_dfm_2_30_26, or_dcpl_850);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_15_sva_8_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2706_enex5 ) begin
      act_regs_data_3_15_sva_8_21_0 <= MUX_v_22_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_3_15_sva_dfm_2_21_0, or_dcpl_850);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_14_sva_8_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2707_enex5 ) begin
      act_regs_data_3_14_sva_8_30_26 <= MUX_v_5_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_3_14_sva_dfm_2_30_26, or_dcpl_852);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_14_sva_8_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2709_enex5 ) begin
      act_regs_data_3_14_sva_8_21_0 <= MUX_v_22_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_3_14_sva_dfm_2_21_0, or_dcpl_852);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_13_sva_8_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2710_enex5 ) begin
      act_regs_data_3_13_sva_8_30_26 <= MUX_v_5_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_3_13_sva_dfm_2_30_26, or_dcpl_855);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_13_sva_8_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2712_enex5 ) begin
      act_regs_data_3_13_sva_8_21_0 <= MUX_v_22_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_3_13_sva_dfm_2_21_0, or_dcpl_855);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_12_sva_8_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2713_enex5 ) begin
      act_regs_data_3_12_sva_8_30_26 <= MUX_v_5_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_3_12_sva_dfm_2_30_26, or_dcpl_857);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_12_sva_8_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2715_enex5 ) begin
      act_regs_data_3_12_sva_8_21_0 <= MUX_v_22_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_3_12_sva_dfm_2_21_0, or_dcpl_857);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_11_sva_8_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2716_enex5 ) begin
      act_regs_data_3_11_sva_8_30_26 <= MUX_v_5_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_3_11_sva_dfm_2_30_26, or_dcpl_860);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_11_sva_8_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2718_enex5 ) begin
      act_regs_data_3_11_sva_8_21_0 <= MUX_v_22_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_3_11_sva_dfm_2_21_0, or_dcpl_860);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_10_sva_8_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2719_enex5 ) begin
      act_regs_data_3_10_sva_8_30_26 <= MUX_v_5_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_3_10_sva_dfm_2_30_26, or_dcpl_862);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_10_sva_8_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2721_enex5 ) begin
      act_regs_data_3_10_sva_8_21_0 <= MUX_v_22_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_3_10_sva_dfm_2_21_0, or_dcpl_862);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_9_sva_8_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2722_enex5 ) begin
      act_regs_data_3_9_sva_8_30_26 <= MUX_v_5_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_3_9_sva_dfm_2_30_26, or_dcpl_865);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_9_sva_8_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2724_enex5 ) begin
      act_regs_data_3_9_sva_8_21_0 <= MUX_v_22_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_3_9_sva_dfm_2_21_0, or_dcpl_865);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_8_sva_8_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2725_enex5 ) begin
      act_regs_data_3_8_sva_8_30_26 <= MUX_v_5_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_3_8_sva_dfm_2_30_26, or_dcpl_867);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_8_sva_8_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2727_enex5 ) begin
      act_regs_data_3_8_sva_8_21_0 <= MUX_v_22_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_3_8_sva_dfm_2_21_0, or_dcpl_867);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_7_sva_8_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2728_enex5 ) begin
      act_regs_data_3_7_sva_8_30_26 <= MUX_v_5_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_3_7_sva_dfm_2_30_26, or_dcpl_869);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_7_sva_8_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2730_enex5 ) begin
      act_regs_data_3_7_sva_8_21_0 <= MUX_v_22_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_3_7_sva_dfm_2_21_0, or_dcpl_869);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_6_sva_8_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2731_enex5 ) begin
      act_regs_data_3_6_sva_8_30_26 <= MUX_v_5_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_3_6_sva_dfm_2_30_26, or_dcpl_870);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_6_sva_8_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2733_enex5 ) begin
      act_regs_data_3_6_sva_8_21_0 <= MUX_v_22_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_3_6_sva_dfm_2_21_0, or_dcpl_870);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_5_sva_8_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2734_enex5 ) begin
      act_regs_data_3_5_sva_8_30_26 <= MUX_v_5_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_3_5_sva_dfm_2_30_26, or_dcpl_871);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_5_sva_8_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2736_enex5 ) begin
      act_regs_data_3_5_sva_8_21_0 <= MUX_v_22_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_3_5_sva_dfm_2_21_0, or_dcpl_871);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_4_sva_8_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2737_enex5 ) begin
      act_regs_data_3_4_sva_8_30_26 <= MUX_v_5_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_3_4_sva_dfm_2_30_26, or_dcpl_872);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_4_sva_8_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2739_enex5 ) begin
      act_regs_data_3_4_sva_8_21_0 <= MUX_v_22_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_3_4_sva_dfm_2_21_0, or_dcpl_872);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_3_sva_8_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2740_enex5 ) begin
      act_regs_data_3_3_sva_8_30_26 <= MUX_v_5_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_3_3_sva_dfm_2_30_26, or_dcpl_873);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_3_sva_8_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2742_enex5 ) begin
      act_regs_data_3_3_sva_8_21_0 <= MUX_v_22_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_3_3_sva_dfm_2_21_0, or_dcpl_873);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_2_sva_8_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2743_enex5 ) begin
      act_regs_data_3_2_sva_8_30_26 <= MUX_v_5_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_3_2_sva_dfm_2_30_26, or_dcpl_874);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_2_sva_8_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2745_enex5 ) begin
      act_regs_data_3_2_sva_8_21_0 <= MUX_v_22_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_3_2_sva_dfm_2_21_0, or_dcpl_874);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_1_sva_8_30_26 <= 5'b00000;
    end
    else if ( act_regs_data_and_2746_enex5 ) begin
      act_regs_data_3_1_sva_8_30_26 <= MUX_v_5_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_3_1_sva_dfm_2_30_26, or_dcpl_875);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_1_sva_8_21_0 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2748_enex5 ) begin
      act_regs_data_3_1_sva_8_21_0 <= MUX_v_22_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_3_1_sva_dfm_2_21_0, or_dcpl_875);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_0_sva_8_31 <= 1'b0;
      act_regs_data_3_0_sva_8_30_26 <= 5'b00000;
      act_regs_data_3_0_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_3_0_sva_8_25 <= 1'b0;
      act_regs_data_3_0_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_124_cse ) begin
      act_regs_data_3_0_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_231_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_nl, and_dcpl_1246);
      act_regs_data_3_0_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_229_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_3_0_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_892_cse
          , act_regs_data_and_893_cse});
      act_regs_data_3_0_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_230_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_3_0_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_892_cse
          , act_regs_data_and_893_cse});
      act_regs_data_3_0_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_69_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_3_0_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_892_cse
          , act_regs_data_and_893_cse});
      act_regs_data_3_0_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_338_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_3_0_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_892_cse
          , act_regs_data_and_893_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_15_sva_8_31 <= 1'b0;
      act_regs_data_2_15_sva_8_30_26 <= 5'b00000;
      act_regs_data_2_15_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_2_15_sva_8_25 <= 1'b0;
      act_regs_data_2_15_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_128_cse ) begin
      act_regs_data_2_15_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_291_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_4_nl, and_dcpl_1246);
      act_regs_data_2_15_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_289_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_2_15_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_898_cse
          , act_regs_data_and_899_cse});
      act_regs_data_2_15_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_290_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_2_15_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_898_cse
          , act_regs_data_and_899_cse});
      act_regs_data_2_15_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_104_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_2_15_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_898_cse
          , act_regs_data_and_899_cse});
      act_regs_data_2_15_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_336_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_2_15_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_898_cse
          , act_regs_data_and_899_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_14_sva_8_31 <= 1'b0;
      act_regs_data_2_14_sva_8_30_26 <= 5'b00000;
      act_regs_data_2_14_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_2_14_sva_8_25 <= 1'b0;
      act_regs_data_2_14_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_132_cse ) begin
      act_regs_data_2_14_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_279_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_8_nl, and_dcpl_1246);
      act_regs_data_2_14_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_277_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_2_14_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_904_cse
          , act_regs_data_and_905_cse});
      act_regs_data_2_14_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_278_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_2_14_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_904_cse
          , act_regs_data_and_905_cse});
      act_regs_data_2_14_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_97_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_2_14_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_904_cse
          , act_regs_data_and_905_cse});
      act_regs_data_2_14_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_334_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_2_14_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_904_cse
          , act_regs_data_and_905_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_13_sva_8_31 <= 1'b0;
      act_regs_data_2_13_sva_8_30_26 <= 5'b00000;
      act_regs_data_2_13_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_2_13_sva_8_25 <= 1'b0;
      act_regs_data_2_13_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_136_cse ) begin
      act_regs_data_2_13_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_267_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_12_nl, and_dcpl_1246);
      act_regs_data_2_13_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_265_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_2_13_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_910_cse
          , act_regs_data_and_911_cse});
      act_regs_data_2_13_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_266_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_2_13_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_910_cse
          , act_regs_data_and_911_cse});
      act_regs_data_2_13_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_90_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_2_13_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_910_cse
          , act_regs_data_and_911_cse});
      act_regs_data_2_13_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_332_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_2_13_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_910_cse
          , act_regs_data_and_911_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_12_sva_8_31 <= 1'b0;
      act_regs_data_2_12_sva_8_30_26 <= 5'b00000;
      act_regs_data_2_12_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_2_12_sva_8_25 <= 1'b0;
      act_regs_data_2_12_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_140_cse ) begin
      act_regs_data_2_12_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_255_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_16_nl, and_dcpl_1246);
      act_regs_data_2_12_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_253_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_2_12_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_916_cse
          , act_regs_data_and_917_cse});
      act_regs_data_2_12_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_254_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_2_12_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_916_cse
          , act_regs_data_and_917_cse});
      act_regs_data_2_12_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_83_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_2_12_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_916_cse
          , act_regs_data_and_917_cse});
      act_regs_data_2_12_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_330_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_2_12_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_916_cse
          , act_regs_data_and_917_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_11_sva_8_31 <= 1'b0;
      act_regs_data_2_11_sva_8_30_26 <= 5'b00000;
      act_regs_data_2_11_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_2_11_sva_8_25 <= 1'b0;
      act_regs_data_2_11_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_144_cse ) begin
      act_regs_data_2_11_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_243_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_20_nl, and_dcpl_1246);
      act_regs_data_2_11_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_241_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_2_11_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_922_cse
          , act_regs_data_and_923_cse});
      act_regs_data_2_11_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_242_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_2_11_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_922_cse
          , act_regs_data_and_923_cse});
      act_regs_data_2_11_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_76_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_2_11_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_922_cse
          , act_regs_data_and_923_cse});
      act_regs_data_2_11_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_328_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_2_11_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_922_cse
          , act_regs_data_and_923_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_10_sva_8_31 <= 1'b0;
      act_regs_data_2_10_sva_8_30_26 <= 5'b00000;
      act_regs_data_2_10_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_2_10_sva_8_25 <= 1'b0;
      act_regs_data_2_10_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_148_cse ) begin
      act_regs_data_2_10_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_132_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_24_nl, and_dcpl_1246);
      act_regs_data_2_10_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_130_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_2_10_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_928_cse
          , act_regs_data_and_929_cse});
      act_regs_data_2_10_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_131_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_2_10_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_928_cse
          , act_regs_data_and_929_cse});
      act_regs_data_2_10_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_12_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_2_10_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_928_cse
          , act_regs_data_and_929_cse});
      act_regs_data_2_10_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_326_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_2_10_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_928_cse
          , act_regs_data_and_929_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_9_sva_8_31 <= 1'b0;
      act_regs_data_2_9_sva_8_30_26 <= 5'b00000;
      act_regs_data_2_9_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_2_9_sva_8_25 <= 1'b0;
      act_regs_data_2_9_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_152_cse ) begin
      act_regs_data_2_9_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_219_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_28_nl, and_dcpl_1246);
      act_regs_data_2_9_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_217_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_2_9_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_934_cse
          , act_regs_data_and_935_cse});
      act_regs_data_2_9_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_218_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_2_9_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_934_cse
          , act_regs_data_and_935_cse});
      act_regs_data_2_9_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_62_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_2_9_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_934_cse
          , act_regs_data_and_935_cse});
      act_regs_data_2_9_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_324_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_2_9_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_934_cse
          , act_regs_data_and_935_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_8_sva_8_31 <= 1'b0;
      act_regs_data_2_8_sva_8_30_26 <= 5'b00000;
      act_regs_data_2_8_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_2_8_sva_8_25 <= 1'b0;
      act_regs_data_2_8_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_156_cse ) begin
      act_regs_data_2_8_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_204_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_32_nl, and_dcpl_1246);
      act_regs_data_2_8_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_202_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_2_8_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_940_cse
          , act_regs_data_and_941_cse});
      act_regs_data_2_8_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_203_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_2_8_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_940_cse
          , act_regs_data_and_941_cse});
      act_regs_data_2_8_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_54_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_2_8_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_940_cse
          , act_regs_data_and_941_cse});
      act_regs_data_2_8_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_322_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_2_8_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_940_cse
          , act_regs_data_and_941_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_7_sva_8_31 <= 1'b0;
      act_regs_data_2_7_sva_8_30_26 <= 5'b00000;
      act_regs_data_2_7_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_2_7_sva_8_25 <= 1'b0;
      act_regs_data_2_7_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_160_cse ) begin
      act_regs_data_2_7_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_192_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_36_nl, and_dcpl_1246);
      act_regs_data_2_7_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_190_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_2_7_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_946_cse
          , act_regs_data_and_947_cse});
      act_regs_data_2_7_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_191_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_2_7_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_946_cse
          , act_regs_data_and_947_cse});
      act_regs_data_2_7_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_47_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_2_7_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_946_cse
          , act_regs_data_and_947_cse});
      act_regs_data_2_7_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_320_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_2_7_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_946_cse
          , act_regs_data_and_947_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_6_sva_8_31 <= 1'b0;
      act_regs_data_2_6_sva_8_30_26 <= 5'b00000;
      act_regs_data_2_6_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_2_6_sva_8_25 <= 1'b0;
      act_regs_data_2_6_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_164_cse ) begin
      act_regs_data_2_6_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_180_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_40_nl, and_dcpl_1246);
      act_regs_data_2_6_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_178_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_2_6_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_952_cse
          , act_regs_data_and_953_cse});
      act_regs_data_2_6_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_179_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_2_6_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_952_cse
          , act_regs_data_and_953_cse});
      act_regs_data_2_6_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_40_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_2_6_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_952_cse
          , act_regs_data_and_953_cse});
      act_regs_data_2_6_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_318_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_2_6_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_952_cse
          , act_regs_data_and_953_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_5_sva_8_31 <= 1'b0;
      act_regs_data_2_5_sva_8_30_26 <= 5'b00000;
      act_regs_data_2_5_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_2_5_sva_8_25 <= 1'b0;
      act_regs_data_2_5_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_168_cse ) begin
      act_regs_data_2_5_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_168_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_44_nl, and_dcpl_1246);
      act_regs_data_2_5_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_166_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_2_5_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_958_cse
          , act_regs_data_and_959_cse});
      act_regs_data_2_5_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_167_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_2_5_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_958_cse
          , act_regs_data_and_959_cse});
      act_regs_data_2_5_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_33_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_2_5_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_958_cse
          , act_regs_data_and_959_cse});
      act_regs_data_2_5_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_316_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_2_5_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_958_cse
          , act_regs_data_and_959_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_4_sva_8_31 <= 1'b0;
      act_regs_data_2_4_sva_8_30_26 <= 5'b00000;
      act_regs_data_2_4_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_2_4_sva_8_25 <= 1'b0;
      act_regs_data_2_4_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_172_cse ) begin
      act_regs_data_2_4_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_156_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_48_nl, and_dcpl_1246);
      act_regs_data_2_4_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_154_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_2_4_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_964_cse
          , act_regs_data_and_965_cse});
      act_regs_data_2_4_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_155_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_2_4_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_964_cse
          , act_regs_data_and_965_cse});
      act_regs_data_2_4_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_26_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_2_4_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_964_cse
          , act_regs_data_and_965_cse});
      act_regs_data_2_4_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_314_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_2_4_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_964_cse
          , act_regs_data_and_965_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_3_sva_8_31 <= 1'b0;
      act_regs_data_2_3_sva_8_30_26 <= 5'b00000;
      act_regs_data_2_3_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_2_3_sva_8_25 <= 1'b0;
      act_regs_data_2_3_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_176_cse ) begin
      act_regs_data_2_3_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_144_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_52_nl, and_dcpl_1246);
      act_regs_data_2_3_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_142_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_2_3_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_970_cse
          , act_regs_data_and_971_cse});
      act_regs_data_2_3_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_143_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_2_3_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_970_cse
          , act_regs_data_and_971_cse});
      act_regs_data_2_3_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_19_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_2_3_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_970_cse
          , act_regs_data_and_971_cse});
      act_regs_data_2_3_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_312_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_2_3_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_970_cse
          , act_regs_data_and_971_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_2_sva_8_31 <= 1'b0;
      act_regs_data_2_2_sva_8_30_26 <= 5'b00000;
      act_regs_data_2_2_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_2_2_sva_8_25 <= 1'b0;
      act_regs_data_2_2_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_180_cse ) begin
      act_regs_data_2_2_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_303_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_56_nl, and_dcpl_1246);
      act_regs_data_2_2_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_301_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_2_2_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_976_cse
          , act_regs_data_and_977_cse});
      act_regs_data_2_2_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_302_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_2_2_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_976_cse
          , act_regs_data_and_977_cse});
      act_regs_data_2_2_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_111_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_2_2_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_976_cse
          , act_regs_data_and_977_cse});
      act_regs_data_2_2_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_310_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_2_2_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_976_cse
          , act_regs_data_and_977_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_1_sva_8_31 <= 1'b0;
      act_regs_data_2_1_sva_8_30_26 <= 5'b00000;
      act_regs_data_2_1_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_2_1_sva_8_25 <= 1'b0;
      act_regs_data_2_1_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_184_cse ) begin
      act_regs_data_2_1_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_120_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_60_nl, and_dcpl_1246);
      act_regs_data_2_1_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_118_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_2_1_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_982_cse
          , act_regs_data_and_983_cse});
      act_regs_data_2_1_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_119_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_2_1_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_982_cse
          , act_regs_data_and_983_cse});
      act_regs_data_2_1_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_5_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_2_1_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_982_cse
          , act_regs_data_and_983_cse});
      act_regs_data_2_1_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_308_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_2_1_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_982_cse
          , act_regs_data_and_983_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_0_sva_8_31 <= 1'b0;
      act_regs_data_2_0_sva_8_30_26 <= 5'b00000;
      act_regs_data_2_0_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_2_0_sva_8_25 <= 1'b0;
      act_regs_data_2_0_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_188_cse ) begin
      act_regs_data_2_0_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_225_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_64_nl, and_dcpl_1246);
      act_regs_data_2_0_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_223_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_2_0_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_988_cse
          , act_regs_data_and_989_cse});
      act_regs_data_2_0_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_224_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_2_0_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_988_cse
          , act_regs_data_and_989_cse});
      act_regs_data_2_0_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_67_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_2_0_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_988_cse
          , act_regs_data_and_989_cse});
      act_regs_data_2_0_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_306_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_2_0_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_988_cse
          , act_regs_data_and_989_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_15_sva_8_31 <= 1'b0;
      act_regs_data_1_15_sva_8_30_26 <= 5'b00000;
      act_regs_data_1_15_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_1_15_sva_8_25 <= 1'b0;
      act_regs_data_1_15_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_192_cse ) begin
      act_regs_data_1_15_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_285_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_68_nl, and_dcpl_1246);
      act_regs_data_1_15_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_283_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_1_15_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_994_cse
          , act_regs_data_and_995_cse});
      act_regs_data_1_15_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_284_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_1_15_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_994_cse
          , act_regs_data_and_995_cse});
      act_regs_data_1_15_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_102_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_1_15_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_994_cse
          , act_regs_data_and_995_cse});
      act_regs_data_1_15_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_305_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_1_15_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_994_cse
          , act_regs_data_and_995_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_14_sva_8_31 <= 1'b0;
      act_regs_data_1_14_sva_8_30_26 <= 5'b00000;
      act_regs_data_1_14_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_1_14_sva_8_25 <= 1'b0;
      act_regs_data_1_14_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_196_cse ) begin
      act_regs_data_1_14_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_273_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_72_nl, and_dcpl_1246);
      act_regs_data_1_14_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_271_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_1_14_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_1000_cse
          , act_regs_data_and_1001_cse});
      act_regs_data_1_14_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_272_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_1_14_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_1000_cse
          , act_regs_data_and_1001_cse});
      act_regs_data_1_14_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_95_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_1_14_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_1000_cse
          , act_regs_data_and_1001_cse});
      act_regs_data_1_14_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_307_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_1_14_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_1000_cse
          , act_regs_data_and_1001_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_13_sva_8_31 <= 1'b0;
      act_regs_data_1_13_sva_8_30_26 <= 5'b00000;
      act_regs_data_1_13_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_1_13_sva_8_25 <= 1'b0;
      act_regs_data_1_13_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_200_cse ) begin
      act_regs_data_1_13_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_261_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_76_nl, and_dcpl_1246);
      act_regs_data_1_13_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_259_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_1_13_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_1006_cse
          , act_regs_data_and_1007_cse});
      act_regs_data_1_13_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_260_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_1_13_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_1006_cse
          , act_regs_data_and_1007_cse});
      act_regs_data_1_13_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_88_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_1_13_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_1006_cse
          , act_regs_data_and_1007_cse});
      act_regs_data_1_13_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_309_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_1_13_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_1006_cse
          , act_regs_data_and_1007_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_12_sva_8_31 <= 1'b0;
      act_regs_data_1_12_sva_8_30_26 <= 5'b00000;
      act_regs_data_1_12_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_1_12_sva_8_25 <= 1'b0;
      act_regs_data_1_12_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_204_cse ) begin
      act_regs_data_1_12_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_249_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_80_nl, and_dcpl_1246);
      act_regs_data_1_12_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_247_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_1_12_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_1012_cse
          , act_regs_data_and_1013_cse});
      act_regs_data_1_12_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_248_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_1_12_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_1012_cse
          , act_regs_data_and_1013_cse});
      act_regs_data_1_12_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_81_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_1_12_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_1012_cse
          , act_regs_data_and_1013_cse});
      act_regs_data_1_12_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_311_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_1_12_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_1012_cse
          , act_regs_data_and_1013_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_11_sva_8_31 <= 1'b0;
      act_regs_data_1_11_sva_8_30_26 <= 5'b00000;
      act_regs_data_1_11_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_1_11_sva_8_25 <= 1'b0;
      act_regs_data_1_11_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_208_cse ) begin
      act_regs_data_1_11_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_237_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_84_nl, and_dcpl_1246);
      act_regs_data_1_11_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_235_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_1_11_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_1018_cse
          , act_regs_data_and_1019_cse});
      act_regs_data_1_11_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_236_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_1_11_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_1018_cse
          , act_regs_data_and_1019_cse});
      act_regs_data_1_11_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_74_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_1_11_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_1018_cse
          , act_regs_data_and_1019_cse});
      act_regs_data_1_11_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_313_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_1_11_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_1018_cse
          , act_regs_data_and_1019_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_10_sva_8_31 <= 1'b0;
      act_regs_data_1_10_sva_8_30_26 <= 5'b00000;
      act_regs_data_1_10_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_1_10_sva_8_25 <= 1'b0;
      act_regs_data_1_10_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_212_cse ) begin
      act_regs_data_1_10_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_126_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_88_nl, and_dcpl_1246);
      act_regs_data_1_10_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_124_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_1_10_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_1024_cse
          , act_regs_data_and_1025_cse});
      act_regs_data_1_10_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_125_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_1_10_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_1024_cse
          , act_regs_data_and_1025_cse});
      act_regs_data_1_10_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_10_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_1_10_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_1024_cse
          , act_regs_data_and_1025_cse});
      act_regs_data_1_10_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_315_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_1_10_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_1024_cse
          , act_regs_data_and_1025_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_9_sva_8_31 <= 1'b0;
      act_regs_data_1_9_sva_8_30_26 <= 5'b00000;
      act_regs_data_1_9_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_1_9_sva_8_25 <= 1'b0;
      act_regs_data_1_9_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_216_cse ) begin
      act_regs_data_1_9_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_213_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_92_nl, and_dcpl_1246);
      act_regs_data_1_9_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_211_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_1_9_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_1030_cse
          , act_regs_data_and_1031_cse});
      act_regs_data_1_9_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_212_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_1_9_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_1030_cse
          , act_regs_data_and_1031_cse});
      act_regs_data_1_9_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_60_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_1_9_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_1030_cse
          , act_regs_data_and_1031_cse});
      act_regs_data_1_9_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_317_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_1_9_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_1030_cse
          , act_regs_data_and_1031_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_8_sva_8_31 <= 1'b0;
      act_regs_data_1_8_sva_8_30_26 <= 5'b00000;
      act_regs_data_1_8_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_1_8_sva_8_25 <= 1'b0;
      act_regs_data_1_8_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_220_cse ) begin
      act_regs_data_1_8_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_198_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_96_nl, and_dcpl_1246);
      act_regs_data_1_8_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_196_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_1_8_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_1036_cse
          , act_regs_data_and_1037_cse});
      act_regs_data_1_8_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_197_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_1_8_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_1036_cse
          , act_regs_data_and_1037_cse});
      act_regs_data_1_8_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_52_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_1_8_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_1036_cse
          , act_regs_data_and_1037_cse});
      act_regs_data_1_8_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_319_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_1_8_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_1036_cse
          , act_regs_data_and_1037_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_7_sva_8_31 <= 1'b0;
      act_regs_data_1_7_sva_8_30_26 <= 5'b00000;
      act_regs_data_1_7_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_1_7_sva_8_25 <= 1'b0;
      act_regs_data_1_7_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_224_cse ) begin
      act_regs_data_1_7_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_186_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_100_nl, and_dcpl_1246);
      act_regs_data_1_7_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_184_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_1_7_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_1042_cse
          , act_regs_data_and_1043_cse});
      act_regs_data_1_7_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_185_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_1_7_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_1042_cse
          , act_regs_data_and_1043_cse});
      act_regs_data_1_7_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_45_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_1_7_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_1042_cse
          , act_regs_data_and_1043_cse});
      act_regs_data_1_7_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_321_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_1_7_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_1042_cse
          , act_regs_data_and_1043_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_6_sva_8_31 <= 1'b0;
      act_regs_data_1_6_sva_8_30_26 <= 5'b00000;
      act_regs_data_1_6_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_1_6_sva_8_25 <= 1'b0;
      act_regs_data_1_6_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_228_cse ) begin
      act_regs_data_1_6_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_174_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_104_nl, and_dcpl_1246);
      act_regs_data_1_6_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_172_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_1_6_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_1048_cse
          , act_regs_data_and_1049_cse});
      act_regs_data_1_6_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_173_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_1_6_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_1048_cse
          , act_regs_data_and_1049_cse});
      act_regs_data_1_6_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_38_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_1_6_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_1048_cse
          , act_regs_data_and_1049_cse});
      act_regs_data_1_6_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_323_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_1_6_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_1048_cse
          , act_regs_data_and_1049_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_5_sva_8_31 <= 1'b0;
      act_regs_data_1_5_sva_8_30_26 <= 5'b00000;
      act_regs_data_1_5_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_1_5_sva_8_25 <= 1'b0;
      act_regs_data_1_5_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_232_cse ) begin
      act_regs_data_1_5_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_162_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_108_nl, and_dcpl_1246);
      act_regs_data_1_5_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_160_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_1_5_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_1054_cse
          , act_regs_data_and_1055_cse});
      act_regs_data_1_5_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_161_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_1_5_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_1054_cse
          , act_regs_data_and_1055_cse});
      act_regs_data_1_5_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_31_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_1_5_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_1054_cse
          , act_regs_data_and_1055_cse});
      act_regs_data_1_5_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_325_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_1_5_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_1054_cse
          , act_regs_data_and_1055_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_4_sva_8_31 <= 1'b0;
      act_regs_data_1_4_sva_8_30_26 <= 5'b00000;
      act_regs_data_1_4_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_1_4_sva_8_25 <= 1'b0;
      act_regs_data_1_4_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_236_cse ) begin
      act_regs_data_1_4_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_150_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_112_nl, and_dcpl_1246);
      act_regs_data_1_4_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_148_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_1_4_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_1060_cse
          , act_regs_data_and_1061_cse});
      act_regs_data_1_4_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_149_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_1_4_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_1060_cse
          , act_regs_data_and_1061_cse});
      act_regs_data_1_4_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_24_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_1_4_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_1060_cse
          , act_regs_data_and_1061_cse});
      act_regs_data_1_4_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_327_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_1_4_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_1060_cse
          , act_regs_data_and_1061_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_3_sva_8_31 <= 1'b0;
      act_regs_data_1_3_sva_8_30_26 <= 5'b00000;
      act_regs_data_1_3_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_1_3_sva_8_25 <= 1'b0;
      act_regs_data_1_3_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_240_cse ) begin
      act_regs_data_1_3_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_138_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_116_nl, and_dcpl_1246);
      act_regs_data_1_3_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_136_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_1_3_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_1066_cse
          , act_regs_data_and_1067_cse});
      act_regs_data_1_3_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_137_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_1_3_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_1066_cse
          , act_regs_data_and_1067_cse});
      act_regs_data_1_3_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_17_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_1_3_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_1066_cse
          , act_regs_data_and_1067_cse});
      act_regs_data_1_3_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_329_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_1_3_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_1066_cse
          , act_regs_data_and_1067_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_2_sva_8_31 <= 1'b0;
      act_regs_data_1_2_sva_8_30_26 <= 5'b00000;
      act_regs_data_1_2_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_1_2_sva_8_25 <= 1'b0;
      act_regs_data_1_2_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_244_cse ) begin
      act_regs_data_1_2_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_297_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_120_nl, and_dcpl_1246);
      act_regs_data_1_2_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_295_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_1_2_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_1072_cse
          , act_regs_data_and_1073_cse});
      act_regs_data_1_2_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_296_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_1_2_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_1072_cse
          , act_regs_data_and_1073_cse});
      act_regs_data_1_2_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_109_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_1_2_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_1072_cse
          , act_regs_data_and_1073_cse});
      act_regs_data_1_2_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_331_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_1_2_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_1072_cse
          , act_regs_data_and_1073_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_1_sva_8_31 <= 1'b0;
      act_regs_data_1_1_sva_8_30_26 <= 5'b00000;
      act_regs_data_1_1_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_1_1_sva_8_25 <= 1'b0;
      act_regs_data_1_1_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_248_cse ) begin
      act_regs_data_1_1_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_114_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_124_nl, and_dcpl_1246);
      act_regs_data_1_1_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_112_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_1_1_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_1078_cse
          , act_regs_data_and_1079_cse});
      act_regs_data_1_1_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_113_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_1_1_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_1078_cse
          , act_regs_data_and_1079_cse});
      act_regs_data_1_1_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_3_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_1_1_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_1078_cse
          , act_regs_data_and_1079_cse});
      act_regs_data_1_1_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_333_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_1_1_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_1078_cse
          , act_regs_data_and_1079_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_0_sva_8_31 <= 1'b0;
      act_regs_data_1_0_sva_8_30_26 <= 5'b00000;
      act_regs_data_1_0_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_1_0_sva_8_25 <= 1'b0;
      act_regs_data_1_0_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_252_cse ) begin
      act_regs_data_1_0_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_222_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_128_nl, and_dcpl_1246);
      act_regs_data_1_0_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_220_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_1_0_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_1084_cse
          , act_regs_data_and_1085_cse});
      act_regs_data_1_0_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_221_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_1_0_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_1084_cse
          , act_regs_data_and_1085_cse});
      act_regs_data_1_0_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_66_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_1_0_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_1084_cse
          , act_regs_data_and_1085_cse});
      act_regs_data_1_0_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_335_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_1_0_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_1084_cse
          , act_regs_data_and_1085_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_15_sva_8_31 <= 1'b0;
      act_regs_data_0_15_sva_8_30_26 <= 5'b00000;
      act_regs_data_0_15_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_0_15_sva_8_25 <= 1'b0;
      act_regs_data_0_15_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_256_cse ) begin
      act_regs_data_0_15_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_282_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_132_nl, and_dcpl_1246);
      act_regs_data_0_15_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_280_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_0_15_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_1090_cse
          , act_regs_data_and_1091_cse});
      act_regs_data_0_15_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_281_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_0_15_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_1090_cse
          , act_regs_data_and_1091_cse});
      act_regs_data_0_15_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_101_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_0_15_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_1090_cse
          , act_regs_data_and_1091_cse});
      act_regs_data_0_15_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_337_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_0_15_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_1090_cse
          , act_regs_data_and_1091_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_14_sva_8_31 <= 1'b0;
      act_regs_data_0_14_sva_8_30_26 <= 5'b00000;
      act_regs_data_0_14_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_0_14_sva_8_25 <= 1'b0;
      act_regs_data_0_14_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_260_cse ) begin
      act_regs_data_0_14_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_270_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_136_nl, and_dcpl_1246);
      act_regs_data_0_14_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_268_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_0_14_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_1096_cse
          , act_regs_data_and_1097_cse});
      act_regs_data_0_14_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_269_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_0_14_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_1096_cse
          , act_regs_data_and_1097_cse});
      act_regs_data_0_14_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_94_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_0_14_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_1096_cse
          , act_regs_data_and_1097_cse});
      act_regs_data_0_14_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_339_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_0_14_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_1096_cse
          , act_regs_data_and_1097_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_13_sva_8_31 <= 1'b0;
      act_regs_data_0_13_sva_8_30_26 <= 5'b00000;
      act_regs_data_0_13_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_0_13_sva_8_25 <= 1'b0;
      act_regs_data_0_13_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_264_cse ) begin
      act_regs_data_0_13_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_258_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_140_nl, and_dcpl_1246);
      act_regs_data_0_13_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_256_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_0_13_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_1102_cse
          , act_regs_data_and_1103_cse});
      act_regs_data_0_13_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_257_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_0_13_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_1102_cse
          , act_regs_data_and_1103_cse});
      act_regs_data_0_13_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_87_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_0_13_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_1102_cse
          , act_regs_data_and_1103_cse});
      act_regs_data_0_13_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_340_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_0_13_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_1102_cse
          , act_regs_data_and_1103_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_12_sva_8_31 <= 1'b0;
      act_regs_data_0_12_sva_8_30_26 <= 5'b00000;
      act_regs_data_0_12_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_0_12_sva_8_25 <= 1'b0;
      act_regs_data_0_12_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_268_cse ) begin
      act_regs_data_0_12_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_246_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_144_nl, and_dcpl_1246);
      act_regs_data_0_12_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_244_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_0_12_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_1108_cse
          , act_regs_data_and_1109_cse});
      act_regs_data_0_12_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_245_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_0_12_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_1108_cse
          , act_regs_data_and_1109_cse});
      act_regs_data_0_12_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_80_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_0_12_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_1108_cse
          , act_regs_data_and_1109_cse});
      act_regs_data_0_12_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_341_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_0_12_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_1108_cse
          , act_regs_data_and_1109_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_11_sva_8_31 <= 1'b0;
      act_regs_data_0_11_sva_8_30_26 <= 5'b00000;
      act_regs_data_0_11_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_0_11_sva_8_25 <= 1'b0;
      act_regs_data_0_11_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_272_cse ) begin
      act_regs_data_0_11_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_234_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_148_nl, and_dcpl_1246);
      act_regs_data_0_11_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_232_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_0_11_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_1114_cse
          , act_regs_data_and_1115_cse});
      act_regs_data_0_11_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_233_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_0_11_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_1114_cse
          , act_regs_data_and_1115_cse});
      act_regs_data_0_11_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_73_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_0_11_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_1114_cse
          , act_regs_data_and_1115_cse});
      act_regs_data_0_11_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_342_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_0_11_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_1114_cse
          , act_regs_data_and_1115_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_10_sva_8_31 <= 1'b0;
      act_regs_data_0_10_sva_8_30_26 <= 5'b00000;
      act_regs_data_0_10_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_0_10_sva_8_25 <= 1'b0;
      act_regs_data_0_10_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_276_cse ) begin
      act_regs_data_0_10_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_129_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_152_nl, and_dcpl_1246);
      act_regs_data_0_10_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_127_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_0_10_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_1120_cse
          , act_regs_data_and_1121_cse});
      act_regs_data_0_10_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_128_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_0_10_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_1120_cse
          , act_regs_data_and_1121_cse});
      act_regs_data_0_10_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_11_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_0_10_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_1120_cse
          , act_regs_data_and_1121_cse});
      act_regs_data_0_10_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_343_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_0_10_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_1120_cse
          , act_regs_data_and_1121_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_9_sva_8_31 <= 1'b0;
      act_regs_data_0_9_sva_8_30_26 <= 5'b00000;
      act_regs_data_0_9_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_0_9_sva_8_25 <= 1'b0;
      act_regs_data_0_9_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_280_cse ) begin
      act_regs_data_0_9_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_210_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_156_nl, and_dcpl_1246);
      act_regs_data_0_9_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_208_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_0_9_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_1126_cse
          , act_regs_data_and_1127_cse});
      act_regs_data_0_9_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_209_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_0_9_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_1126_cse
          , act_regs_data_and_1127_cse});
      act_regs_data_0_9_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_59_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_0_9_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_1126_cse
          , act_regs_data_and_1127_cse});
      act_regs_data_0_9_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_344_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_0_9_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_1126_cse
          , act_regs_data_and_1127_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_8_sva_8_31 <= 1'b0;
      act_regs_data_0_8_sva_8_30_26 <= 5'b00000;
      act_regs_data_0_8_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_0_8_sva_8_25 <= 1'b0;
      act_regs_data_0_8_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_284_cse ) begin
      act_regs_data_0_8_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_201_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_160_nl, and_dcpl_1246);
      act_regs_data_0_8_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_199_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_0_8_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_1132_cse
          , act_regs_data_and_1133_cse});
      act_regs_data_0_8_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_200_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_0_8_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_1132_cse
          , act_regs_data_and_1133_cse});
      act_regs_data_0_8_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_53_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_0_8_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_1132_cse
          , act_regs_data_and_1133_cse});
      act_regs_data_0_8_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_345_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_0_8_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_1132_cse
          , act_regs_data_and_1133_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_7_sva_8_31 <= 1'b0;
      act_regs_data_0_7_sva_8_30_26 <= 5'b00000;
      act_regs_data_0_7_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_0_7_sva_8_25 <= 1'b0;
      act_regs_data_0_7_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_288_cse ) begin
      act_regs_data_0_7_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_189_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_164_nl, and_dcpl_1246);
      act_regs_data_0_7_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_187_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_0_7_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_1138_cse
          , act_regs_data_and_1139_cse});
      act_regs_data_0_7_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_188_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_0_7_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_1138_cse
          , act_regs_data_and_1139_cse});
      act_regs_data_0_7_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_46_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_0_7_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_1138_cse
          , act_regs_data_and_1139_cse});
      act_regs_data_0_7_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_346_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_0_7_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_1138_cse
          , act_regs_data_and_1139_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_6_sva_8_31 <= 1'b0;
      act_regs_data_0_6_sva_8_30_26 <= 5'b00000;
      act_regs_data_0_6_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_0_6_sva_8_25 <= 1'b0;
      act_regs_data_0_6_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_292_cse ) begin
      act_regs_data_0_6_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_177_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_168_nl, and_dcpl_1246);
      act_regs_data_0_6_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_175_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_0_6_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_1144_cse
          , act_regs_data_and_1145_cse});
      act_regs_data_0_6_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_176_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_0_6_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_1144_cse
          , act_regs_data_and_1145_cse});
      act_regs_data_0_6_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_39_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_0_6_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_1144_cse
          , act_regs_data_and_1145_cse});
      act_regs_data_0_6_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_347_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_0_6_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_1144_cse
          , act_regs_data_and_1145_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_5_sva_8_31 <= 1'b0;
      act_regs_data_0_5_sva_8_30_26 <= 5'b00000;
      act_regs_data_0_5_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_0_5_sva_8_25 <= 1'b0;
      act_regs_data_0_5_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_296_cse ) begin
      act_regs_data_0_5_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_165_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_172_nl, and_dcpl_1246);
      act_regs_data_0_5_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_163_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_0_5_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_1150_cse
          , act_regs_data_and_1151_cse});
      act_regs_data_0_5_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_164_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_0_5_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_1150_cse
          , act_regs_data_and_1151_cse});
      act_regs_data_0_5_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_32_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_0_5_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_1150_cse
          , act_regs_data_and_1151_cse});
      act_regs_data_0_5_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_348_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_0_5_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_1150_cse
          , act_regs_data_and_1151_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_4_sva_8_31 <= 1'b0;
      act_regs_data_0_4_sva_8_30_26 <= 5'b00000;
      act_regs_data_0_4_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_0_4_sva_8_25 <= 1'b0;
      act_regs_data_0_4_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_300_cse ) begin
      act_regs_data_0_4_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_153_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_176_nl, and_dcpl_1246);
      act_regs_data_0_4_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_151_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_0_4_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_1156_cse
          , act_regs_data_and_1157_cse});
      act_regs_data_0_4_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_152_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_0_4_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_1156_cse
          , act_regs_data_and_1157_cse});
      act_regs_data_0_4_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_25_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_0_4_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_1156_cse
          , act_regs_data_and_1157_cse});
      act_regs_data_0_4_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_349_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_0_4_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_1156_cse
          , act_regs_data_and_1157_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_3_sva_8_31 <= 1'b0;
      act_regs_data_0_3_sva_8_30_26 <= 5'b00000;
      act_regs_data_0_3_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_0_3_sva_8_25 <= 1'b0;
      act_regs_data_0_3_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_304_cse ) begin
      act_regs_data_0_3_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_141_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_180_nl, and_dcpl_1246);
      act_regs_data_0_3_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_139_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_0_3_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_1162_cse
          , act_regs_data_and_1163_cse});
      act_regs_data_0_3_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_140_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_0_3_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_1162_cse
          , act_regs_data_and_1163_cse});
      act_regs_data_0_3_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_18_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_0_3_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_1162_cse
          , act_regs_data_and_1163_cse});
      act_regs_data_0_3_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_350_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_0_3_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_1162_cse
          , act_regs_data_and_1163_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_2_sva_8_31 <= 1'b0;
      act_regs_data_0_2_sva_8_30_26 <= 5'b00000;
      act_regs_data_0_2_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_0_2_sva_8_25 <= 1'b0;
      act_regs_data_0_2_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_308_cse ) begin
      act_regs_data_0_2_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_294_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_184_nl, and_dcpl_1246);
      act_regs_data_0_2_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_292_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_0_2_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_1168_cse
          , act_regs_data_and_1169_cse});
      act_regs_data_0_2_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_293_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_0_2_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_1168_cse
          , act_regs_data_and_1169_cse});
      act_regs_data_0_2_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_108_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_0_2_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_1168_cse
          , act_regs_data_and_1169_cse});
      act_regs_data_0_2_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_351_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_0_2_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_1168_cse
          , act_regs_data_and_1169_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_1_sva_8_31 <= 1'b0;
      act_regs_data_0_1_sva_8_30_26 <= 5'b00000;
      act_regs_data_0_1_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_0_1_sva_8_25 <= 1'b0;
      act_regs_data_0_1_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_312_cse ) begin
      act_regs_data_0_1_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_117_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_188_nl, and_dcpl_1246);
      act_regs_data_0_1_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_115_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_0_1_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_1174_cse
          , act_regs_data_and_1175_cse});
      act_regs_data_0_1_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_116_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_0_1_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_1174_cse
          , act_regs_data_and_1175_cse});
      act_regs_data_0_1_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_4_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_0_1_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_1174_cse
          , act_regs_data_and_1175_cse});
      act_regs_data_0_1_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_352_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_0_1_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_1174_cse
          , act_regs_data_and_1175_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_0_sva_8_31 <= 1'b0;
      act_regs_data_0_0_sva_8_30_26 <= 5'b00000;
      act_regs_data_0_0_sva_8_21_0 <= 22'b0000000000000000000000;
      act_regs_data_0_0_sva_8_25 <= 1'b0;
      act_regs_data_0_0_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_316_cse ) begin
      act_regs_data_0_0_sva_8_31 <= MUX_s_1_2_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_228_nl,
          ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_192_nl, and_dcpl_1246);
      act_regs_data_0_0_sva_8_30_26 <= MUX1HOT_v_5_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_226_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          act_regs_data_0_0_sva_dfm_2_30_26, {(~ and_dcpl_1246) , act_regs_data_and_1180_cse
          , act_regs_data_and_1181_cse});
      act_regs_data_0_0_sva_8_21_0 <= MUX1HOT_v_22_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_227_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          act_regs_data_0_0_sva_dfm_2_21_0, {(~ and_dcpl_1246) , act_regs_data_and_1180_cse
          , act_regs_data_and_1181_cse});
      act_regs_data_0_0_sva_8_25 <= MUX1HOT_s_1_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_68_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_0_0_sva_dfm_2_25_22_rsp_0, {(~ and_dcpl_1246) , act_regs_data_and_1180_cse
          , act_regs_data_and_1181_cse});
      act_regs_data_0_0_sva_8_24_22 <= MUX1HOT_v_3_3_2(nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_353_nl,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_0_0_sva_dfm_2_25_22_rsp_1, {(~ and_dcpl_1246) , act_regs_data_and_1180_cse
          , act_regs_data_and_1181_cse});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_CheckStart_start_reg_sva <= 1'b0;
    end
    else if ( ActUnitRun_wen & mux_451_nl ) begin
      ActUnit_CheckStart_start_reg_sva <= MUX1HOT_s_1_3_2(ActUnit_RunInst_switch_lp_and_48_tmp_1,
          start_PopNB_mioi_data_rsc_z_mxwt, while_and_64_nl, {and_dcpl_331 , and_dcpl_1244
          , and_dcpl_1104});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      Silu_for_y_8_lpi_1_dfm_4_31 <= 1'b0;
      Silu_for_y_8_lpi_1_dfm_4_21_0 <= 22'b0000000000000000000000;
      Silu_for_y_7_lpi_1_dfm_4_31 <= 1'b0;
      Silu_for_y_7_lpi_1_dfm_4_21_0 <= 22'b0000000000000000000000;
      Silu_for_y_6_lpi_1_dfm_4_31 <= 1'b0;
      Silu_for_y_6_lpi_1_dfm_4_21_0 <= 22'b0000000000000000000000;
      Silu_for_y_5_lpi_1_dfm_4_31 <= 1'b0;
      Silu_for_y_5_lpi_1_dfm_4_21_0 <= 22'b0000000000000000000000;
      Silu_for_y_4_lpi_1_dfm_4_31 <= 1'b0;
      Silu_for_y_4_lpi_1_dfm_4_21_0 <= 22'b0000000000000000000000;
      Silu_for_y_3_lpi_1_dfm_4_31 <= 1'b0;
      Silu_for_y_3_lpi_1_dfm_4_21_0 <= 22'b0000000000000000000000;
      Silu_for_y_2_lpi_1_dfm_4_31 <= 1'b0;
      Silu_for_y_2_lpi_1_dfm_4_21_0 <= 22'b0000000000000000000000;
      Silu_for_y_1_lpi_1_dfm_4_31 <= 1'b0;
      Silu_for_y_1_lpi_1_dfm_4_21_0 <= 22'b0000000000000000000000;
      Silu_for_y_8_lpi_1_dfm_4_25 <= 1'b0;
      Silu_for_y_8_lpi_1_dfm_4_24_22 <= 3'b000;
      Silu_for_y_7_lpi_1_dfm_4_25 <= 1'b0;
      Silu_for_y_7_lpi_1_dfm_4_24_22 <= 3'b000;
      Silu_for_y_6_lpi_1_dfm_4_25 <= 1'b0;
      Silu_for_y_6_lpi_1_dfm_4_24_22 <= 3'b000;
      Silu_for_y_5_lpi_1_dfm_4_25 <= 1'b0;
      Silu_for_y_5_lpi_1_dfm_4_24_22 <= 3'b000;
      Silu_for_y_4_lpi_1_dfm_4_25 <= 1'b0;
      Silu_for_y_4_lpi_1_dfm_4_24_22 <= 3'b000;
      Silu_for_y_3_lpi_1_dfm_4_25 <= 1'b0;
      Silu_for_y_3_lpi_1_dfm_4_24_22 <= 3'b000;
      Silu_for_y_2_lpi_1_dfm_4_25 <= 1'b0;
      Silu_for_y_2_lpi_1_dfm_4_24_22 <= 3'b000;
      Silu_for_y_1_lpi_1_dfm_4_25 <= 1'b0;
      Silu_for_y_1_lpi_1_dfm_4_24_22 <= 3'b000;
    end
    else if ( Silu_for_y_and_2_cse ) begin
      Silu_for_y_8_lpi_1_dfm_4_31 <= Silu_for_else_mux_32_nl & (~(Silu_for_else_and_39_ssc_1
          | Silu_for_else_else_else_and_14_ssc_1 | Silu_for_else_else_else_and_15_ssc_1))
          & Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
      Silu_for_y_8_lpi_1_dfm_4_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000, ({Silu_for_else_Silu_for_else_mux1h_39_nl
          , Silu_for_else_Silu_for_else_mux1h_48_nl}), Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
      Silu_for_y_7_lpi_1_dfm_4_31 <= Silu_for_else_mux_33_nl & (~(Silu_for_else_and_38_ssc_1
          | Silu_for_else_else_else_and_12_ssc_1 | Silu_for_else_else_else_and_13_ssc_1))
          & Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
      Silu_for_y_7_lpi_1_dfm_4_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000, ({Silu_for_else_Silu_for_else_mux1h_38_nl
          , Silu_for_else_Silu_for_else_mux1h_50_nl}), Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
      Silu_for_y_6_lpi_1_dfm_4_31 <= Silu_for_else_mux_34_nl & (~(Silu_for_else_and_37_ssc_1
          | Silu_for_else_else_else_and_10_ssc_1 | Silu_for_else_else_else_and_11_ssc_1))
          & Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
      Silu_for_y_6_lpi_1_dfm_4_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000, ({Silu_for_else_Silu_for_else_mux1h_37_nl
          , Silu_for_else_Silu_for_else_mux1h_52_nl}), Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
      Silu_for_y_5_lpi_1_dfm_4_31 <= Silu_for_else_mux_35_nl & (~(Silu_for_else_and_36_ssc_1
          | Silu_for_else_else_else_and_8_ssc_1 | Silu_for_else_else_else_and_9_ssc_1))
          & Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
      Silu_for_y_5_lpi_1_dfm_4_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000, ({Silu_for_else_Silu_for_else_mux1h_36_nl
          , Silu_for_else_Silu_for_else_mux1h_54_nl}), Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
      Silu_for_y_4_lpi_1_dfm_4_31 <= Silu_for_else_mux_36_nl & (~(Silu_for_else_and_35_ssc_1
          | Silu_for_else_else_else_and_6_ssc_1 | Silu_for_else_else_else_and_7_ssc_1))
          & Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
      Silu_for_y_4_lpi_1_dfm_4_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000, ({Silu_for_else_Silu_for_else_mux1h_35_nl
          , Silu_for_else_Silu_for_else_mux1h_56_nl}), Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
      Silu_for_y_3_lpi_1_dfm_4_31 <= Silu_for_else_mux_37_nl & (~(Silu_for_else_and_34_ssc_1
          | Silu_for_else_else_else_and_4_ssc_1 | Silu_for_else_else_else_and_5_ssc_1))
          & Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
      Silu_for_y_3_lpi_1_dfm_4_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000, ({Silu_for_else_Silu_for_else_mux1h_34_nl
          , Silu_for_else_Silu_for_else_mux1h_58_nl}), Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
      Silu_for_y_2_lpi_1_dfm_4_31 <= Silu_for_else_mux_38_nl & (~(Silu_for_else_and_33_ssc_1
          | Silu_for_else_else_else_and_2_ssc_1 | Silu_for_else_else_else_and_3_ssc_1))
          & Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
      Silu_for_y_2_lpi_1_dfm_4_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000, ({Silu_for_else_Silu_for_else_mux1h_33_nl
          , Silu_for_else_Silu_for_else_mux1h_60_nl}), Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
      Silu_for_y_1_lpi_1_dfm_4_31 <= Silu_for_else_mux_39_nl & (~(Silu_for_else_and_32_ssc_1
          | Silu_for_else_else_else_and_ssc_1 | Silu_for_else_else_else_and_1_ssc_1))
          & Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
      Silu_for_y_1_lpi_1_dfm_4_21_0 <= MUX_v_22_2_2(22'b0000000000000000000000, ({Silu_for_else_Silu_for_else_mux1h_32_nl
          , Silu_for_else_Silu_for_else_mux1h_62_nl}), Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
      Silu_for_y_8_lpi_1_dfm_4_25 <= Silu_for_else_Silu_for_else_mux1h_23_nl & (~
          Silu_for_else_and_39_ssc_1) & Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
      Silu_for_y_8_lpi_1_dfm_4_24_22 <= MUX_v_3_2_2(3'b000, Silu_for_else_Silu_for_else_mux1h_49_nl,
          Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
      Silu_for_y_7_lpi_1_dfm_4_25 <= Silu_for_else_Silu_for_else_mux1h_22_nl & (~
          Silu_for_else_and_38_ssc_1) & Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
      Silu_for_y_7_lpi_1_dfm_4_24_22 <= MUX_v_3_2_2(3'b000, Silu_for_else_Silu_for_else_mux1h_51_nl,
          Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
      Silu_for_y_6_lpi_1_dfm_4_25 <= Silu_for_else_Silu_for_else_mux1h_21_nl & (~
          Silu_for_else_and_37_ssc_1) & Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
      Silu_for_y_6_lpi_1_dfm_4_24_22 <= MUX_v_3_2_2(3'b000, Silu_for_else_Silu_for_else_mux1h_53_nl,
          Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
      Silu_for_y_5_lpi_1_dfm_4_25 <= Silu_for_else_Silu_for_else_mux1h_20_nl & (~
          Silu_for_else_and_36_ssc_1) & Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
      Silu_for_y_5_lpi_1_dfm_4_24_22 <= MUX_v_3_2_2(3'b000, Silu_for_else_Silu_for_else_mux1h_55_nl,
          Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
      Silu_for_y_4_lpi_1_dfm_4_25 <= Silu_for_else_Silu_for_else_mux1h_19_nl & (~
          Silu_for_else_and_35_ssc_1) & Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
      Silu_for_y_4_lpi_1_dfm_4_24_22 <= MUX_v_3_2_2(3'b000, Silu_for_else_Silu_for_else_mux1h_57_nl,
          Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
      Silu_for_y_3_lpi_1_dfm_4_25 <= Silu_for_else_Silu_for_else_mux1h_18_nl & (~
          Silu_for_else_and_34_ssc_1) & Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
      Silu_for_y_3_lpi_1_dfm_4_24_22 <= MUX_v_3_2_2(3'b000, Silu_for_else_Silu_for_else_mux1h_59_nl,
          Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
      Silu_for_y_2_lpi_1_dfm_4_25 <= Silu_for_else_Silu_for_else_mux1h_17_nl & (~
          Silu_for_else_and_33_ssc_1) & Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
      Silu_for_y_2_lpi_1_dfm_4_24_22 <= MUX_v_3_2_2(3'b000, Silu_for_else_Silu_for_else_mux1h_61_nl,
          Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
      Silu_for_y_1_lpi_1_dfm_4_25 <= Silu_for_else_Silu_for_else_mux1h_16_nl & (~
          Silu_for_else_and_32_ssc_1) & Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs;
      Silu_for_y_1_lpi_1_dfm_4_24_22 <= MUX_v_3_2_2(3'b000, Silu_for_else_Silu_for_else_mux1h_63_nl,
          Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_1_30_26 <= 5'b00000;
    end
    else if ( and_1909_tmp ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_1_30_26 <= MUX_v_5_2_2(5'b00000,
          ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_70_nl, not_8877_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_1_30_26 <= 5'b00000;
    end
    else if ( and_1915_tmp ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_1_30_26 <= MUX_v_5_2_2(5'b00000,
          ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_75_nl, not_8878_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_1_30_26 <= 5'b00000;
    end
    else if ( and_1921_tmp ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_1_30_26 <= MUX_v_5_2_2(5'b00000,
          ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_80_nl, not_8879_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_1_30_26 <= 5'b00000;
    end
    else if ( and_1927_tmp ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_1_30_26 <= MUX_v_5_2_2(5'b00000,
          ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_85_nl, not_8880_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_1_30_26 <= 5'b00000;
    end
    else if ( and_1933_tmp ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_1_30_26 <= MUX_v_5_2_2(5'b00000,
          ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_90_nl, not_8881_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_1_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_817 | and_dcpl_1090)) | and_dcpl_1236)
        ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_1_31 <= MUX_s_1_2_2(ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_31_3,
          nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_123_nl, and_dcpl_1236);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_1_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_826 | and_dcpl_1090)) | and_dcpl_1244
        | and_dcpl_1236) ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_1_31 <= ActUnit_PushOutput_if_output_port_reg_data_data_mux_nl
          & (~ and_dcpl_1244);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_1_sva_1_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_828 | and_dcpl_1090)) | and_dcpl_1244
        | and_dcpl_1236) ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_1_sva_1_31 <= ActUnit_PushOutput_if_output_port_reg_data_data_mux_1_nl
          & (~ and_dcpl_1244);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_1_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_829 | and_dcpl_1090)) | and_dcpl_1244
        | and_dcpl_1236) ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_1_31 <= ActUnit_PushOutput_if_output_port_reg_data_data_mux_2_nl
          & (~ and_dcpl_1244);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_1_31 <= 1'b0;
      ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_1_30_26 <= 5'b00000;
    end
    else if ( ActUnit_PushOutput_if_output_port_reg_data_data_and_22_cse ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_1_31 <= ActUnit_PushOutput_if_output_port_reg_data_data_mux_3_nl
          & (~ and_dcpl_1244);
      ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_1_30_26 <= MUX_v_5_2_2(5'b00000,
          ActUnit_PushOutput_if_output_port_reg_data_data_mux_4_nl, not_8882_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_1_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_831 | and_dcpl_1090)) | and_dcpl_1244
        | and_dcpl_1236) ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_1_31 <= ActUnit_PushOutput_if_output_port_reg_data_data_mux_5_nl
          & (~ and_dcpl_1244);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_1_31 <= 1'b0;
      ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_1_30_26 <= 5'b00000;
    end
    else if ( ActUnit_PushOutput_if_output_port_reg_data_data_and_25_cse ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_1_31 <= ActUnit_PushOutput_if_output_port_reg_data_data_mux_6_nl
          & (~ and_dcpl_1244);
      ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_1_30_26 <= MUX_v_5_2_2(5'b00000,
          ActUnit_PushOutput_if_output_port_reg_data_data_mux_7_nl, not_8883_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_1_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_835 | and_dcpl_1090)) | and_dcpl_1244
        | and_dcpl_1236) ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_1_31 <= ActUnit_PushOutput_if_output_port_reg_data_data_mux_8_nl
          & (~ and_dcpl_1244);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_1_31 <= 1'b0;
      ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_1_30_26 <= 5'b00000;
    end
    else if ( ActUnit_PushOutput_if_output_port_reg_data_data_and_28_cse ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_1_31 <= ActUnit_PushOutput_if_output_port_reg_data_data_mux_9_nl
          & (~ and_dcpl_1244);
      ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_1_30_26 <= MUX_v_5_2_2(5'b00000,
          ActUnit_PushOutput_if_output_port_reg_data_data_mux_10_nl, not_8884_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_1_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_838 | and_dcpl_1090)) | and_dcpl_1244
        | and_dcpl_1236) ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_1_31 <= ActUnit_PushOutput_if_output_port_reg_data_data_mux_11_nl
          & (~ and_dcpl_1244);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_1_31 <= 1'b0;
      ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_1_30_26 <= 5'b00000;
    end
    else if ( ActUnit_PushOutput_if_output_port_reg_data_data_and_31_cse ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_1_31 <= ActUnit_PushOutput_if_output_port_reg_data_data_mux_12_nl
          & (~ and_dcpl_1244);
      ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_1_30_26 <= MUX_v_5_2_2(5'b00000,
          ActUnit_PushOutput_if_output_port_reg_data_data_mux_13_nl, not_8885_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_1_31 <= 1'b0;
      ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_1_30_26 <= 5'b00000;
      ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_1_25 <= 1'b0;
      ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_1_24_22 <= 3'b000;
    end
    else if ( ActUnit_PushOutput_if_output_port_reg_data_data_and_33_cse ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_1_31 <= ActUnit_PushOutput_if_output_port_reg_data_data_mux_14_nl
          & (~ and_dcpl_1244);
      ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_1_30_26 <= MUX_v_5_2_2(5'b00000,
          ActUnit_PushOutput_if_output_port_reg_data_data_mux_15_nl, not_8886_nl);
      ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_1_25 <= ActUnit_PushOutput_if_for_i_mux_nl
          & (~ or_dcpl);
      ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_1_24_22 <= MUX_v_3_2_2(3'b000,
          ActUnit_PushOutput_if_for_i_mux_1_nl, not_8896_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_1_31 <= 1'b0;
      ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_1_30_26 <= 5'b00000;
    end
    else if ( ActUnit_PushOutput_if_output_port_reg_data_data_and_36_cse ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_1_31 <= ActUnit_PushOutput_if_output_port_reg_data_data_mux_16_nl
          & (~ and_dcpl_1244);
      ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_1_30_26 <= MUX_v_5_2_2(5'b00000,
          ActUnit_PushOutput_if_output_port_reg_data_data_mux_17_nl, not_8888_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_1_31 <= 1'b0;
      ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_1_30_26 <= 5'b00000;
    end
    else if ( ActUnit_PushOutput_if_output_port_reg_data_data_and_38_cse ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_1_31 <= ActUnit_PushOutput_if_output_port_reg_data_data_mux_18_nl
          & (~ and_dcpl_1244);
      ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_1_30_26 <= MUX_v_5_2_2(5'b00000,
          ActUnit_PushOutput_if_output_port_reg_data_data_mux_19_nl, not_8889_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_1_31 <= 1'b0;
      ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_1_30_26 <= 5'b00000;
    end
    else if ( ActUnit_PushOutput_if_output_port_reg_data_data_and_40_cse ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_1_31 <= ActUnit_PushOutput_if_output_port_reg_data_data_mux_20_nl
          & (~ and_dcpl_1244);
      ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_1_30_26 <= MUX_v_5_2_2(5'b00000,
          ActUnit_PushOutput_if_output_port_reg_data_data_mux_21_nl, not_8890_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_0_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_936 | or_dcpl_866 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_0_0_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_213_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_1_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_936 | or_dcpl_864 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_0_1_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_214_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_2_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_936 | or_dcpl_861 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_0_2_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_215_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_3_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_936 | or_dcpl_859 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_0_3_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_216_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_4_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_936 | or_dcpl_856 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_0_4_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_217_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_5_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_936 | or_dcpl_854 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_0_5_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_218_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_6_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_936 | or_dcpl_851 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_0_6_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_219_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_7_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_936 | or_dcpl_847 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_0_7_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_220_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_8_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_946 | or_dcpl_866 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_0_8_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_221_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_9_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_946 | or_dcpl_864 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_0_9_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_222_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_10_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_946 | or_dcpl_861 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_0_10_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_223_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_11_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_946 | or_dcpl_859 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_0_11_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_224_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_12_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_946 | or_dcpl_856 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_0_12_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_225_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_13_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_946 | or_dcpl_854 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_0_13_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_226_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_14_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_946 | or_dcpl_851 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_0_14_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_227_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_15_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_946 | or_dcpl_847 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_0_15_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_228_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_0_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_956 | or_dcpl_866 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_1_0_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_229_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_1_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_956 | or_dcpl_864 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_1_1_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_230_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_2_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_956 | or_dcpl_861 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_1_2_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_231_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_3_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_956 | or_dcpl_859 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_1_3_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_232_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_4_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_956 | or_dcpl_856 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_1_4_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_233_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_5_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_956 | or_dcpl_854 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_1_5_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_234_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_6_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_956 | or_dcpl_851 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_1_6_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_235_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_7_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_956 | or_dcpl_847 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_1_7_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_236_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_8_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_965 | or_dcpl_866 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_1_8_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_237_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_9_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_965 | or_dcpl_864 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_1_9_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_238_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_10_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_965 | or_dcpl_861 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_1_10_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_239_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_11_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_965 | or_dcpl_859 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_1_11_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_240_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_12_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_965 | or_dcpl_856 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_1_12_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_241_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_13_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_965 | or_dcpl_854 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_1_13_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_242_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_14_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_965 | or_dcpl_851 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_1_14_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_243_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_15_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_965 | or_dcpl_847 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_1_15_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_244_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_0_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_975 | or_dcpl_866 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_2_0_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_245_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_1_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_975 | or_dcpl_864 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_2_1_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_246_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_2_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_975 | or_dcpl_861 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_2_2_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_247_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_3_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_975 | or_dcpl_859 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_2_3_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_248_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_4_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_975 | or_dcpl_856 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_2_4_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_249_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_5_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_975 | or_dcpl_854 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_2_5_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_250_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_6_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_975 | or_dcpl_851 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_2_6_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_251_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_7_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_975 | or_dcpl_847 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_2_7_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_252_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_8_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_985 | or_dcpl_866 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_2_8_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_253_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_9_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_985 | or_dcpl_864 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_2_9_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_254_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_10_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_985 | or_dcpl_861 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_2_10_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_255_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_11_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_985 | or_dcpl_859 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_2_11_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_256_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_12_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_985 | or_dcpl_856 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_2_12_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_257_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_13_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_985 | or_dcpl_854 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_2_13_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_258_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_14_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_985 | or_dcpl_851 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_2_14_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_259_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_15_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_985 | or_dcpl_847 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_2_15_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_260_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_0_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_994 | or_dcpl_866 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_3_0_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_261_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_1_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_994 | or_dcpl_864 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_3_1_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_262_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_2_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_994 | or_dcpl_861 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_3_2_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_263_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_3_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_994 | or_dcpl_859 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_3_3_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_264_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_4_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_994 | or_dcpl_856 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_3_4_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_265_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_5_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_994 | or_dcpl_854 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_3_5_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_266_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_6_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_994 | or_dcpl_851 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_3_6_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_267_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_7_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_994 | or_dcpl_847 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_3_7_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_268_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_8_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_1003 | or_dcpl_866 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_3_8_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_269_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_9_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_1003 | or_dcpl_864 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_3_9_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_270_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_10_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_1003 | or_dcpl_861 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_3_10_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_271_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_11_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_1003 | or_dcpl_859 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_3_11_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_272_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_12_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_1003 | or_dcpl_856 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_3_12_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_273_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_13_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_1003 | or_dcpl_854 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_3_13_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_274_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_14_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_1003 | or_dcpl_851 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_3_14_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_275_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_15_sva_dfm_2_31 <= 1'b0;
    end
    else if ( ActUnitRun_wen & ((~(or_dcpl_1003 | or_dcpl_847 | not_tmp_640)) | and_dcpl_1244)
        ) begin
      act_regs_data_3_15_sva_dfm_2_31 <= MUX_s_1_2_2(while_and_276_nl, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
          and_dcpl_1246);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_0_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_0_0_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_0_0_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_1935_cse ) begin
      act_regs_data_0_0_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(reg_act_regs_data_0_0_ftd_3,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[21:0]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_1_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_1_lpi_1_dfm_21_0,
          Silu_for_y_1_lpi_1_dfm_4_21_0, Gelu_for_y_1_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
      act_regs_data_0_0_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(reg_act_regs_data_0_0_ftd_2_3,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[25]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_1_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_1_lpi_1_dfm_25,
          Silu_for_y_1_lpi_1_dfm_4_25, Gelu_for_y_1_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
      act_regs_data_0_0_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(reg_act_regs_data_0_0_ftd_2_2_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[24:22]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_1_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_1_lpi_1_dfm_24_22,
          Silu_for_y_1_lpi_1_dfm_4_24_22, Gelu_for_y_1_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_1_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_0_1_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_0_1_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_1937_cse ) begin
      act_regs_data_0_1_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(reg_act_regs_data_0_1_ftd_3,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[53:32]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_2_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_2_lpi_1_dfm_21_0,
          Silu_for_y_2_lpi_1_dfm_4_21_0, Gelu_for_y_2_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
      act_regs_data_0_1_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(reg_act_regs_data_0_1_ftd_2_3,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[57]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_2_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_2_lpi_1_dfm_25,
          Silu_for_y_2_lpi_1_dfm_4_25, Gelu_for_y_2_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
      act_regs_data_0_1_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(reg_act_regs_data_0_1_ftd_2_2_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[56:54]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_2_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_2_lpi_1_dfm_24_22,
          Silu_for_y_2_lpi_1_dfm_4_24_22, Gelu_for_y_2_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_2_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_0_2_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_0_2_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_1939_cse ) begin
      act_regs_data_0_2_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_0_2_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[85:64]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_3_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_3_lpi_1_dfm_21_0,
          Silu_for_y_3_lpi_1_dfm_4_21_0, Gelu_for_y_3_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
      act_regs_data_0_2_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_0_2_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[89]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_3_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_3_lpi_1_dfm_25,
          Silu_for_y_3_lpi_1_dfm_4_25, Gelu_for_y_3_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
      act_regs_data_0_2_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_0_2_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[88:86]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_3_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_3_lpi_1_dfm_24_22,
          Silu_for_y_3_lpi_1_dfm_4_24_22, Gelu_for_y_3_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_3_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_0_3_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_0_3_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_1941_cse ) begin
      act_regs_data_0_3_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_0_3_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[117:96]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_4_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_4_lpi_1_dfm_21_0,
          Silu_for_y_4_lpi_1_dfm_4_21_0, Gelu_for_y_4_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
      act_regs_data_0_3_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_0_3_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[121]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_4_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_4_lpi_1_dfm_25,
          Silu_for_y_4_lpi_1_dfm_4_25, Gelu_for_y_4_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
      act_regs_data_0_3_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_0_3_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[120:118]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_4_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_4_lpi_1_dfm_24_22,
          Silu_for_y_4_lpi_1_dfm_4_24_22, Gelu_for_y_4_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_4_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_0_4_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_0_4_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_1943_cse ) begin
      act_regs_data_0_4_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_0_4_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[149:128]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_5_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_5_lpi_1_dfm_21_0,
          Silu_for_y_5_lpi_1_dfm_4_21_0, Gelu_for_y_5_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
      act_regs_data_0_4_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_0_4_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[153]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_5_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_5_lpi_1_dfm_25,
          Silu_for_y_5_lpi_1_dfm_4_25, Gelu_for_y_5_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
      act_regs_data_0_4_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_0_4_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[152:150]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_5_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_5_lpi_1_dfm_24_22,
          Silu_for_y_5_lpi_1_dfm_4_24_22, Gelu_for_y_5_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_5_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_0_5_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_0_5_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_1945_cse ) begin
      act_regs_data_0_5_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_0_5_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[181:160]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_6_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_6_lpi_1_dfm_21_0,
          Silu_for_y_6_lpi_1_dfm_4_21_0, Gelu_for_y_6_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
      act_regs_data_0_5_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_0_5_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[185]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_6_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_6_lpi_1_dfm_25,
          Silu_for_y_6_lpi_1_dfm_4_25, Gelu_for_y_6_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
      act_regs_data_0_5_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_0_5_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[184:182]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_6_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_6_lpi_1_dfm_24_22,
          Silu_for_y_6_lpi_1_dfm_4_24_22, Gelu_for_y_6_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_6_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_0_6_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_0_6_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_1947_cse ) begin
      act_regs_data_0_6_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_0_6_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[213:192]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_7_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_7_lpi_1_dfm_21_0,
          Silu_for_y_7_lpi_1_dfm_4_21_0, Gelu_for_y_7_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
      act_regs_data_0_6_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_0_6_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[217]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_7_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_7_lpi_1_dfm_25,
          Silu_for_y_7_lpi_1_dfm_4_25, Gelu_for_y_7_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
      act_regs_data_0_6_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_0_6_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[216:214]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_7_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_7_lpi_1_dfm_24_22,
          Silu_for_y_7_lpi_1_dfm_4_24_22, Gelu_for_y_7_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_7_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_0_7_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_0_7_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_1949_cse ) begin
      act_regs_data_0_7_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_0_7_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[245:224]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_8_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_8_lpi_1_dfm_21_0,
          Silu_for_y_8_lpi_1_dfm_4_21_0, Gelu_for_y_8_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
      act_regs_data_0_7_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_0_7_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[249]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_8_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_8_lpi_1_dfm_25,
          Silu_for_y_8_lpi_1_dfm_4_25, Gelu_for_y_8_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
      act_regs_data_0_7_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_0_7_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[248:246]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_8_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_8_lpi_1_dfm_24_22,
          Silu_for_y_8_lpi_1_dfm_4_24_22, Gelu_for_y_8_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_8_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_0_8_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_0_8_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_1951_cse ) begin
      act_regs_data_0_8_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_0_8_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[277:256]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_9_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_9_lpi_1_dfm_21_0,
          Silu_for_y_9_lpi_1_dfm_4_21_0_1, Gelu_for_y_9_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
      act_regs_data_0_8_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_0_8_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[281]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_9_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_9_lpi_1_dfm_25,
          Silu_for_y_9_lpi_1_dfm_4_25, Gelu_for_y_9_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
      act_regs_data_0_8_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_0_8_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[280:278]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_9_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_9_lpi_1_dfm_24_22,
          Silu_for_y_9_lpi_1_dfm_4_24_22, Gelu_for_y_9_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_9_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_0_9_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_0_9_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_1953_cse ) begin
      act_regs_data_0_9_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_0_9_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[309:288]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_10_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_10_lpi_1_dfm_21_0,
          Silu_for_y_10_lpi_1_dfm_4_21_0_1, Gelu_for_y_10_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
      act_regs_data_0_9_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_0_9_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[313]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_10_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_10_lpi_1_dfm_25,
          Silu_for_y_10_lpi_1_dfm_4_25, Gelu_for_y_10_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
      act_regs_data_0_9_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_0_9_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[312:310]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_10_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_10_lpi_1_dfm_24_22,
          Silu_for_y_10_lpi_1_dfm_4_24_22, Gelu_for_y_10_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_10_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_0_10_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_0_10_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_1955_cse ) begin
      act_regs_data_0_10_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(reg_act_regs_data_0_10_ftd_3,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[341:320]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_11_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_11_lpi_1_dfm_21_0,
          Silu_for_y_11_lpi_1_dfm_4_21_0_1, Gelu_for_y_11_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
      act_regs_data_0_10_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(reg_act_regs_data_0_10_ftd_2_3,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[345]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_11_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_11_lpi_1_dfm_25,
          Silu_for_y_11_lpi_1_dfm_4_25, Gelu_for_y_11_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
      act_regs_data_0_10_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(reg_act_regs_data_0_10_ftd_2_2_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[344:342]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_11_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_11_lpi_1_dfm_24_22,
          Silu_for_y_11_lpi_1_dfm_4_24_22, Gelu_for_y_11_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_11_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_0_11_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_0_11_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_1957_cse ) begin
      act_regs_data_0_11_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(reg_act_regs_data_0_11_ftd_3,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[373:352]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_12_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_12_lpi_1_dfm_21_0,
          Silu_for_y_12_lpi_1_dfm_4_21_0_1, Gelu_for_y_12_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
      act_regs_data_0_11_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(reg_act_regs_data_0_11_ftd_2_3,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[377]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_12_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_12_lpi_1_dfm_25,
          Silu_for_y_12_lpi_1_dfm_4_25, Gelu_for_y_12_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
      act_regs_data_0_11_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(reg_act_regs_data_0_11_ftd_2_2_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[376:374]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_12_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_12_lpi_1_dfm_24_22,
          Silu_for_y_12_lpi_1_dfm_4_24_22, Gelu_for_y_12_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_12_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_0_12_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_0_12_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_1959_cse ) begin
      act_regs_data_0_12_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(reg_act_regs_data_0_12_ftd_3,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[405:384]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_13_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_13_lpi_1_dfm_21_0,
          Silu_for_y_13_lpi_1_dfm_4_21_0_1, Gelu_for_y_13_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
      act_regs_data_0_12_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(reg_act_regs_data_0_12_ftd_2_3,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[409]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_13_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_13_lpi_1_dfm_25,
          Silu_for_y_13_lpi_1_dfm_4_25, Gelu_for_y_13_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
      act_regs_data_0_12_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(reg_act_regs_data_0_12_ftd_2_2_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[408:406]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_13_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_13_lpi_1_dfm_24_22,
          Silu_for_y_13_lpi_1_dfm_4_24_22, Gelu_for_y_13_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_13_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_0_13_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_0_13_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_1961_cse ) begin
      act_regs_data_0_13_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(reg_act_regs_data_0_13_ftd_3,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[437:416]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_14_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_14_lpi_1_dfm_21_0,
          Silu_for_y_14_lpi_1_dfm_4_21_0_1, Gelu_for_y_14_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
      act_regs_data_0_13_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(reg_act_regs_data_0_13_ftd_2_3,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[441]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_14_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_14_lpi_1_dfm_25,
          Silu_for_y_14_lpi_1_dfm_4_25, Gelu_for_y_14_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
      act_regs_data_0_13_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(reg_act_regs_data_0_13_ftd_2_2_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[440:438]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_14_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_14_lpi_1_dfm_24_22,
          Silu_for_y_14_lpi_1_dfm_4_24_22, Gelu_for_y_14_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_14_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_0_14_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_0_14_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_1963_cse ) begin
      act_regs_data_0_14_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_0_14_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[469:448]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_15_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_15_lpi_1_dfm_21_0,
          Silu_for_y_15_lpi_1_dfm_4_21_0_1, Gelu_for_y_15_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
      act_regs_data_0_14_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_0_14_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[473]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_15_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_15_lpi_1_dfm_25,
          Silu_for_y_15_lpi_1_dfm_4_25, Gelu_for_y_15_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
      act_regs_data_0_14_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_0_14_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[472:470]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_15_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_15_lpi_1_dfm_24_22,
          Silu_for_y_15_lpi_1_dfm_4_24_22, Gelu_for_y_15_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_15_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_0_15_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_0_15_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_1965_cse ) begin
      act_regs_data_0_15_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_0_15_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[501:480]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_lpi_1_dfm_21_0, Silu_for_y_lpi_1_dfm_4_21_0_1,
          Gelu_for_y_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
      act_regs_data_0_15_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_0_15_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[505]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_lpi_1_dfm_25, Silu_for_y_lpi_1_dfm_4_25,
          Gelu_for_y_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
      act_regs_data_0_15_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_0_15_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[504:502]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_lpi_1_dfm_24_22,
          Silu_for_y_lpi_1_dfm_4_24_22, Gelu_for_y_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_0_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_1_0_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_1_0_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_1967_cse ) begin
      act_regs_data_1_0_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_1_0_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[21:0]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_1_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_1_lpi_1_dfm_21_0,
          Silu_for_y_1_lpi_1_dfm_4_21_0, Gelu_for_y_1_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
      act_regs_data_1_0_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_1_0_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[25]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_1_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_1_lpi_1_dfm_25,
          Silu_for_y_1_lpi_1_dfm_4_25, Gelu_for_y_1_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
      act_regs_data_1_0_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_1_0_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[24:22]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_1_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_1_lpi_1_dfm_24_22,
          Silu_for_y_1_lpi_1_dfm_4_24_22, Gelu_for_y_1_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_1_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_1_1_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_1_1_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_1969_cse ) begin
      act_regs_data_1_1_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_1_1_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[53:32]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_2_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_2_lpi_1_dfm_21_0,
          Silu_for_y_2_lpi_1_dfm_4_21_0, Gelu_for_y_2_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
      act_regs_data_1_1_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_1_1_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[57]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_2_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_2_lpi_1_dfm_25,
          Silu_for_y_2_lpi_1_dfm_4_25, Gelu_for_y_2_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
      act_regs_data_1_1_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_1_1_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[56:54]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_2_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_2_lpi_1_dfm_24_22,
          Silu_for_y_2_lpi_1_dfm_4_24_22, Gelu_for_y_2_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_2_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_1_2_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_1_2_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_1971_cse ) begin
      act_regs_data_1_2_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_1_2_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[85:64]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_3_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_3_lpi_1_dfm_21_0,
          Silu_for_y_3_lpi_1_dfm_4_21_0, Gelu_for_y_3_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
      act_regs_data_1_2_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_1_2_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[89]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_3_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_3_lpi_1_dfm_25,
          Silu_for_y_3_lpi_1_dfm_4_25, Gelu_for_y_3_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
      act_regs_data_1_2_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_1_2_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[88:86]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_3_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_3_lpi_1_dfm_24_22,
          Silu_for_y_3_lpi_1_dfm_4_24_22, Gelu_for_y_3_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_3_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_1_3_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_1_3_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_1973_cse ) begin
      act_regs_data_1_3_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_1_3_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[117:96]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_4_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_4_lpi_1_dfm_21_0,
          Silu_for_y_4_lpi_1_dfm_4_21_0, Gelu_for_y_4_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
      act_regs_data_1_3_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_1_3_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[121]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_4_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_4_lpi_1_dfm_25,
          Silu_for_y_4_lpi_1_dfm_4_25, Gelu_for_y_4_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
      act_regs_data_1_3_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_1_3_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[120:118]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_4_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_4_lpi_1_dfm_24_22,
          Silu_for_y_4_lpi_1_dfm_4_24_22, Gelu_for_y_4_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_4_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_1_4_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_1_4_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_1975_cse ) begin
      act_regs_data_1_4_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_1_4_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[149:128]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_5_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_5_lpi_1_dfm_21_0,
          Silu_for_y_5_lpi_1_dfm_4_21_0, Gelu_for_y_5_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
      act_regs_data_1_4_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_1_4_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[153]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_5_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_5_lpi_1_dfm_25,
          Silu_for_y_5_lpi_1_dfm_4_25, Gelu_for_y_5_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
      act_regs_data_1_4_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_1_4_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[152:150]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_5_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_5_lpi_1_dfm_24_22,
          Silu_for_y_5_lpi_1_dfm_4_24_22, Gelu_for_y_5_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_5_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_1_5_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_1_5_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_1977_cse ) begin
      act_regs_data_1_5_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_1_5_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[181:160]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_6_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_6_lpi_1_dfm_21_0,
          Silu_for_y_6_lpi_1_dfm_4_21_0, Gelu_for_y_6_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
      act_regs_data_1_5_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_1_5_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[185]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_6_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_6_lpi_1_dfm_25,
          Silu_for_y_6_lpi_1_dfm_4_25, Gelu_for_y_6_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
      act_regs_data_1_5_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_1_5_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[184:182]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_6_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_6_lpi_1_dfm_24_22,
          Silu_for_y_6_lpi_1_dfm_4_24_22, Gelu_for_y_6_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_6_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_1_6_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_1_6_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_1979_cse ) begin
      act_regs_data_1_6_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_1_6_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[213:192]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_7_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_7_lpi_1_dfm_21_0,
          Silu_for_y_7_lpi_1_dfm_4_21_0, Gelu_for_y_7_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
      act_regs_data_1_6_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_1_6_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[217]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_7_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_7_lpi_1_dfm_25,
          Silu_for_y_7_lpi_1_dfm_4_25, Gelu_for_y_7_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
      act_regs_data_1_6_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_1_6_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[216:214]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_7_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_7_lpi_1_dfm_24_22,
          Silu_for_y_7_lpi_1_dfm_4_24_22, Gelu_for_y_7_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_7_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_1_7_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_1_7_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_1981_cse ) begin
      act_regs_data_1_7_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_1_7_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[245:224]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_8_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_8_lpi_1_dfm_21_0,
          Silu_for_y_8_lpi_1_dfm_4_21_0, Gelu_for_y_8_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
      act_regs_data_1_7_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_1_7_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[249]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_8_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_8_lpi_1_dfm_25,
          Silu_for_y_8_lpi_1_dfm_4_25, Gelu_for_y_8_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
      act_regs_data_1_7_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_1_7_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[248:246]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_8_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_8_lpi_1_dfm_24_22,
          Silu_for_y_8_lpi_1_dfm_4_24_22, Gelu_for_y_8_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_8_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_1_8_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_1_8_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_1983_cse ) begin
      act_regs_data_1_8_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_1_8_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[277:256]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_9_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_9_lpi_1_dfm_21_0,
          Silu_for_y_9_lpi_1_dfm_4_21_0_1, Gelu_for_y_9_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
      act_regs_data_1_8_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_1_8_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[281]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_9_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_9_lpi_1_dfm_25,
          Silu_for_y_9_lpi_1_dfm_4_25, Gelu_for_y_9_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
      act_regs_data_1_8_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_1_8_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[280:278]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_9_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_9_lpi_1_dfm_24_22,
          Silu_for_y_9_lpi_1_dfm_4_24_22, Gelu_for_y_9_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_9_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_1_9_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_1_9_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_1985_cse ) begin
      act_regs_data_1_9_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_1_9_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[309:288]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_10_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_10_lpi_1_dfm_21_0,
          Silu_for_y_10_lpi_1_dfm_4_21_0_1, Gelu_for_y_10_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
      act_regs_data_1_9_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_1_9_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[313]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_10_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_10_lpi_1_dfm_25,
          Silu_for_y_10_lpi_1_dfm_4_25, Gelu_for_y_10_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
      act_regs_data_1_9_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_1_9_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[312:310]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_10_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_10_lpi_1_dfm_24_22,
          Silu_for_y_10_lpi_1_dfm_4_24_22, Gelu_for_y_10_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_10_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_1_10_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_1_10_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_1987_cse ) begin
      act_regs_data_1_10_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_1_10_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[341:320]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_11_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_11_lpi_1_dfm_21_0,
          Silu_for_y_11_lpi_1_dfm_4_21_0_1, Gelu_for_y_11_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
      act_regs_data_1_10_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_1_10_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[345]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_11_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_11_lpi_1_dfm_25,
          Silu_for_y_11_lpi_1_dfm_4_25, Gelu_for_y_11_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
      act_regs_data_1_10_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_1_10_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[344:342]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_11_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_11_lpi_1_dfm_24_22,
          Silu_for_y_11_lpi_1_dfm_4_24_22, Gelu_for_y_11_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_11_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_1_11_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_1_11_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_1989_cse ) begin
      act_regs_data_1_11_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_1_11_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[373:352]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_12_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_12_lpi_1_dfm_21_0,
          Silu_for_y_12_lpi_1_dfm_4_21_0_1, Gelu_for_y_12_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
      act_regs_data_1_11_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_1_11_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[377]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_12_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_12_lpi_1_dfm_25,
          Silu_for_y_12_lpi_1_dfm_4_25, Gelu_for_y_12_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
      act_regs_data_1_11_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_1_11_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[376:374]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_12_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_12_lpi_1_dfm_24_22,
          Silu_for_y_12_lpi_1_dfm_4_24_22, Gelu_for_y_12_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_12_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_1_12_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_1_12_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_1991_cse ) begin
      act_regs_data_1_12_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_1_12_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[405:384]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_13_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_13_lpi_1_dfm_21_0,
          Silu_for_y_13_lpi_1_dfm_4_21_0_1, Gelu_for_y_13_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
      act_regs_data_1_12_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_1_12_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[409]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_13_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_13_lpi_1_dfm_25,
          Silu_for_y_13_lpi_1_dfm_4_25, Gelu_for_y_13_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
      act_regs_data_1_12_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_1_12_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[408:406]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_13_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_13_lpi_1_dfm_24_22,
          Silu_for_y_13_lpi_1_dfm_4_24_22, Gelu_for_y_13_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_13_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_1_13_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_1_13_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_1993_cse ) begin
      act_regs_data_1_13_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_1_13_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[437:416]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_14_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_14_lpi_1_dfm_21_0,
          Silu_for_y_14_lpi_1_dfm_4_21_0_1, Gelu_for_y_14_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
      act_regs_data_1_13_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_1_13_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[441]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_14_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_14_lpi_1_dfm_25,
          Silu_for_y_14_lpi_1_dfm_4_25, Gelu_for_y_14_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
      act_regs_data_1_13_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_1_13_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[440:438]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_14_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_14_lpi_1_dfm_24_22,
          Silu_for_y_14_lpi_1_dfm_4_24_22, Gelu_for_y_14_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_14_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_1_14_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_1_14_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_1995_cse ) begin
      act_regs_data_1_14_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_1_14_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[469:448]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_15_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_15_lpi_1_dfm_21_0,
          Silu_for_y_15_lpi_1_dfm_4_21_0_1, Gelu_for_y_15_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
      act_regs_data_1_14_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_1_14_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[473]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_15_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_15_lpi_1_dfm_25,
          Silu_for_y_15_lpi_1_dfm_4_25, Gelu_for_y_15_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
      act_regs_data_1_14_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_1_14_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[472:470]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_15_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_15_lpi_1_dfm_24_22,
          Silu_for_y_15_lpi_1_dfm_4_24_22, Gelu_for_y_15_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_15_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_1_15_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_1_15_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_1997_cse ) begin
      act_regs_data_1_15_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_1_15_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[501:480]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_lpi_1_dfm_21_0, Silu_for_y_lpi_1_dfm_4_21_0_1,
          Gelu_for_y_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
      act_regs_data_1_15_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_1_15_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[505]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_lpi_1_dfm_25, Silu_for_y_lpi_1_dfm_4_25,
          Gelu_for_y_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
      act_regs_data_1_15_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_1_15_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[504:502]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_lpi_1_dfm_24_22,
          Silu_for_y_lpi_1_dfm_4_24_22, Gelu_for_y_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_0_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_2_0_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_2_0_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_1999_cse ) begin
      act_regs_data_2_0_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_2_0_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[21:0]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_1_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_1_lpi_1_dfm_21_0,
          Silu_for_y_1_lpi_1_dfm_4_21_0, Gelu_for_y_1_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
      act_regs_data_2_0_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_2_0_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[25]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_1_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_1_lpi_1_dfm_25,
          Silu_for_y_1_lpi_1_dfm_4_25, Gelu_for_y_1_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
      act_regs_data_2_0_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_2_0_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[24:22]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_1_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_1_lpi_1_dfm_24_22,
          Silu_for_y_1_lpi_1_dfm_4_24_22, Gelu_for_y_1_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_1_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_2_1_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_2_1_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_2001_cse ) begin
      act_regs_data_2_1_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_2_1_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[53:32]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_2_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_2_lpi_1_dfm_21_0,
          Silu_for_y_2_lpi_1_dfm_4_21_0, Gelu_for_y_2_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
      act_regs_data_2_1_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_2_1_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[57]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_2_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_2_lpi_1_dfm_25,
          Silu_for_y_2_lpi_1_dfm_4_25, Gelu_for_y_2_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
      act_regs_data_2_1_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_2_1_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[56:54]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_2_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_2_lpi_1_dfm_24_22,
          Silu_for_y_2_lpi_1_dfm_4_24_22, Gelu_for_y_2_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_2_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_2_2_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_2_2_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_2003_cse ) begin
      act_regs_data_2_2_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_2_2_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[85:64]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_3_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_3_lpi_1_dfm_21_0,
          Silu_for_y_3_lpi_1_dfm_4_21_0, Gelu_for_y_3_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
      act_regs_data_2_2_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_2_2_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[89]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_3_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_3_lpi_1_dfm_25,
          Silu_for_y_3_lpi_1_dfm_4_25, Gelu_for_y_3_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
      act_regs_data_2_2_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_2_2_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[88:86]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_3_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_3_lpi_1_dfm_24_22,
          Silu_for_y_3_lpi_1_dfm_4_24_22, Gelu_for_y_3_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_3_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_2_3_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_2_3_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_2005_cse ) begin
      act_regs_data_2_3_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_2_3_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[117:96]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_4_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_4_lpi_1_dfm_21_0,
          Silu_for_y_4_lpi_1_dfm_4_21_0, Gelu_for_y_4_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
      act_regs_data_2_3_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_2_3_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[121]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_4_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_4_lpi_1_dfm_25,
          Silu_for_y_4_lpi_1_dfm_4_25, Gelu_for_y_4_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
      act_regs_data_2_3_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_2_3_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[120:118]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_4_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_4_lpi_1_dfm_24_22,
          Silu_for_y_4_lpi_1_dfm_4_24_22, Gelu_for_y_4_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_4_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_2_4_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_2_4_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_2007_cse ) begin
      act_regs_data_2_4_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_2_4_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[149:128]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_5_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_5_lpi_1_dfm_21_0,
          Silu_for_y_5_lpi_1_dfm_4_21_0, Gelu_for_y_5_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
      act_regs_data_2_4_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_2_4_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[153]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_5_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_5_lpi_1_dfm_25,
          Silu_for_y_5_lpi_1_dfm_4_25, Gelu_for_y_5_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
      act_regs_data_2_4_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_2_4_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[152:150]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_5_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_5_lpi_1_dfm_24_22,
          Silu_for_y_5_lpi_1_dfm_4_24_22, Gelu_for_y_5_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_5_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_2_5_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_2_5_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_2009_cse ) begin
      act_regs_data_2_5_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_2_5_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[181:160]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_6_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_6_lpi_1_dfm_21_0,
          Silu_for_y_6_lpi_1_dfm_4_21_0, Gelu_for_y_6_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
      act_regs_data_2_5_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_2_5_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[185]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_6_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_6_lpi_1_dfm_25,
          Silu_for_y_6_lpi_1_dfm_4_25, Gelu_for_y_6_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
      act_regs_data_2_5_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_2_5_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[184:182]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_6_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_6_lpi_1_dfm_24_22,
          Silu_for_y_6_lpi_1_dfm_4_24_22, Gelu_for_y_6_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_6_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_2_6_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_2_6_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_2011_cse ) begin
      act_regs_data_2_6_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_2_6_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[213:192]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_7_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_7_lpi_1_dfm_21_0,
          Silu_for_y_7_lpi_1_dfm_4_21_0, Gelu_for_y_7_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
      act_regs_data_2_6_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_2_6_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[217]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_7_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_7_lpi_1_dfm_25,
          Silu_for_y_7_lpi_1_dfm_4_25, Gelu_for_y_7_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
      act_regs_data_2_6_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_2_6_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[216:214]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_7_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_7_lpi_1_dfm_24_22,
          Silu_for_y_7_lpi_1_dfm_4_24_22, Gelu_for_y_7_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_7_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_2_7_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_2_7_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_2013_cse ) begin
      act_regs_data_2_7_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_2_7_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[245:224]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_8_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_8_lpi_1_dfm_21_0,
          Silu_for_y_8_lpi_1_dfm_4_21_0, Gelu_for_y_8_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
      act_regs_data_2_7_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_2_7_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[249]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_8_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_8_lpi_1_dfm_25,
          Silu_for_y_8_lpi_1_dfm_4_25, Gelu_for_y_8_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
      act_regs_data_2_7_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_2_7_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[248:246]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_8_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_8_lpi_1_dfm_24_22,
          Silu_for_y_8_lpi_1_dfm_4_24_22, Gelu_for_y_8_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_8_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_2_8_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_2_8_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_2015_cse ) begin
      act_regs_data_2_8_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_2_8_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[277:256]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_9_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_9_lpi_1_dfm_21_0,
          Silu_for_y_9_lpi_1_dfm_4_21_0_1, Gelu_for_y_9_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
      act_regs_data_2_8_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_2_8_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[281]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_9_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_9_lpi_1_dfm_25,
          Silu_for_y_9_lpi_1_dfm_4_25, Gelu_for_y_9_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
      act_regs_data_2_8_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_2_8_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[280:278]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_9_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_9_lpi_1_dfm_24_22,
          Silu_for_y_9_lpi_1_dfm_4_24_22, Gelu_for_y_9_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_9_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_2_9_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_2_9_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_2017_cse ) begin
      act_regs_data_2_9_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_2_9_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[309:288]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_10_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_10_lpi_1_dfm_21_0,
          Silu_for_y_10_lpi_1_dfm_4_21_0_1, Gelu_for_y_10_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
      act_regs_data_2_9_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_2_9_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[313]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_10_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_10_lpi_1_dfm_25,
          Silu_for_y_10_lpi_1_dfm_4_25, Gelu_for_y_10_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
      act_regs_data_2_9_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_2_9_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[312:310]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_10_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_10_lpi_1_dfm_24_22,
          Silu_for_y_10_lpi_1_dfm_4_24_22, Gelu_for_y_10_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_10_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_2_10_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_2_10_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_2019_cse ) begin
      act_regs_data_2_10_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_2_10_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[341:320]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_11_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_11_lpi_1_dfm_21_0,
          Silu_for_y_11_lpi_1_dfm_4_21_0_1, Gelu_for_y_11_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
      act_regs_data_2_10_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_2_10_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[345]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_11_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_11_lpi_1_dfm_25,
          Silu_for_y_11_lpi_1_dfm_4_25, Gelu_for_y_11_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
      act_regs_data_2_10_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_2_10_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[344:342]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_11_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_11_lpi_1_dfm_24_22,
          Silu_for_y_11_lpi_1_dfm_4_24_22, Gelu_for_y_11_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_11_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_2_11_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_2_11_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_2021_cse ) begin
      act_regs_data_2_11_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_2_11_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[373:352]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_12_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_12_lpi_1_dfm_21_0,
          Silu_for_y_12_lpi_1_dfm_4_21_0_1, Gelu_for_y_12_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
      act_regs_data_2_11_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_2_11_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[377]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_12_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_12_lpi_1_dfm_25,
          Silu_for_y_12_lpi_1_dfm_4_25, Gelu_for_y_12_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
      act_regs_data_2_11_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_2_11_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[376:374]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_12_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_12_lpi_1_dfm_24_22,
          Silu_for_y_12_lpi_1_dfm_4_24_22, Gelu_for_y_12_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_12_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_2_12_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_2_12_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_2023_cse ) begin
      act_regs_data_2_12_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_2_12_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[405:384]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_13_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_13_lpi_1_dfm_21_0,
          Silu_for_y_13_lpi_1_dfm_4_21_0_1, Gelu_for_y_13_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
      act_regs_data_2_12_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_2_12_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[409]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_13_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_13_lpi_1_dfm_25,
          Silu_for_y_13_lpi_1_dfm_4_25, Gelu_for_y_13_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
      act_regs_data_2_12_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_2_12_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[408:406]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_13_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_13_lpi_1_dfm_24_22,
          Silu_for_y_13_lpi_1_dfm_4_24_22, Gelu_for_y_13_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_13_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_2_13_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_2_13_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_2025_cse ) begin
      act_regs_data_2_13_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_2_13_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[437:416]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_14_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_14_lpi_1_dfm_21_0,
          Silu_for_y_14_lpi_1_dfm_4_21_0_1, Gelu_for_y_14_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
      act_regs_data_2_13_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_2_13_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[441]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_14_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_14_lpi_1_dfm_25,
          Silu_for_y_14_lpi_1_dfm_4_25, Gelu_for_y_14_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
      act_regs_data_2_13_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_2_13_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[440:438]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_14_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_14_lpi_1_dfm_24_22,
          Silu_for_y_14_lpi_1_dfm_4_24_22, Gelu_for_y_14_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_14_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_2_14_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_2_14_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_2027_cse ) begin
      act_regs_data_2_14_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_2_14_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[469:448]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_15_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_15_lpi_1_dfm_21_0,
          Silu_for_y_15_lpi_1_dfm_4_21_0_1, Gelu_for_y_15_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
      act_regs_data_2_14_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_2_14_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[473]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_15_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_15_lpi_1_dfm_25,
          Silu_for_y_15_lpi_1_dfm_4_25, Gelu_for_y_15_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
      act_regs_data_2_14_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_2_14_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[472:470]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_15_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_15_lpi_1_dfm_24_22,
          Silu_for_y_15_lpi_1_dfm_4_24_22, Gelu_for_y_15_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_15_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_2_15_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_2_15_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_2029_cse ) begin
      act_regs_data_2_15_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_2_15_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[501:480]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_lpi_1_dfm_21_0, Silu_for_y_lpi_1_dfm_4_21_0_1,
          Gelu_for_y_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
      act_regs_data_2_15_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_2_15_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[505]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_lpi_1_dfm_25, Silu_for_y_lpi_1_dfm_4_25,
          Gelu_for_y_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
      act_regs_data_2_15_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_2_15_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[504:502]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_lpi_1_dfm_24_22,
          Silu_for_y_lpi_1_dfm_4_24_22, Gelu_for_y_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_0_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_3_0_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_3_0_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_2031_cse ) begin
      act_regs_data_3_0_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_3_0_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[21:0]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_1_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_1_lpi_1_dfm_21_0,
          Silu_for_y_1_lpi_1_dfm_4_21_0, Gelu_for_y_1_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
      act_regs_data_3_0_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_3_0_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[25]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_1_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_1_lpi_1_dfm_25,
          Silu_for_y_1_lpi_1_dfm_4_25, Gelu_for_y_1_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
      act_regs_data_3_0_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_3_0_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[24:22]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_1_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_1_lpi_1_dfm_24_22,
          Silu_for_y_1_lpi_1_dfm_4_24_22, Gelu_for_y_1_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_1_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_3_1_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_3_1_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_2033_cse ) begin
      act_regs_data_3_1_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_3_1_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[53:32]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_2_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_2_lpi_1_dfm_21_0,
          Silu_for_y_2_lpi_1_dfm_4_21_0, Gelu_for_y_2_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
      act_regs_data_3_1_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_3_1_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[57]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_2_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_2_lpi_1_dfm_25,
          Silu_for_y_2_lpi_1_dfm_4_25, Gelu_for_y_2_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
      act_regs_data_3_1_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_3_1_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[56:54]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_2_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_2_lpi_1_dfm_24_22,
          Silu_for_y_2_lpi_1_dfm_4_24_22, Gelu_for_y_2_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_2_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_3_2_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_3_2_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_2035_cse ) begin
      act_regs_data_3_2_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_3_2_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[85:64]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_3_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_3_lpi_1_dfm_21_0,
          Silu_for_y_3_lpi_1_dfm_4_21_0, Gelu_for_y_3_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
      act_regs_data_3_2_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_3_2_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[89]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_3_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_3_lpi_1_dfm_25,
          Silu_for_y_3_lpi_1_dfm_4_25, Gelu_for_y_3_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
      act_regs_data_3_2_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_3_2_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[88:86]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_3_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_3_lpi_1_dfm_24_22,
          Silu_for_y_3_lpi_1_dfm_4_24_22, Gelu_for_y_3_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_3_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_3_3_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_3_3_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_2037_cse ) begin
      act_regs_data_3_3_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_3_3_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[117:96]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_4_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_4_lpi_1_dfm_21_0,
          Silu_for_y_4_lpi_1_dfm_4_21_0, Gelu_for_y_4_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
      act_regs_data_3_3_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_3_3_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[121]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_4_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_4_lpi_1_dfm_25,
          Silu_for_y_4_lpi_1_dfm_4_25, Gelu_for_y_4_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
      act_regs_data_3_3_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_3_3_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[120:118]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_4_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_4_lpi_1_dfm_24_22,
          Silu_for_y_4_lpi_1_dfm_4_24_22, Gelu_for_y_4_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_4_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_3_4_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_3_4_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_2039_cse ) begin
      act_regs_data_3_4_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_3_4_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[149:128]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_5_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_5_lpi_1_dfm_21_0,
          Silu_for_y_5_lpi_1_dfm_4_21_0, Gelu_for_y_5_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
      act_regs_data_3_4_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_3_4_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[153]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_5_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_5_lpi_1_dfm_25,
          Silu_for_y_5_lpi_1_dfm_4_25, Gelu_for_y_5_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
      act_regs_data_3_4_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_3_4_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[152:150]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_5_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_5_lpi_1_dfm_24_22,
          Silu_for_y_5_lpi_1_dfm_4_24_22, Gelu_for_y_5_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_5_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_3_5_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_3_5_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_2041_cse ) begin
      act_regs_data_3_5_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_3_5_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[181:160]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_6_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_6_lpi_1_dfm_21_0,
          Silu_for_y_6_lpi_1_dfm_4_21_0, Gelu_for_y_6_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
      act_regs_data_3_5_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_3_5_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[185]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_6_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_6_lpi_1_dfm_25,
          Silu_for_y_6_lpi_1_dfm_4_25, Gelu_for_y_6_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
      act_regs_data_3_5_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_3_5_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[184:182]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_6_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_6_lpi_1_dfm_24_22,
          Silu_for_y_6_lpi_1_dfm_4_24_22, Gelu_for_y_6_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_6_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_3_6_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_3_6_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_2043_cse ) begin
      act_regs_data_3_6_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_3_6_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[213:192]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_7_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_7_lpi_1_dfm_21_0,
          Silu_for_y_7_lpi_1_dfm_4_21_0, Gelu_for_y_7_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
      act_regs_data_3_6_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_3_6_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[217]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_7_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_7_lpi_1_dfm_25,
          Silu_for_y_7_lpi_1_dfm_4_25, Gelu_for_y_7_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
      act_regs_data_3_6_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_3_6_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[216:214]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_7_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_7_lpi_1_dfm_24_22,
          Silu_for_y_7_lpi_1_dfm_4_24_22, Gelu_for_y_7_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_7_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_3_7_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_3_7_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_2045_cse ) begin
      act_regs_data_3_7_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_3_7_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[245:224]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_8_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_8_lpi_1_dfm_21_0,
          Silu_for_y_8_lpi_1_dfm_4_21_0, Gelu_for_y_8_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
      act_regs_data_3_7_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_3_7_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[249]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_8_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_8_lpi_1_dfm_25,
          Silu_for_y_8_lpi_1_dfm_4_25, Gelu_for_y_8_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
      act_regs_data_3_7_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_3_7_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[248:246]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_8_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_8_lpi_1_dfm_24_22,
          Silu_for_y_8_lpi_1_dfm_4_24_22, Gelu_for_y_8_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_8_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_3_8_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_3_8_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_2047_cse ) begin
      act_regs_data_3_8_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_3_8_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[277:256]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_9_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_9_lpi_1_dfm_21_0,
          Silu_for_y_9_lpi_1_dfm_4_21_0_1, Gelu_for_y_9_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
      act_regs_data_3_8_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_3_8_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[281]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_9_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_9_lpi_1_dfm_25,
          Silu_for_y_9_lpi_1_dfm_4_25, Gelu_for_y_9_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
      act_regs_data_3_8_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_3_8_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[280:278]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_9_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_9_lpi_1_dfm_24_22,
          Silu_for_y_9_lpi_1_dfm_4_24_22, Gelu_for_y_9_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_9_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_3_9_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_3_9_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_2049_cse ) begin
      act_regs_data_3_9_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_3_9_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[309:288]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_10_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_10_lpi_1_dfm_21_0,
          Silu_for_y_10_lpi_1_dfm_4_21_0_1, Gelu_for_y_10_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
      act_regs_data_3_9_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_3_9_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[313]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_10_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_10_lpi_1_dfm_25,
          Silu_for_y_10_lpi_1_dfm_4_25, Gelu_for_y_10_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
      act_regs_data_3_9_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_3_9_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[312:310]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_10_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_10_lpi_1_dfm_24_22,
          Silu_for_y_10_lpi_1_dfm_4_24_22, Gelu_for_y_10_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_10_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_3_10_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_3_10_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_2051_cse ) begin
      act_regs_data_3_10_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_3_10_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[341:320]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_11_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_11_lpi_1_dfm_21_0,
          Silu_for_y_11_lpi_1_dfm_4_21_0_1, Gelu_for_y_11_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
      act_regs_data_3_10_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_3_10_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[345]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_11_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_11_lpi_1_dfm_25,
          Silu_for_y_11_lpi_1_dfm_4_25, Gelu_for_y_11_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
      act_regs_data_3_10_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_3_10_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[344:342]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_11_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_11_lpi_1_dfm_24_22,
          Silu_for_y_11_lpi_1_dfm_4_24_22, Gelu_for_y_11_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_11_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_3_11_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_3_11_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_2053_cse ) begin
      act_regs_data_3_11_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_3_11_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[373:352]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_12_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_12_lpi_1_dfm_21_0,
          Silu_for_y_12_lpi_1_dfm_4_21_0_1, Gelu_for_y_12_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
      act_regs_data_3_11_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_3_11_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[377]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_12_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_12_lpi_1_dfm_25,
          Silu_for_y_12_lpi_1_dfm_4_25, Gelu_for_y_12_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
      act_regs_data_3_11_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_3_11_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[376:374]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_12_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_12_lpi_1_dfm_24_22,
          Silu_for_y_12_lpi_1_dfm_4_24_22, Gelu_for_y_12_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_12_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_3_12_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_3_12_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_2055_cse ) begin
      act_regs_data_3_12_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_3_12_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[405:384]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_13_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_13_lpi_1_dfm_21_0,
          Silu_for_y_13_lpi_1_dfm_4_21_0_1, Gelu_for_y_13_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
      act_regs_data_3_12_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_3_12_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[409]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_13_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_13_lpi_1_dfm_25,
          Silu_for_y_13_lpi_1_dfm_4_25, Gelu_for_y_13_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
      act_regs_data_3_12_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_3_12_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[408:406]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_13_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_13_lpi_1_dfm_24_22,
          Silu_for_y_13_lpi_1_dfm_4_24_22, Gelu_for_y_13_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_13_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_3_13_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_3_13_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_2057_cse ) begin
      act_regs_data_3_13_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_3_13_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[437:416]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_14_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_14_lpi_1_dfm_21_0,
          Silu_for_y_14_lpi_1_dfm_4_21_0_1, Gelu_for_y_14_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
      act_regs_data_3_13_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_3_13_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[441]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_14_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_14_lpi_1_dfm_25,
          Silu_for_y_14_lpi_1_dfm_4_25, Gelu_for_y_14_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
      act_regs_data_3_13_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_3_13_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[440:438]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_14_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_14_lpi_1_dfm_24_22,
          Silu_for_y_14_lpi_1_dfm_4_24_22, Gelu_for_y_14_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_14_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_3_14_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_3_14_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_2059_cse ) begin
      act_regs_data_3_14_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_3_14_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[469:448]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_15_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_15_lpi_1_dfm_21_0,
          Silu_for_y_15_lpi_1_dfm_4_21_0_1, Gelu_for_y_15_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
      act_regs_data_3_14_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_3_14_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[473]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_15_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_15_lpi_1_dfm_25,
          Silu_for_y_15_lpi_1_dfm_4_25, Gelu_for_y_15_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
      act_regs_data_3_14_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_3_14_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[472:470]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_15_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_15_lpi_1_dfm_24_22,
          Silu_for_y_15_lpi_1_dfm_4_24_22, Gelu_for_y_15_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_15_sva_dfm_2_21_0 <= 22'b0000000000000000000000;
      act_regs_data_3_15_sva_dfm_2_25_22_rsp_0 <= 1'b0;
      act_regs_data_3_15_sva_dfm_2_25_22_rsp_1 <= 3'b000;
    end
    else if ( and_2061_cse ) begin
      act_regs_data_3_15_sva_dfm_2_21_0 <= MUX1HOT_v_22_8_2(act_regs_data_3_15_sva_21_0,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[501:480]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_21_0,
          Tanh_for_y_25_0_lpi_1_dfm_1_21_0, Relu_for_y_qr_30_0_lpi_1_dfm_21_0, Silu_for_y_lpi_1_dfm_4_21_0_1,
          Gelu_for_y_lpi_1_dfm_4_21_0_1, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[21:0]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
      act_regs_data_3_15_sva_dfm_2_25_22_rsp_0 <= MUX1HOT_s_1_8_2(act_regs_data_3_15_sva_25,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[505]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25,
          reg_Tanh_for_y_25_0_lpi_1_dfm_1_ftd, Relu_for_y_qr_30_0_lpi_1_dfm_25, Silu_for_y_lpi_1_dfm_4_25,
          Gelu_for_y_lpi_1_dfm_4_25, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
      act_regs_data_3_15_sva_dfm_2_25_22_rsp_1 <= MUX1HOT_v_3_8_2(act_regs_data_3_15_sva_24_22,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[504:502]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22,
          reg_Tanh_for_y_25_0_lpi_1_dfm_1_ftd_1, Relu_for_y_qr_30_0_lpi_1_dfm_24_22,
          Silu_for_y_lpi_1_dfm_4_24_22, Gelu_for_y_lpi_1_dfm_4_24_22, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_0_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2063_tmp ) begin
      act_regs_data_0_0_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(reg_act_regs_data_0_0_ftd_1,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[30:26]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_1_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_1_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_1_lpi_1_dfm_30_26, ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_30_26,
          Gelu_for_y_1_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_1_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2065_tmp ) begin
      act_regs_data_0_1_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(reg_act_regs_data_0_1_ftd_1,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[62:58]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_2_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_2_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_2_lpi_1_dfm_30_26, ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_1_30_26,
          Gelu_for_y_2_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_2_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2067_tmp ) begin
      act_regs_data_0_2_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_0_2_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[94:90]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_3_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_3_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_3_lpi_1_dfm_30_26, rva_out_reg_data_71_64_sva_dfm_6_4_0,
          Gelu_for_y_3_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_3_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2069_tmp ) begin
      act_regs_data_0_3_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_0_3_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[126:122]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_4_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_4_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_4_lpi_1_dfm_30_26, ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_1_30_26,
          Gelu_for_y_4_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_4_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2071_tmp ) begin
      act_regs_data_0_4_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_0_4_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[158:154]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_5_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_5_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_5_lpi_1_dfm_30_26, ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_1_30_26,
          Gelu_for_y_5_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_5_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2073_tmp ) begin
      act_regs_data_0_5_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_0_5_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[190:186]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_6_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_6_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_6_lpi_1_dfm_30_26, ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_1_30_26,
          Gelu_for_y_6_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_6_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2075_tmp ) begin
      act_regs_data_0_6_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_0_6_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[222:218]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_7_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_7_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_7_lpi_1_dfm_30_26, ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_1_30_26,
          Gelu_for_y_7_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_7_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2077_tmp ) begin
      act_regs_data_0_7_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_0_7_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[254:250]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_8_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_8_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_8_lpi_1_dfm_30_26, ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_1_30_26,
          Gelu_for_y_8_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_8_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2079_tmp ) begin
      act_regs_data_0_8_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_0_8_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[286:282]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_9_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_9_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_9_lpi_1_dfm_30_26, Silu_for_y_9_lpi_1_dfm_4_30_26_1,
          Gelu_for_y_9_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_9_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2081_tmp ) begin
      act_regs_data_0_9_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_0_9_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[318:314]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_10_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_10_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_10_lpi_1_dfm_30_26, Silu_for_y_10_lpi_1_dfm_4_30_26_1,
          Gelu_for_y_10_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_10_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2083_tmp ) begin
      act_regs_data_0_10_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(reg_act_regs_data_0_10_ftd_1,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[350:346]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_11_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_11_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_11_lpi_1_dfm_30_26, Silu_for_y_11_lpi_1_dfm_4_30_26_1,
          Gelu_for_y_11_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_11_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2085_tmp ) begin
      act_regs_data_0_11_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(reg_act_regs_data_0_11_ftd_1,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[382:378]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_12_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_12_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_12_lpi_1_dfm_30_26, Silu_for_y_12_lpi_1_dfm_4_30_26_1,
          Gelu_for_y_12_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_12_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2087_tmp ) begin
      act_regs_data_0_12_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(reg_act_regs_data_0_12_ftd_1,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[414:410]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_13_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_13_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_13_lpi_1_dfm_30_26, Silu_for_y_13_lpi_1_dfm_4_30_26_1,
          Gelu_for_y_13_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_13_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2089_tmp ) begin
      act_regs_data_0_13_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(reg_act_regs_data_0_13_ftd_1,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[446:442]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_14_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_14_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_14_lpi_1_dfm_30_26, Silu_for_y_14_lpi_1_dfm_4_30_26_1,
          Gelu_for_y_14_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_14_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2091_tmp ) begin
      act_regs_data_0_14_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_0_14_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[478:474]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_15_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_15_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_15_lpi_1_dfm_30_26, Silu_for_y_15_lpi_1_dfm_4_30_26_1,
          Gelu_for_y_15_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_15_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2093_tmp ) begin
      act_regs_data_0_15_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_0_15_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[510:506]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_lpi_1_dfm_30_26, Silu_for_y_lpi_1_dfm_4_30_26_1, Gelu_for_y_lpi_1_dfm_4_30_26,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1186_cse , act_regs_data_and_1187_cse , act_regs_data_and_1188_cse
          , act_regs_data_and_1189_cse , act_regs_data_and_1190_cse , act_regs_data_and_1191_cse
          , act_regs_data_and_1192_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_0_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2095_tmp ) begin
      act_regs_data_1_0_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_1_0_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[30:26]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_1_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_1_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_1_lpi_1_dfm_30_26, ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_30_26,
          Gelu_for_y_1_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_1_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2097_tmp ) begin
      act_regs_data_1_1_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_1_1_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[62:58]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_2_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_2_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_2_lpi_1_dfm_30_26, ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_1_30_26,
          Gelu_for_y_2_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_2_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2099_tmp ) begin
      act_regs_data_1_2_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_1_2_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[94:90]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_3_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_3_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_3_lpi_1_dfm_30_26, rva_out_reg_data_71_64_sva_dfm_6_4_0,
          Gelu_for_y_3_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_3_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2101_tmp ) begin
      act_regs_data_1_3_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_1_3_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[126:122]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_4_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_4_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_4_lpi_1_dfm_30_26, ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_1_30_26,
          Gelu_for_y_4_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_4_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2103_tmp ) begin
      act_regs_data_1_4_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_1_4_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[158:154]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_5_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_5_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_5_lpi_1_dfm_30_26, ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_1_30_26,
          Gelu_for_y_5_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_5_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2105_tmp ) begin
      act_regs_data_1_5_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_1_5_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[190:186]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_6_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_6_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_6_lpi_1_dfm_30_26, ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_1_30_26,
          Gelu_for_y_6_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_6_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2107_tmp ) begin
      act_regs_data_1_6_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_1_6_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[222:218]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_7_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_7_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_7_lpi_1_dfm_30_26, ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_1_30_26,
          Gelu_for_y_7_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_7_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2109_tmp ) begin
      act_regs_data_1_7_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_1_7_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[254:250]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_8_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_8_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_8_lpi_1_dfm_30_26, ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_1_30_26,
          Gelu_for_y_8_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_8_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2111_tmp ) begin
      act_regs_data_1_8_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_1_8_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[286:282]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_9_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_9_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_9_lpi_1_dfm_30_26, Silu_for_y_9_lpi_1_dfm_4_30_26_1,
          Gelu_for_y_9_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_9_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2113_tmp ) begin
      act_regs_data_1_9_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_1_9_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[318:314]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_10_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_10_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_10_lpi_1_dfm_30_26, Silu_for_y_10_lpi_1_dfm_4_30_26_1,
          Gelu_for_y_10_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_10_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2115_tmp ) begin
      act_regs_data_1_10_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_1_10_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[350:346]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_11_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_11_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_11_lpi_1_dfm_30_26, Silu_for_y_11_lpi_1_dfm_4_30_26_1,
          Gelu_for_y_11_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_11_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2117_tmp ) begin
      act_regs_data_1_11_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_1_11_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[382:378]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_12_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_12_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_12_lpi_1_dfm_30_26, Silu_for_y_12_lpi_1_dfm_4_30_26_1,
          Gelu_for_y_12_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_12_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2119_tmp ) begin
      act_regs_data_1_12_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_1_12_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[414:410]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_13_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_13_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_13_lpi_1_dfm_30_26, Silu_for_y_13_lpi_1_dfm_4_30_26_1,
          Gelu_for_y_13_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_13_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2121_tmp ) begin
      act_regs_data_1_13_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_1_13_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[446:442]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_14_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_14_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_14_lpi_1_dfm_30_26, Silu_for_y_14_lpi_1_dfm_4_30_26_1,
          Gelu_for_y_14_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_14_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2123_tmp ) begin
      act_regs_data_1_14_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_1_14_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[478:474]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_15_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_15_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_15_lpi_1_dfm_30_26, Silu_for_y_15_lpi_1_dfm_4_30_26_1,
          Gelu_for_y_15_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_15_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2125_tmp ) begin
      act_regs_data_1_15_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_1_15_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[510:506]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_lpi_1_dfm_30_26, Silu_for_y_lpi_1_dfm_4_30_26_1, Gelu_for_y_lpi_1_dfm_4_30_26,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1298_cse , act_regs_data_and_1299_cse , act_regs_data_and_1300_cse
          , act_regs_data_and_1301_cse , act_regs_data_and_1302_cse , act_regs_data_and_1303_cse
          , act_regs_data_and_1304_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_0_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2127_tmp ) begin
      act_regs_data_2_0_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_2_0_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[30:26]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_1_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_1_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_1_lpi_1_dfm_30_26, ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_30_26,
          Gelu_for_y_1_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_1_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2129_tmp ) begin
      act_regs_data_2_1_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_2_1_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[62:58]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_2_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_2_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_2_lpi_1_dfm_30_26, ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_1_30_26,
          Gelu_for_y_2_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_2_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2131_tmp ) begin
      act_regs_data_2_2_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_2_2_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[94:90]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_3_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_3_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_3_lpi_1_dfm_30_26, rva_out_reg_data_71_64_sva_dfm_6_4_0,
          Gelu_for_y_3_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_3_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2133_tmp ) begin
      act_regs_data_2_3_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_2_3_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[126:122]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_4_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_4_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_4_lpi_1_dfm_30_26, ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_1_30_26,
          Gelu_for_y_4_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_4_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2135_tmp ) begin
      act_regs_data_2_4_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_2_4_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[158:154]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_5_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_5_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_5_lpi_1_dfm_30_26, ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_1_30_26,
          Gelu_for_y_5_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_5_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2137_tmp ) begin
      act_regs_data_2_5_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_2_5_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[190:186]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_6_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_6_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_6_lpi_1_dfm_30_26, ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_1_30_26,
          Gelu_for_y_6_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_6_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2139_tmp ) begin
      act_regs_data_2_6_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_2_6_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[222:218]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_7_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_7_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_7_lpi_1_dfm_30_26, ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_1_30_26,
          Gelu_for_y_7_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_7_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2141_tmp ) begin
      act_regs_data_2_7_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_2_7_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[254:250]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_8_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_8_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_8_lpi_1_dfm_30_26, ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_1_30_26,
          Gelu_for_y_8_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_8_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2143_tmp ) begin
      act_regs_data_2_8_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_2_8_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[286:282]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_9_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_9_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_9_lpi_1_dfm_30_26, Silu_for_y_9_lpi_1_dfm_4_30_26_1,
          Gelu_for_y_9_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_9_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2145_tmp ) begin
      act_regs_data_2_9_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_2_9_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[318:314]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_10_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_10_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_10_lpi_1_dfm_30_26, Silu_for_y_10_lpi_1_dfm_4_30_26_1,
          Gelu_for_y_10_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_10_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2147_tmp ) begin
      act_regs_data_2_10_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_2_10_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[350:346]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_11_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_11_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_11_lpi_1_dfm_30_26, Silu_for_y_11_lpi_1_dfm_4_30_26_1,
          Gelu_for_y_11_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_11_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2149_tmp ) begin
      act_regs_data_2_11_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_2_11_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[382:378]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_12_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_12_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_12_lpi_1_dfm_30_26, Silu_for_y_12_lpi_1_dfm_4_30_26_1,
          Gelu_for_y_12_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_12_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2151_tmp ) begin
      act_regs_data_2_12_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_2_12_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[414:410]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_13_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_13_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_13_lpi_1_dfm_30_26, Silu_for_y_13_lpi_1_dfm_4_30_26_1,
          Gelu_for_y_13_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_13_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2153_tmp ) begin
      act_regs_data_2_13_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_2_13_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[446:442]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_14_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_14_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_14_lpi_1_dfm_30_26, Silu_for_y_14_lpi_1_dfm_4_30_26_1,
          Gelu_for_y_14_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_14_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2155_tmp ) begin
      act_regs_data_2_14_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_2_14_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[478:474]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_15_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_15_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_15_lpi_1_dfm_30_26, Silu_for_y_15_lpi_1_dfm_4_30_26_1,
          Gelu_for_y_15_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_15_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2157_tmp ) begin
      act_regs_data_2_15_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_2_15_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[510:506]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_lpi_1_dfm_30_26, Silu_for_y_lpi_1_dfm_4_30_26_1, Gelu_for_y_lpi_1_dfm_4_30_26,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1410_cse , act_regs_data_and_1411_cse , act_regs_data_and_1412_cse
          , act_regs_data_and_1413_cse , act_regs_data_and_1414_cse , act_regs_data_and_1415_cse
          , act_regs_data_and_1416_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_0_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2159_tmp ) begin
      act_regs_data_3_0_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_3_0_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[30:26]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_1_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_1_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_1_lpi_1_dfm_30_26, ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_30_26,
          Gelu_for_y_1_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_1_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2161_tmp ) begin
      act_regs_data_3_1_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_3_1_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[62:58]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_2_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_2_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_2_lpi_1_dfm_30_26, ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_1_30_26,
          Gelu_for_y_2_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_2_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2163_tmp ) begin
      act_regs_data_3_2_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_3_2_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[94:90]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_3_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_3_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_3_lpi_1_dfm_30_26, rva_out_reg_data_71_64_sva_dfm_6_4_0,
          Gelu_for_y_3_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_3_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2165_tmp ) begin
      act_regs_data_3_3_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_3_3_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[126:122]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_4_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_4_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_4_lpi_1_dfm_30_26, ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_1_30_26,
          Gelu_for_y_4_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_4_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2167_tmp ) begin
      act_regs_data_3_4_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_3_4_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[158:154]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_5_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_5_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_5_lpi_1_dfm_30_26, ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_1_30_26,
          Gelu_for_y_5_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_5_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2169_tmp ) begin
      act_regs_data_3_5_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_3_5_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[190:186]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_6_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_6_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_6_lpi_1_dfm_30_26, ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_1_30_26,
          Gelu_for_y_6_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_6_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2171_tmp ) begin
      act_regs_data_3_6_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_3_6_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[222:218]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_7_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_7_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_7_lpi_1_dfm_30_26, ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_1_30_26,
          Gelu_for_y_7_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_7_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2173_tmp ) begin
      act_regs_data_3_7_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_3_7_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[254:250]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_8_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_8_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_8_lpi_1_dfm_30_26, ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_1_30_26,
          Gelu_for_y_8_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_8_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2175_tmp ) begin
      act_regs_data_3_8_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_3_8_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[286:282]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_9_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_9_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_9_lpi_1_dfm_30_26, Silu_for_y_9_lpi_1_dfm_4_30_26_1,
          Gelu_for_y_9_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_9_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2177_tmp ) begin
      act_regs_data_3_9_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_3_9_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[318:314]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_10_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_10_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_10_lpi_1_dfm_30_26, Silu_for_y_10_lpi_1_dfm_4_30_26_1,
          Gelu_for_y_10_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_10_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2179_tmp ) begin
      act_regs_data_3_10_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_3_10_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[350:346]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_11_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_11_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_11_lpi_1_dfm_30_26, Silu_for_y_11_lpi_1_dfm_4_30_26_1,
          Gelu_for_y_11_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_11_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2181_tmp ) begin
      act_regs_data_3_11_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_3_11_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[382:378]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_12_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_12_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_12_lpi_1_dfm_30_26, Silu_for_y_12_lpi_1_dfm_4_30_26_1,
          Gelu_for_y_12_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_12_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2183_tmp ) begin
      act_regs_data_3_12_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_3_12_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[414:410]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_13_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_13_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_13_lpi_1_dfm_30_26, Silu_for_y_13_lpi_1_dfm_4_30_26_1,
          Gelu_for_y_13_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_13_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2185_tmp ) begin
      act_regs_data_3_13_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_3_13_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[446:442]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_14_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_14_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_14_lpi_1_dfm_30_26, Silu_for_y_14_lpi_1_dfm_4_30_26_1,
          Gelu_for_y_14_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_14_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2187_tmp ) begin
      act_regs_data_3_14_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_3_14_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[478:474]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_15_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_15_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_15_lpi_1_dfm_30_26, Silu_for_y_15_lpi_1_dfm_4_30_26_1,
          Gelu_for_y_15_lpi_1_dfm_4_30_26, (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_15_sva_dfm_2_30_26 <= 5'b00000;
    end
    else if ( and_2189_tmp ) begin
      act_regs_data_3_15_sva_dfm_2_30_26 <= MUX1HOT_v_5_8_2(act_regs_data_3_15_sva_30_26,
          (ActUnit_RunInst_case_3_act_port_reg_data_sva[510:506]), nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_30_26,
          ({{4{reg_Tanh_for_y_25_0_lpi_1_dfm_1_ftd}}, reg_Tanh_for_y_25_0_lpi_1_dfm_1_ftd}),
          Relu_for_y_qr_30_0_lpi_1_dfm_30_26, Silu_for_y_lpi_1_dfm_4_30_26_1, Gelu_for_y_lpi_1_dfm_4_30_26,
          (ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[30:26]),
          {act_regs_data_and_1522_cse , act_regs_data_and_1523_cse , act_regs_data_and_1524_cse
          , act_regs_data_and_1525_cse , act_regs_data_and_1526_cse , act_regs_data_and_1527_cse
          , act_regs_data_and_1528_cse , and_dcpl_1246});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_get_slc_2U_NVUINT8_return_3_sva <= 2'b00;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp ) begin
      nvhls_get_slc_2U_NVUINT8_return_3_sva <= nvhls_get_slc_2U_NVUINT8_return_3_sva_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_config_InstIncr_if_act_config_InstIncr_if_if_nor_mdf_sva <= 1'b0;
    end
    else if ( ActUnitRun_wen & (~((~ is_start_sva) | (~ act_config_InstIncr_if_equal_1_tmp)
        | (operator_6_false_acc_tmp[6:5]!=2'b00))) & while_asn_262_itm & is_incr_lpi_1_dfm_1
        ) begin
      act_config_InstIncr_if_act_config_InstIncr_if_if_nor_mdf_sva <= act_config_InstIncr_if_act_config_InstIncr_if_if_nor_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_else_1_mux_1_itm <= 1'b0;
    end
    else if ( ActUnitRun_wen & while_asn_262_itm ) begin
      while_else_1_mux_1_itm <= MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4, act_config_InstIncr_mux_2_nl,
          is_incr_lpi_1_dfm_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_23_4_ftd_12
          <= 8'b00000000;
    end
    else if ( mux_1474_nl & (~((fsm_output[3]) | is_start_sva)) & ActUnitRun_wen
        & (fsm_output[2:0]==3'b011) ) begin
      reg_ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_23_4_ftd_12
          <= ActUnit_DecodeAxi_Connections_InBlocking_RVSink_spec_Axi_rvaCfg_Write_Connections_SYN_PORT_PopNB_rva_in_reg_addr_sva_23_4_mx1_tmp_7_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_13_ftd_1 <= 5'b00000;
    end
    else if ( act_regs_data_and_2749_enex5 ) begin
      reg_act_regs_data_0_13_ftd_1 <= MUX1HOT_v_5_3_2(act_regs_data_0_13_sva_dfm_2_30_26,
          ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_1_30_26, act_regs_data_0_13_sva_8_30_26,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_13_ftd_3 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2751_enex5 ) begin
      reg_act_regs_data_0_13_ftd_3 <= MUX1HOT_v_22_3_2(act_regs_data_0_13_sva_dfm_2_21_0,
          reg_Silu_for_16_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1,
          act_regs_data_0_13_sva_8_21_0, {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1
          , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_12_ftd_1 <= 5'b00000;
    end
    else if ( act_regs_data_and_2752_enex5 ) begin
      reg_act_regs_data_0_12_ftd_1 <= MUX1HOT_v_5_3_2(act_regs_data_0_12_sva_dfm_2_30_26,
          ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_1_30_26, act_regs_data_0_12_sva_8_30_26,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_12_ftd_3 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2754_enex5 ) begin
      reg_act_regs_data_0_12_ftd_3 <= MUX1HOT_v_22_3_2(act_regs_data_0_12_sva_dfm_2_21_0,
          reg_Silu_for_15_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1,
          act_regs_data_0_12_sva_8_21_0, {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1
          , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_11_ftd_1 <= 5'b00000;
    end
    else if ( act_regs_data_and_2755_enex5 ) begin
      reg_act_regs_data_0_11_ftd_1 <= MUX1HOT_v_5_3_2(act_regs_data_0_11_sva_dfm_2_30_26,
          ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_1_30_26, act_regs_data_0_11_sva_8_30_26,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_11_ftd_3 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2757_enex5 ) begin
      reg_act_regs_data_0_11_ftd_3 <= MUX1HOT_v_22_3_2(act_regs_data_0_11_sva_dfm_2_21_0,
          reg_Silu_for_14_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1,
          act_regs_data_0_11_sva_8_21_0, {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1
          , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_10_ftd_1 <= 5'b00000;
    end
    else if ( act_regs_data_and_2758_enex5 ) begin
      reg_act_regs_data_0_10_ftd_1 <= MUX1HOT_v_5_3_2(act_regs_data_0_10_sva_dfm_2_30_26,
          ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_1_30_26, act_regs_data_0_10_sva_8_30_26,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_10_ftd_3 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2760_enex5 ) begin
      reg_act_regs_data_0_10_ftd_3 <= MUX1HOT_v_22_3_2(act_regs_data_0_10_sva_dfm_2_21_0,
          reg_Silu_for_13_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1,
          act_regs_data_0_10_sva_8_21_0, {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1
          , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_1_ftd_1 <= 5'b00000;
    end
    else if ( act_regs_data_and_2761_enex5 ) begin
      reg_act_regs_data_0_1_ftd_1 <= MUX1HOT_v_5_3_2(act_regs_data_0_1_sva_dfm_2_30_26,
          rva_out_reg_data_71_64_sva_dfm_6_4_0, act_regs_data_0_1_sva_8_30_26, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_1_ftd_3 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2763_enex5 ) begin
      reg_act_regs_data_0_1_ftd_3 <= MUX1HOT_v_22_3_2(act_regs_data_0_1_sva_dfm_2_21_0,
          reg_Silu_for_12_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1,
          act_regs_data_0_1_sva_8_21_0, {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1
          , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_0_ftd_1 <= 5'b00000;
    end
    else if ( act_regs_data_and_2764_enex5 ) begin
      reg_act_regs_data_0_0_ftd_1 <= MUX1HOT_v_5_3_2(act_regs_data_0_0_sva_dfm_2_30_26,
          ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_1_30_26, act_regs_data_0_0_sva_8_30_26,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_0_ftd_3 <= 22'b0000000000000000000000;
    end
    else if ( act_regs_data_and_2766_enex5 ) begin
      reg_act_regs_data_0_0_ftd_3 <= MUX1HOT_v_22_3_2(act_regs_data_0_0_sva_dfm_2_21_0,
          reg_Silu_for_11_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1,
          act_regs_data_0_0_sva_8_21_0, {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1
          , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_RunInst_case_14_nv_scvector_cctor_data_0_1_ftd_1 <= 22'b0000000000000000000000;
    end
    else if ( ActUnit_RunInst_switch_lp_and_817_enex5 ) begin
      reg_ActUnit_RunInst_case_14_nv_scvector_cctor_data_0_1_ftd_1 <= nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_RunInst_case_14_nv_scvector_cctor_data_0_ftd_1_30_26 <= 5'b00000;
    end
    else if ( ActUnit_RunInst_switch_lp_and_818_enex5 ) begin
      reg_ActUnit_RunInst_case_14_nv_scvector_cctor_data_0_ftd_1_30_26 <= nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_2_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1
          <= 22'b0000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_15_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_2_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1
          <= nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_2_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          <= 5'b00000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_16_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_2_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          <= nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1
          <= 22'b0000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_18_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1
          <= nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          <= 5'b00000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_19_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          <= nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1
          <= 22'b0000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_21_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1
          <= nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          <= 5'b00000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_22_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          <= nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1
          <= 22'b0000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_24_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1
          <= nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          <= 5'b00000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_25_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          <= nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1
          <= 22'b0000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_27_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1
          <= nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          <= 5'b00000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_28_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          <= nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1
          <= 22'b0000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_30_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1
          <= nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          <= 5'b00000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_31_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          <= nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1
          <= 22'b0000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_33_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1
          <= nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          <= 5'b00000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_34_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          <= nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1
          <= 22'b0000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_36_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1
          <= nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          <= 5'b00000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_37_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          <= nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1
          <= 22'b0000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_39_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1
          <= nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          <= 5'b00000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_40_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          <= nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1
          <= 22'b0000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_42_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1
          <= nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          <= 5'b00000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_43_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          <= nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1
          <= 22'b0000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_45_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1
          <= nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          <= 5'b00000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_46_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          <= nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1
          <= 22'b0000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_48_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1
          <= nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          <= 5'b00000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_49_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          <= nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1
          <= 22'b0000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_51_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1
          <= nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          <= 5'b00000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_52_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          <= nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1
          <= 22'b0000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_54_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1
          <= nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          <= 5'b00000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_55_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          <= nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1
          <= 22'b0000000000000000000000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_57_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1
          <= nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_3_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          <= 5'b00000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_58_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26
          <= nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_1_itm;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Silu_for_10_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd
          <= 3'b000;
    end
    else if ( Silu_for_else_else_else_if_and_1_ssc & and_dcpl_9 & (~ (act_config_in_InstFetch_return_sva_7_2[2]))
        & Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
        & Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
        & Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
        & (~ operator_32_8_true_AC_TRN_AC_WRAP_3_less_6_tmp) ) begin
      reg_Silu_for_10_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd
          <= Silu_for_10_else_else_else_if_acc_itm_25_1_1[24:22];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Silu_for_10_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1
          <= 22'b0000000000000000000000;
    end
    else if ( Silu_for_else_else_else_if_and_1_ssc ) begin
      reg_Silu_for_10_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1
          <= MUX1HOT_v_22_3_2((Silu_for_10_else_else_else_if_acc_itm_25_1_1[21:0]),
          (Silu_for_1_else_if_Silu_for_else_if_mul_cmp_7_z[44:23]), ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_21_0_mx0w1,
          {and_dcpl_331 , and_dcpl_1112 , and_dcpl_1235});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Silu_for_11_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd
          <= 3'b000;
    end
    else if ( Silu_for_else_else_else_if_and_2_ssc & and_dcpl_9 & (~ (act_config_in_InstFetch_return_sva_7_2[2]))
        & Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
        & Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
        & (~ operator_32_8_true_AC_TRN_AC_WRAP_3_less_5_tmp) & Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
        ) begin
      reg_Silu_for_11_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd
          <= Silu_for_11_else_else_else_if_acc_itm_25_1_1[24:22];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Silu_for_11_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1
          <= 22'b0000000000000000000000;
    end
    else if ( Silu_for_else_else_else_if_and_tmp ) begin
      reg_Silu_for_11_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1
          <= MUX1HOT_v_22_4_2((Silu_for_11_else_else_else_if_acc_itm_25_1_1[21:0]),
          (Silu_for_1_else_if_Silu_for_else_if_mul_cmp_z[44:23]), ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_21_0_mx0w1,
          nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_122_nl, {(~
          Silu_for_else_else_else_if_or_13_rgt) , and_dcpl_1112 , and_dcpl_1390 ,
          and_dcpl_1236});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Silu_for_12_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd
          <= 3'b000;
    end
    else if ( Silu_for_else_else_else_if_and_3_ssc & and_dcpl_9 & (~ (act_config_in_InstFetch_return_sva_7_2[2]))
        & Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
        & Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
        & (~ operator_32_8_true_AC_TRN_AC_WRAP_3_less_4_tmp) & Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
        ) begin
      reg_Silu_for_12_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd
          <= Silu_for_12_else_else_else_if_acc_itm_25_1_1[24:22];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Silu_for_12_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1
          <= 22'b0000000000000000000000;
    end
    else if ( and_2324_tmp ) begin
      reg_Silu_for_12_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1
          <= MUX_v_22_2_2((Silu_for_12_else_else_else_if_acc_itm_25_1_1[21:0]), and_1777_nl,
          Silu_for_else_else_else_if_or_14_cse);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Silu_for_13_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd
          <= 3'b000;
    end
    else if ( Silu_for_else_else_else_if_and_3_ssc & and_dcpl_9 & (~ (act_config_in_InstFetch_return_sva_7_2[2]))
        & Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
        & Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
        & (~ operator_32_8_true_AC_TRN_AC_WRAP_3_less_3_tmp) & Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
        ) begin
      reg_Silu_for_13_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd
          <= Silu_for_13_else_else_else_if_acc_itm_25_1_1[24:22];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Silu_for_13_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1
          <= 22'b0000000000000000000000;
    end
    else if ( and_2325_tmp ) begin
      reg_Silu_for_13_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1
          <= MUX_v_22_2_2((Silu_for_13_else_else_else_if_acc_itm_25_1_1[21:0]), and_1782_nl,
          Silu_for_else_else_else_if_or_14_cse);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Silu_for_14_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd
          <= 3'b000;
    end
    else if ( Silu_for_else_else_else_if_and_3_ssc & and_dcpl_9 & (~ (act_config_in_InstFetch_return_sva_7_2[2]))
        & Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
        & Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
        & Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
        & (~ operator_32_8_true_AC_TRN_AC_WRAP_3_less_2_tmp) ) begin
      reg_Silu_for_14_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd
          <= Silu_for_14_else_else_else_if_acc_itm_25_1_1[24:22];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Silu_for_14_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1
          <= 22'b0000000000000000000000;
    end
    else if ( and_2326_tmp ) begin
      reg_Silu_for_14_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1
          <= MUX_v_22_2_2((Silu_for_14_else_else_else_if_acc_itm_25_1_1[21:0]), and_1786_nl,
          Silu_for_else_else_else_if_or_14_cse);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Silu_for_15_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd
          <= 3'b000;
    end
    else if ( Silu_for_else_else_else_if_and_3_ssc & and_dcpl_9 & (~ (act_config_in_InstFetch_return_sva_7_2[2]))
        & Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
        & Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
        & Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
        & (~ operator_32_8_true_AC_TRN_AC_WRAP_3_less_1_tmp) ) begin
      reg_Silu_for_15_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd
          <= Silu_for_15_else_else_else_if_acc_itm_25_1_1[24:22];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Silu_for_15_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1
          <= 22'b0000000000000000000000;
    end
    else if ( and_2327_tmp ) begin
      reg_Silu_for_15_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1
          <= MUX_v_22_2_2((Silu_for_15_else_else_else_if_acc_itm_25_1_1[21:0]), and_1790_nl,
          Silu_for_else_else_else_if_or_14_cse);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Silu_for_16_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd
          <= 3'b000;
    end
    else if ( Silu_for_else_else_else_if_and_3_ssc & and_dcpl_9 & (~ (act_config_in_InstFetch_return_sva_7_2[2]))
        & Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs
        & Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
        & Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs
        & (~ operator_32_8_true_AC_TRN_AC_WRAP_3_less_tmp) ) begin
      reg_Silu_for_16_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd
          <= Silu_for_16_else_else_else_if_acc_itm_25_1_1[24:22];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Silu_for_16_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1
          <= 22'b0000000000000000000000;
    end
    else if ( and_2328_tmp ) begin
      reg_Silu_for_16_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_ftd_1
          <= MUX_v_22_2_2((Silu_for_16_else_else_else_if_acc_itm_25_1_1[21:0]), and_1794_nl,
          Silu_for_else_else_else_if_or_14_cse);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2530_enex5 ) begin
      reg_is_start_enexo <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2530_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_15_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2189_tmp | act_regs_data_and_2530_enex5 ) begin
      reg_act_regs_data_3_15_sva_dfm_2_30_26_enexo <= and_2189_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2530_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_15_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2704_enex5 | act_regs_data_and_2530_enex5 ) begin
      reg_act_regs_data_3_15_sva_8_30_26_enexo <= act_regs_data_and_2704_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_2_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_180_cse | act_regs_data_and_2530_enex5 ) begin
      reg_act_regs_data_2_2_sva_8_30_26_enexo <= act_regs_data_and_180_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_1 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2531_enex5 ) begin
      reg_is_start_enexo_1 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_15_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_2061_cse | act_regs_data_and_2531_enex5 ) begin
      reg_act_regs_data_3_15_sva_dfm_2_25_22_enexo <= and_2061_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_1 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2531_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_1 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_1 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2531_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_1 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_15_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2705_enex5 | act_regs_data_and_2531_enex5 ) begin
      reg_act_regs_data_3_15_sva_8_25_22_enexo <= act_regs_data_and_2705_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_2_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_180_cse | act_regs_data_and_2531_enex5 ) begin
      reg_act_regs_data_2_2_sva_8_25_22_enexo <= act_regs_data_and_180_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_2 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2532_enex5 ) begin
      reg_is_start_enexo_2 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_2 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2532_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_2 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_15_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_2061_cse | act_regs_data_and_2532_enex5 ) begin
      reg_act_regs_data_3_15_sva_dfm_2_21_0_enexo <= and_2061_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_2 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2532_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_2 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_15_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2706_enex5 | act_regs_data_and_2532_enex5 ) begin
      reg_act_regs_data_3_15_sva_8_21_0_enexo <= act_regs_data_and_2706_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_2_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_180_cse | act_regs_data_and_2532_enex5 ) begin
      reg_act_regs_data_2_2_sva_8_21_0_enexo <= act_regs_data_and_180_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_3 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2533_enex5 ) begin
      reg_is_start_enexo_3 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_3 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2533_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_3 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_15_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_128_cse | act_regs_data_and_2533_enex5 ) begin
      reg_act_regs_data_2_15_sva_8_30_26_enexo <= act_regs_data_and_128_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_14_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2187_tmp | act_regs_data_and_2533_enex5 ) begin
      reg_act_regs_data_3_14_sva_dfm_2_30_26_enexo <= and_2187_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_3 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2533_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_3 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_14_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2707_enex5 | act_regs_data_and_2533_enex5 ) begin
      reg_act_regs_data_3_14_sva_8_30_26_enexo <= act_regs_data_and_2707_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_4 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2534_enex5 ) begin
      reg_is_start_enexo_4 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_14_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_2059_cse | act_regs_data_and_2534_enex5 ) begin
      reg_act_regs_data_3_14_sva_dfm_2_25_22_enexo <= and_2059_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_4 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2534_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_4 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_15_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_128_cse | act_regs_data_and_2534_enex5 ) begin
      reg_act_regs_data_2_15_sva_8_25_22_enexo <= act_regs_data_and_128_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_4 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2534_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_4 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_14_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2708_enex5 | act_regs_data_and_2534_enex5 ) begin
      reg_act_regs_data_3_14_sva_8_25_22_enexo <= act_regs_data_and_2708_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_5 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2535_enex5 ) begin
      reg_is_start_enexo_5 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_5 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2535_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_5 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_15_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_128_cse | act_regs_data_and_2535_enex5 ) begin
      reg_act_regs_data_2_15_sva_8_21_0_enexo <= act_regs_data_and_128_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_14_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_2059_cse | act_regs_data_and_2535_enex5 ) begin
      reg_act_regs_data_3_14_sva_dfm_2_21_0_enexo <= and_2059_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_5 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2535_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_5 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_14_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2709_enex5 | act_regs_data_and_2535_enex5 ) begin
      reg_act_regs_data_3_14_sva_8_21_0_enexo <= act_regs_data_and_2709_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_6 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2536_enex5 ) begin
      reg_is_start_enexo_6 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_6 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2536_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_6 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_14_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_132_cse | act_regs_data_and_2536_enex5 ) begin
      reg_act_regs_data_2_14_sva_8_30_26_enexo <= act_regs_data_and_132_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_13_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2185_tmp | act_regs_data_and_2536_enex5 ) begin
      reg_act_regs_data_3_13_sva_dfm_2_30_26_enexo <= and_2185_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_6 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2536_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_6 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_13_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2710_enex5 | act_regs_data_and_2536_enex5 ) begin
      reg_act_regs_data_3_13_sva_8_30_26_enexo <= act_regs_data_and_2710_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_7 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2537_enex5 ) begin
      reg_is_start_enexo_7 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_13_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_2057_cse | act_regs_data_and_2537_enex5 ) begin
      reg_act_regs_data_3_13_sva_dfm_2_25_22_enexo <= and_2057_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_7 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2537_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_7 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_14_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_132_cse | act_regs_data_and_2537_enex5 ) begin
      reg_act_regs_data_2_14_sva_8_25_22_enexo <= act_regs_data_and_132_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_7 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2537_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_7 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_13_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2711_enex5 | act_regs_data_and_2537_enex5 ) begin
      reg_act_regs_data_3_13_sva_8_25_22_enexo <= act_regs_data_and_2711_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_8 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2538_enex5 ) begin
      reg_is_start_enexo_8 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_8 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2538_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_8 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_14_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_132_cse | act_regs_data_and_2538_enex5 ) begin
      reg_act_regs_data_2_14_sva_8_21_0_enexo <= act_regs_data_and_132_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_13_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_2057_cse | act_regs_data_and_2538_enex5 ) begin
      reg_act_regs_data_3_13_sva_dfm_2_21_0_enexo <= and_2057_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_8 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2538_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_8 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_13_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2712_enex5 | act_regs_data_and_2538_enex5 ) begin
      reg_act_regs_data_3_13_sva_8_21_0_enexo <= act_regs_data_and_2712_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_9 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2539_enex5 ) begin
      reg_is_start_enexo_9 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_9 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2539_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_9 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_13_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_136_cse | act_regs_data_and_2539_enex5 ) begin
      reg_act_regs_data_2_13_sva_8_30_26_enexo <= act_regs_data_and_136_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_12_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2183_tmp | act_regs_data_and_2539_enex5 ) begin
      reg_act_regs_data_3_12_sva_dfm_2_30_26_enexo <= and_2183_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_9 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2539_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_9 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_12_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2713_enex5 | act_regs_data_and_2539_enex5 ) begin
      reg_act_regs_data_3_12_sva_8_30_26_enexo <= act_regs_data_and_2713_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_10 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2540_enex5 ) begin
      reg_is_start_enexo_10 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_12_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_2055_cse | act_regs_data_and_2540_enex5 ) begin
      reg_act_regs_data_3_12_sva_dfm_2_25_22_enexo <= and_2055_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_10 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2540_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_10 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_13_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_136_cse | act_regs_data_and_2540_enex5 ) begin
      reg_act_regs_data_2_13_sva_8_25_22_enexo <= act_regs_data_and_136_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_10 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2540_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_10 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_12_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2714_enex5 | act_regs_data_and_2540_enex5 ) begin
      reg_act_regs_data_3_12_sva_8_25_22_enexo <= act_regs_data_and_2714_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_11 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2541_enex5 ) begin
      reg_is_start_enexo_11 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_11 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2541_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_11 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_13_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_136_cse | act_regs_data_and_2541_enex5 ) begin
      reg_act_regs_data_2_13_sva_8_21_0_enexo <= act_regs_data_and_136_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_12_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_2055_cse | act_regs_data_and_2541_enex5 ) begin
      reg_act_regs_data_3_12_sva_dfm_2_21_0_enexo <= and_2055_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_11 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2541_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_11 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_12_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2715_enex5 | act_regs_data_and_2541_enex5 ) begin
      reg_act_regs_data_3_12_sva_8_21_0_enexo <= act_regs_data_and_2715_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_12 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2542_enex5 ) begin
      reg_is_start_enexo_12 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_12 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2542_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_12 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_12_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_140_cse | act_regs_data_and_2542_enex5 ) begin
      reg_act_regs_data_2_12_sva_8_30_26_enexo <= act_regs_data_and_140_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_11_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2181_tmp | act_regs_data_and_2542_enex5 ) begin
      reg_act_regs_data_3_11_sva_dfm_2_30_26_enexo <= and_2181_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_12 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2542_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_12 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_11_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2716_enex5 | act_regs_data_and_2542_enex5 ) begin
      reg_act_regs_data_3_11_sva_8_30_26_enexo <= act_regs_data_and_2716_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_13 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2543_enex5 ) begin
      reg_is_start_enexo_13 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_11_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_2053_cse | act_regs_data_and_2543_enex5 ) begin
      reg_act_regs_data_3_11_sva_dfm_2_25_22_enexo <= and_2053_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_13 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2543_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_13 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_12_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_140_cse | act_regs_data_and_2543_enex5 ) begin
      reg_act_regs_data_2_12_sva_8_25_22_enexo <= act_regs_data_and_140_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_13 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2543_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_13 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_11_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2717_enex5 | act_regs_data_and_2543_enex5 ) begin
      reg_act_regs_data_3_11_sva_8_25_22_enexo <= act_regs_data_and_2717_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_14 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2544_enex5 ) begin
      reg_is_start_enexo_14 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_14 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2544_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_14 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_12_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_140_cse | act_regs_data_and_2544_enex5 ) begin
      reg_act_regs_data_2_12_sva_8_21_0_enexo <= act_regs_data_and_140_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_11_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_2053_cse | act_regs_data_and_2544_enex5 ) begin
      reg_act_regs_data_3_11_sva_dfm_2_21_0_enexo <= and_2053_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_14 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2544_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_14 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_11_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2718_enex5 | act_regs_data_and_2544_enex5 ) begin
      reg_act_regs_data_3_11_sva_8_21_0_enexo <= act_regs_data_and_2718_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_15 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2545_enex5 ) begin
      reg_is_start_enexo_15 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_15 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2545_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_15 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_11_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_144_cse | act_regs_data_and_2545_enex5 ) begin
      reg_act_regs_data_2_11_sva_8_30_26_enexo <= act_regs_data_and_144_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_10_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2179_tmp | act_regs_data_and_2545_enex5 ) begin
      reg_act_regs_data_3_10_sva_dfm_2_30_26_enexo <= and_2179_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_15 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2545_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_15 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_10_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2719_enex5 | act_regs_data_and_2545_enex5 ) begin
      reg_act_regs_data_3_10_sva_8_30_26_enexo <= act_regs_data_and_2719_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_16 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2546_enex5 ) begin
      reg_is_start_enexo_16 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_10_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_2051_cse | act_regs_data_and_2546_enex5 ) begin
      reg_act_regs_data_3_10_sva_dfm_2_25_22_enexo <= and_2051_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_16 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2546_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_16 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_11_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_144_cse | act_regs_data_and_2546_enex5 ) begin
      reg_act_regs_data_2_11_sva_8_25_22_enexo <= act_regs_data_and_144_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_16 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2546_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_16 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_10_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2720_enex5 | act_regs_data_and_2546_enex5 ) begin
      reg_act_regs_data_3_10_sva_8_25_22_enexo <= act_regs_data_and_2720_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_17 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2547_enex5 ) begin
      reg_is_start_enexo_17 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_17 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2547_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_17 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_11_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_144_cse | act_regs_data_and_2547_enex5 ) begin
      reg_act_regs_data_2_11_sva_8_21_0_enexo <= act_regs_data_and_144_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_10_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_2051_cse | act_regs_data_and_2547_enex5 ) begin
      reg_act_regs_data_3_10_sva_dfm_2_21_0_enexo <= and_2051_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_17 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2547_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_17 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_10_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2721_enex5 | act_regs_data_and_2547_enex5 ) begin
      reg_act_regs_data_3_10_sva_8_21_0_enexo <= act_regs_data_and_2721_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_18 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2548_enex5 ) begin
      reg_is_start_enexo_18 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_18 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2548_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_18 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_0_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_124_cse | act_regs_data_and_2548_enex5 ) begin
      reg_act_regs_data_3_0_sva_8_30_26_enexo <= act_regs_data_and_124_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_9_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2177_tmp | act_regs_data_and_2548_enex5 ) begin
      reg_act_regs_data_3_9_sva_dfm_2_30_26_enexo <= and_2177_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_9_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2722_enex5 | act_regs_data_and_2548_enex5 ) begin
      reg_act_regs_data_3_9_sva_8_30_26_enexo <= act_regs_data_and_2722_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_18 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2548_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_18 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_19 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2549_enex5 ) begin
      reg_is_start_enexo_19 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_9_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_2049_cse | act_regs_data_and_2549_enex5 ) begin
      reg_act_regs_data_3_9_sva_dfm_2_25_22_enexo <= and_2049_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_19 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2549_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_19 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_0_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_124_cse | act_regs_data_and_2549_enex5 ) begin
      reg_act_regs_data_3_0_sva_8_25_22_enexo <= act_regs_data_and_124_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_9_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2723_enex5 | act_regs_data_and_2549_enex5 ) begin
      reg_act_regs_data_3_9_sva_8_25_22_enexo <= act_regs_data_and_2723_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_19 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2549_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_19 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_20 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2550_enex5 ) begin
      reg_is_start_enexo_20 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_20 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2550_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_20 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_0_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_124_cse | act_regs_data_and_2550_enex5 ) begin
      reg_act_regs_data_3_0_sva_8_21_0_enexo <= act_regs_data_and_124_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_9_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_2049_cse | act_regs_data_and_2550_enex5 ) begin
      reg_act_regs_data_3_9_sva_dfm_2_21_0_enexo <= and_2049_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_9_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2724_enex5 | act_regs_data_and_2550_enex5 ) begin
      reg_act_regs_data_3_9_sva_8_21_0_enexo <= act_regs_data_and_2724_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_20 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2550_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_20 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_21 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2551_enex5 ) begin
      reg_is_start_enexo_21 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_21 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2551_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_21 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_9_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_152_cse | act_regs_data_and_2551_enex5 ) begin
      reg_act_regs_data_2_9_sva_8_30_26_enexo <= act_regs_data_and_152_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_8_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2175_tmp | act_regs_data_and_2551_enex5 ) begin
      reg_act_regs_data_3_8_sva_dfm_2_30_26_enexo <= and_2175_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_8_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2725_enex5 | act_regs_data_and_2551_enex5 ) begin
      reg_act_regs_data_3_8_sva_8_30_26_enexo <= act_regs_data_and_2725_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_21 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2551_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_21 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_22 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2552_enex5 ) begin
      reg_is_start_enexo_22 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_8_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_2047_cse | act_regs_data_and_2552_enex5 ) begin
      reg_act_regs_data_3_8_sva_dfm_2_25_22_enexo <= and_2047_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_22 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2552_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_22 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_9_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_152_cse | act_regs_data_and_2552_enex5 ) begin
      reg_act_regs_data_2_9_sva_8_25_22_enexo <= act_regs_data_and_152_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_8_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2726_enex5 | act_regs_data_and_2552_enex5 ) begin
      reg_act_regs_data_3_8_sva_8_25_22_enexo <= act_regs_data_and_2726_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_22 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2552_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_22 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_23 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2553_enex5 ) begin
      reg_is_start_enexo_23 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_23 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2553_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_23 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_9_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_152_cse | act_regs_data_and_2553_enex5 ) begin
      reg_act_regs_data_2_9_sva_8_21_0_enexo <= act_regs_data_and_152_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_8_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_2047_cse | act_regs_data_and_2553_enex5 ) begin
      reg_act_regs_data_3_8_sva_dfm_2_21_0_enexo <= and_2047_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_8_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2727_enex5 | act_regs_data_and_2553_enex5 ) begin
      reg_act_regs_data_3_8_sva_8_21_0_enexo <= act_regs_data_and_2727_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_23 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2553_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_23 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_24 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2554_enex5 ) begin
      reg_is_start_enexo_24 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_24 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2554_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_24 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_8_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_156_cse | act_regs_data_and_2554_enex5 ) begin
      reg_act_regs_data_2_8_sva_8_30_26_enexo <= act_regs_data_and_156_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_7_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2173_tmp | act_regs_data_and_2554_enex5 ) begin
      reg_act_regs_data_3_7_sva_dfm_2_30_26_enexo <= and_2173_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_7_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2728_enex5 | act_regs_data_and_2554_enex5 ) begin
      reg_act_regs_data_3_7_sva_8_30_26_enexo <= act_regs_data_and_2728_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_24 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2554_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_24 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_25 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2555_enex5 ) begin
      reg_is_start_enexo_25 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_7_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_2045_cse | act_regs_data_and_2555_enex5 ) begin
      reg_act_regs_data_3_7_sva_dfm_2_25_22_enexo <= and_2045_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_25 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2555_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_25 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_8_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_156_cse | act_regs_data_and_2555_enex5 ) begin
      reg_act_regs_data_2_8_sva_8_25_22_enexo <= act_regs_data_and_156_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_7_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2729_enex5 | act_regs_data_and_2555_enex5 ) begin
      reg_act_regs_data_3_7_sva_8_25_22_enexo <= act_regs_data_and_2729_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_25 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2555_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_25 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_26 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2556_enex5 ) begin
      reg_is_start_enexo_26 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_26 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2556_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_26 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_8_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_156_cse | act_regs_data_and_2556_enex5 ) begin
      reg_act_regs_data_2_8_sva_8_21_0_enexo <= act_regs_data_and_156_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_7_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_2045_cse | act_regs_data_and_2556_enex5 ) begin
      reg_act_regs_data_3_7_sva_dfm_2_21_0_enexo <= and_2045_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_7_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2730_enex5 | act_regs_data_and_2556_enex5 ) begin
      reg_act_regs_data_3_7_sva_8_21_0_enexo <= act_regs_data_and_2730_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_26 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2556_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_26 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_27 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2557_enex5 ) begin
      reg_is_start_enexo_27 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_27 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2557_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_27 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_7_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_160_cse | act_regs_data_and_2557_enex5 ) begin
      reg_act_regs_data_2_7_sva_8_30_26_enexo <= act_regs_data_and_160_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_6_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2171_tmp | act_regs_data_and_2557_enex5 ) begin
      reg_act_regs_data_3_6_sva_dfm_2_30_26_enexo <= and_2171_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_6_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2731_enex5 | act_regs_data_and_2557_enex5 ) begin
      reg_act_regs_data_3_6_sva_8_30_26_enexo <= act_regs_data_and_2731_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_27 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2557_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_27 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_28 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2558_enex5 ) begin
      reg_is_start_enexo_28 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_6_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_2043_cse | act_regs_data_and_2558_enex5 ) begin
      reg_act_regs_data_3_6_sva_dfm_2_25_22_enexo <= and_2043_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_28 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2558_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_28 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_7_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_160_cse | act_regs_data_and_2558_enex5 ) begin
      reg_act_regs_data_2_7_sva_8_25_22_enexo <= act_regs_data_and_160_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_6_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2732_enex5 | act_regs_data_and_2558_enex5 ) begin
      reg_act_regs_data_3_6_sva_8_25_22_enexo <= act_regs_data_and_2732_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_28 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2558_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_28 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_29 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2559_enex5 ) begin
      reg_is_start_enexo_29 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_29 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2559_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_29 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_7_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_160_cse | act_regs_data_and_2559_enex5 ) begin
      reg_act_regs_data_2_7_sva_8_21_0_enexo <= act_regs_data_and_160_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_6_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_2043_cse | act_regs_data_and_2559_enex5 ) begin
      reg_act_regs_data_3_6_sva_dfm_2_21_0_enexo <= and_2043_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_6_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2733_enex5 | act_regs_data_and_2559_enex5 ) begin
      reg_act_regs_data_3_6_sva_8_21_0_enexo <= act_regs_data_and_2733_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_29 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2559_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_29 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_30 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2560_enex5 ) begin
      reg_is_start_enexo_30 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_30 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2560_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_30 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_6_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_164_cse | act_regs_data_and_2560_enex5 ) begin
      reg_act_regs_data_2_6_sva_8_30_26_enexo <= act_regs_data_and_164_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_5_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2169_tmp | act_regs_data_and_2560_enex5 ) begin
      reg_act_regs_data_3_5_sva_dfm_2_30_26_enexo <= and_2169_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_5_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2734_enex5 | act_regs_data_and_2560_enex5 ) begin
      reg_act_regs_data_3_5_sva_8_30_26_enexo <= act_regs_data_and_2734_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_30 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2560_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_30 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_31 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2561_enex5 ) begin
      reg_is_start_enexo_31 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_5_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_2041_cse | act_regs_data_and_2561_enex5 ) begin
      reg_act_regs_data_3_5_sva_dfm_2_25_22_enexo <= and_2041_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_31 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2561_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_31 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_6_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_164_cse | act_regs_data_and_2561_enex5 ) begin
      reg_act_regs_data_2_6_sva_8_25_22_enexo <= act_regs_data_and_164_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_5_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2735_enex5 | act_regs_data_and_2561_enex5 ) begin
      reg_act_regs_data_3_5_sva_8_25_22_enexo <= act_regs_data_and_2735_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_31 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2561_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_31 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_32 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2562_enex5 ) begin
      reg_is_start_enexo_32 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_32 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2562_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_32 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_6_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_164_cse | act_regs_data_and_2562_enex5 ) begin
      reg_act_regs_data_2_6_sva_8_21_0_enexo <= act_regs_data_and_164_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_5_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_2041_cse | act_regs_data_and_2562_enex5 ) begin
      reg_act_regs_data_3_5_sva_dfm_2_21_0_enexo <= and_2041_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_5_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2736_enex5 | act_regs_data_and_2562_enex5 ) begin
      reg_act_regs_data_3_5_sva_8_21_0_enexo <= act_regs_data_and_2736_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_32 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2562_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_32 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_33 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2563_enex5 ) begin
      reg_is_start_enexo_33 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_33 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2563_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_33 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_5_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_168_cse | act_regs_data_and_2563_enex5 ) begin
      reg_act_regs_data_2_5_sva_8_30_26_enexo <= act_regs_data_and_168_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_4_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2167_tmp | act_regs_data_and_2563_enex5 ) begin
      reg_act_regs_data_3_4_sva_dfm_2_30_26_enexo <= and_2167_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_4_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2737_enex5 | act_regs_data_and_2563_enex5 ) begin
      reg_act_regs_data_3_4_sva_8_30_26_enexo <= act_regs_data_and_2737_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_33 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2563_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_33 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_34 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2564_enex5 ) begin
      reg_is_start_enexo_34 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_4_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_2039_cse | act_regs_data_and_2564_enex5 ) begin
      reg_act_regs_data_3_4_sva_dfm_2_25_22_enexo <= and_2039_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_34 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2564_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_34 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_5_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_168_cse | act_regs_data_and_2564_enex5 ) begin
      reg_act_regs_data_2_5_sva_8_25_22_enexo <= act_regs_data_and_168_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_4_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2738_enex5 | act_regs_data_and_2564_enex5 ) begin
      reg_act_regs_data_3_4_sva_8_25_22_enexo <= act_regs_data_and_2738_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_34 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2564_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_34 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_35 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2565_enex5 ) begin
      reg_is_start_enexo_35 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_35 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2565_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_35 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_4_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_2039_cse | act_regs_data_and_2565_enex5 ) begin
      reg_act_regs_data_3_4_sva_dfm_2_21_0_enexo <= and_2039_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_4_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2739_enex5 | act_regs_data_and_2565_enex5 ) begin
      reg_act_regs_data_3_4_sva_8_21_0_enexo <= act_regs_data_and_2739_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_35 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2565_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_35 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_5_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_168_cse | act_regs_data_and_2565_enex5 ) begin
      reg_act_regs_data_2_5_sva_8_21_0_enexo <= act_regs_data_and_168_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_36 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2566_enex5 ) begin
      reg_is_start_enexo_36 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_36 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2566_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_36 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_3_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2165_tmp | act_regs_data_and_2566_enex5 ) begin
      reg_act_regs_data_3_3_sva_dfm_2_30_26_enexo <= and_2165_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_3_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2740_enex5 | act_regs_data_and_2566_enex5 ) begin
      reg_act_regs_data_3_3_sva_8_30_26_enexo <= act_regs_data_and_2740_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_36 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2566_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_36 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_4_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_172_cse | act_regs_data_and_2566_enex5 ) begin
      reg_act_regs_data_2_4_sva_8_30_26_enexo <= act_regs_data_and_172_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_37 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2567_enex5 ) begin
      reg_is_start_enexo_37 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_3_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_2037_cse | act_regs_data_and_2567_enex5 ) begin
      reg_act_regs_data_3_3_sva_dfm_2_25_22_enexo <= and_2037_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_37 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2567_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_37 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_3_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2741_enex5 | act_regs_data_and_2567_enex5 ) begin
      reg_act_regs_data_3_3_sva_8_25_22_enexo <= act_regs_data_and_2741_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_37 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2567_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_37 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_4_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_172_cse | act_regs_data_and_2567_enex5 ) begin
      reg_act_regs_data_2_4_sva_8_25_22_enexo <= act_regs_data_and_172_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_38 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2568_enex5 ) begin
      reg_is_start_enexo_38 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_38 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2568_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_38 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_3_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_2037_cse | act_regs_data_and_2568_enex5 ) begin
      reg_act_regs_data_3_3_sva_dfm_2_21_0_enexo <= and_2037_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_3_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2742_enex5 | act_regs_data_and_2568_enex5 ) begin
      reg_act_regs_data_3_3_sva_8_21_0_enexo <= act_regs_data_and_2742_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_38 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2568_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_38 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_4_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_172_cse | act_regs_data_and_2568_enex5 ) begin
      reg_act_regs_data_2_4_sva_8_21_0_enexo <= act_regs_data_and_172_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_39 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2569_enex5 ) begin
      reg_is_start_enexo_39 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_39 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2569_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_39 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_2_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2163_tmp | act_regs_data_and_2569_enex5 ) begin
      reg_act_regs_data_3_2_sva_dfm_2_30_26_enexo <= and_2163_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_2_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2743_enex5 | act_regs_data_and_2569_enex5 ) begin
      reg_act_regs_data_3_2_sva_8_30_26_enexo <= act_regs_data_and_2743_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_39 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2569_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_39 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_3_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_176_cse | act_regs_data_and_2569_enex5 ) begin
      reg_act_regs_data_2_3_sva_8_30_26_enexo <= act_regs_data_and_176_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_40 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2570_enex5 ) begin
      reg_is_start_enexo_40 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_2_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_2035_cse | act_regs_data_and_2570_enex5 ) begin
      reg_act_regs_data_3_2_sva_dfm_2_25_22_enexo <= and_2035_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_40 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2570_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_40 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_2_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2744_enex5 | act_regs_data_and_2570_enex5 ) begin
      reg_act_regs_data_3_2_sva_8_25_22_enexo <= act_regs_data_and_2744_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_40 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2570_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_40 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_3_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_176_cse | act_regs_data_and_2570_enex5 ) begin
      reg_act_regs_data_2_3_sva_8_25_22_enexo <= act_regs_data_and_176_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_41 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2571_enex5 ) begin
      reg_is_start_enexo_41 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_41 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2571_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_41 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_2_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_2035_cse | act_regs_data_and_2571_enex5 ) begin
      reg_act_regs_data_3_2_sva_dfm_2_21_0_enexo <= and_2035_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_2_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2745_enex5 | act_regs_data_and_2571_enex5 ) begin
      reg_act_regs_data_3_2_sva_8_21_0_enexo <= act_regs_data_and_2745_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_41 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2571_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_41 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_3_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_176_cse | act_regs_data_and_2571_enex5 ) begin
      reg_act_regs_data_2_3_sva_8_21_0_enexo <= act_regs_data_and_176_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_42 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2572_enex5 ) begin
      reg_is_start_enexo_42 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_42 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2572_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_42 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_10_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_148_cse | act_regs_data_and_2572_enex5 ) begin
      reg_act_regs_data_2_10_sva_8_30_26_enexo <= act_regs_data_and_148_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_1_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2161_tmp | act_regs_data_and_2572_enex5 ) begin
      reg_act_regs_data_3_1_sva_dfm_2_30_26_enexo <= and_2161_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_1_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2746_enex5 | act_regs_data_and_2572_enex5 ) begin
      reg_act_regs_data_3_1_sva_8_30_26_enexo <= act_regs_data_and_2746_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_42 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2572_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_42 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_43 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2573_enex5 ) begin
      reg_is_start_enexo_43 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_1_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_2033_cse | act_regs_data_and_2573_enex5 ) begin
      reg_act_regs_data_3_1_sva_dfm_2_25_22_enexo <= and_2033_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_43 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2573_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_43 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_10_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_148_cse | act_regs_data_and_2573_enex5 ) begin
      reg_act_regs_data_2_10_sva_8_25_22_enexo <= act_regs_data_and_148_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_1_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2747_enex5 | act_regs_data_and_2573_enex5 ) begin
      reg_act_regs_data_3_1_sva_8_25_22_enexo <= act_regs_data_and_2747_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_43 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2573_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_43 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_44 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2574_enex5 ) begin
      reg_is_start_enexo_44 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_44 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2574_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_44 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_10_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_148_cse | act_regs_data_and_2574_enex5 ) begin
      reg_act_regs_data_2_10_sva_8_21_0_enexo <= act_regs_data_and_148_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_1_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_2033_cse | act_regs_data_and_2574_enex5 ) begin
      reg_act_regs_data_3_1_sva_dfm_2_21_0_enexo <= and_2033_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_1_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2748_enex5 | act_regs_data_and_2574_enex5 ) begin
      reg_act_regs_data_3_1_sva_8_21_0_enexo <= act_regs_data_and_2748_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_44 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2574_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_44 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_45 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2575_enex5 ) begin
      reg_is_start_enexo_45 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_45 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2575_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_45 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_0_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_124_cse | act_regs_data_and_2575_enex5 ) begin
      reg_act_regs_data_3_0_sva_8_30_26_enexo_1 <= act_regs_data_and_124_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_0_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2159_tmp | act_regs_data_and_2575_enex5 ) begin
      reg_act_regs_data_3_0_sva_dfm_2_30_26_enexo <= and_2159_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_45 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2575_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_45 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_1_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_184_cse | act_regs_data_and_2575_enex5 ) begin
      reg_act_regs_data_2_1_sva_8_30_26_enexo <= act_regs_data_and_184_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_46 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2576_enex5 ) begin
      reg_is_start_enexo_46 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_0_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_2031_cse | act_regs_data_and_2576_enex5 ) begin
      reg_act_regs_data_3_0_sva_dfm_2_25_22_enexo <= and_2031_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_46 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2576_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_46 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_0_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_124_cse | act_regs_data_and_2576_enex5 ) begin
      reg_act_regs_data_3_0_sva_8_25_22_enexo_1 <= act_regs_data_and_124_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_46 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2576_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_46 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_1_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_184_cse | act_regs_data_and_2576_enex5 ) begin
      reg_act_regs_data_2_1_sva_8_25_22_enexo <= act_regs_data_and_184_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_47 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2577_enex5 ) begin
      reg_is_start_enexo_47 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_47 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2577_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_47 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_0_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_124_cse | act_regs_data_and_2577_enex5 ) begin
      reg_act_regs_data_3_0_sva_8_21_0_enexo_1 <= act_regs_data_and_124_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_0_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_2031_cse | act_regs_data_and_2577_enex5 ) begin
      reg_act_regs_data_3_0_sva_dfm_2_21_0_enexo <= and_2031_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_47 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2577_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_47 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_1_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_184_cse | act_regs_data_and_2577_enex5 ) begin
      reg_act_regs_data_2_1_sva_8_21_0_enexo <= act_regs_data_and_184_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_48 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2578_enex5 ) begin
      reg_is_start_enexo_48 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_48 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2578_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_48 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_2_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_244_cse | act_regs_data_and_2578_enex5 ) begin
      reg_act_regs_data_1_2_sva_8_30_26_enexo <= act_regs_data_and_244_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_15_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_128_cse | act_regs_data_and_2578_enex5 ) begin
      reg_act_regs_data_2_15_sva_8_30_26_enexo_1 <= act_regs_data_and_128_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_15_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2157_tmp | act_regs_data_and_2578_enex5 ) begin
      reg_act_regs_data_2_15_sva_dfm_2_30_26_enexo <= and_2157_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_48 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2578_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_48 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_49 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2579_enex5 ) begin
      reg_is_start_enexo_49 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_15_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_2029_cse | act_regs_data_and_2579_enex5 ) begin
      reg_act_regs_data_2_15_sva_dfm_2_25_22_enexo <= and_2029_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_49 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2579_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_49 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_2_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_244_cse | act_regs_data_and_2579_enex5 ) begin
      reg_act_regs_data_1_2_sva_8_25_22_enexo <= act_regs_data_and_244_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_15_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_128_cse | act_regs_data_and_2579_enex5 ) begin
      reg_act_regs_data_2_15_sva_8_25_22_enexo_1 <= act_regs_data_and_128_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_49 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2579_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_49 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_50 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2580_enex5 ) begin
      reg_is_start_enexo_50 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_50 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2580_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_50 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_2_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_244_cse | act_regs_data_and_2580_enex5 ) begin
      reg_act_regs_data_1_2_sva_8_21_0_enexo <= act_regs_data_and_244_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_15_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_128_cse | act_regs_data_and_2580_enex5 ) begin
      reg_act_regs_data_2_15_sva_8_21_0_enexo_1 <= act_regs_data_and_128_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_15_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_2029_cse | act_regs_data_and_2580_enex5 ) begin
      reg_act_regs_data_2_15_sva_dfm_2_21_0_enexo <= and_2029_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_50 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2580_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_50 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_51 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2581_enex5 ) begin
      reg_is_start_enexo_51 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_51 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2581_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_51 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_14_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_132_cse | act_regs_data_and_2581_enex5 ) begin
      reg_act_regs_data_2_14_sva_8_30_26_enexo_1 <= act_regs_data_and_132_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_14_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2155_tmp | act_regs_data_and_2581_enex5 ) begin
      reg_act_regs_data_2_14_sva_dfm_2_30_26_enexo <= and_2155_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_51 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2581_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_51 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_15_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_192_cse | act_regs_data_and_2581_enex5 ) begin
      reg_act_regs_data_1_15_sva_8_30_26_enexo <= act_regs_data_and_192_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_52 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2582_enex5 ) begin
      reg_is_start_enexo_52 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_14_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_2027_cse | act_regs_data_and_2582_enex5 ) begin
      reg_act_regs_data_2_14_sva_dfm_2_25_22_enexo <= and_2027_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_52 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2582_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_52 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_14_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_132_cse | act_regs_data_and_2582_enex5 ) begin
      reg_act_regs_data_2_14_sva_8_25_22_enexo_1 <= act_regs_data_and_132_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_52 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2582_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_52 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_15_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_192_cse | act_regs_data_and_2582_enex5 ) begin
      reg_act_regs_data_1_15_sva_8_25_22_enexo <= act_regs_data_and_192_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_53 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2583_enex5 ) begin
      reg_is_start_enexo_53 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_53 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2583_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_53 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_14_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_132_cse | act_regs_data_and_2583_enex5 ) begin
      reg_act_regs_data_2_14_sva_8_21_0_enexo_1 <= act_regs_data_and_132_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_14_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_2027_cse | act_regs_data_and_2583_enex5 ) begin
      reg_act_regs_data_2_14_sva_dfm_2_21_0_enexo <= and_2027_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_53 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2583_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_53 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_15_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_192_cse | act_regs_data_and_2583_enex5 ) begin
      reg_act_regs_data_1_15_sva_8_21_0_enexo <= act_regs_data_and_192_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_54 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2584_enex5 ) begin
      reg_is_start_enexo_54 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_54 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2584_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_54 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_13_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_136_cse | act_regs_data_and_2584_enex5 ) begin
      reg_act_regs_data_2_13_sva_8_30_26_enexo_1 <= act_regs_data_and_136_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_13_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2153_tmp | act_regs_data_and_2584_enex5 ) begin
      reg_act_regs_data_2_13_sva_dfm_2_30_26_enexo <= and_2153_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_54 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2584_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_54 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_14_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_196_cse | act_regs_data_and_2584_enex5 ) begin
      reg_act_regs_data_1_14_sva_8_30_26_enexo <= act_regs_data_and_196_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_55 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2585_enex5 ) begin
      reg_is_start_enexo_55 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_13_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_2025_cse | act_regs_data_and_2585_enex5 ) begin
      reg_act_regs_data_2_13_sva_dfm_2_25_22_enexo <= and_2025_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_55 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2585_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_55 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_13_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_136_cse | act_regs_data_and_2585_enex5 ) begin
      reg_act_regs_data_2_13_sva_8_25_22_enexo_1 <= act_regs_data_and_136_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_55 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2585_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_55 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_14_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_196_cse | act_regs_data_and_2585_enex5 ) begin
      reg_act_regs_data_1_14_sva_8_25_22_enexo <= act_regs_data_and_196_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_56 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2586_enex5 ) begin
      reg_is_start_enexo_56 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_56 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2586_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_56 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_13_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_136_cse | act_regs_data_and_2586_enex5 ) begin
      reg_act_regs_data_2_13_sva_8_21_0_enexo_1 <= act_regs_data_and_136_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_13_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_2025_cse | act_regs_data_and_2586_enex5 ) begin
      reg_act_regs_data_2_13_sva_dfm_2_21_0_enexo <= and_2025_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_56 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2586_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_56 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_14_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_196_cse | act_regs_data_and_2586_enex5 ) begin
      reg_act_regs_data_1_14_sva_8_21_0_enexo <= act_regs_data_and_196_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_57 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2587_enex5 ) begin
      reg_is_start_enexo_57 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_57 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2587_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_57 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_12_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_140_cse | act_regs_data_and_2587_enex5 ) begin
      reg_act_regs_data_2_12_sva_8_30_26_enexo_1 <= act_regs_data_and_140_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_12_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2151_tmp | act_regs_data_and_2587_enex5 ) begin
      reg_act_regs_data_2_12_sva_dfm_2_30_26_enexo <= and_2151_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_57 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2587_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_57 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_13_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_200_cse | act_regs_data_and_2587_enex5 ) begin
      reg_act_regs_data_1_13_sva_8_30_26_enexo <= act_regs_data_and_200_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_58 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2588_enex5 ) begin
      reg_is_start_enexo_58 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_12_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_2023_cse | act_regs_data_and_2588_enex5 ) begin
      reg_act_regs_data_2_12_sva_dfm_2_25_22_enexo <= and_2023_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_58 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2588_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_58 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_12_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_140_cse | act_regs_data_and_2588_enex5 ) begin
      reg_act_regs_data_2_12_sva_8_25_22_enexo_1 <= act_regs_data_and_140_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_58 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2588_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_58 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_13_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_200_cse | act_regs_data_and_2588_enex5 ) begin
      reg_act_regs_data_1_13_sva_8_25_22_enexo <= act_regs_data_and_200_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_59 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2589_enex5 ) begin
      reg_is_start_enexo_59 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_59 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2589_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_59 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_12_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_140_cse | act_regs_data_and_2589_enex5 ) begin
      reg_act_regs_data_2_12_sva_8_21_0_enexo_1 <= act_regs_data_and_140_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_12_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_2023_cse | act_regs_data_and_2589_enex5 ) begin
      reg_act_regs_data_2_12_sva_dfm_2_21_0_enexo <= and_2023_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_59 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2589_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_59 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_13_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_200_cse | act_regs_data_and_2589_enex5 ) begin
      reg_act_regs_data_1_13_sva_8_21_0_enexo <= act_regs_data_and_200_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_60 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2590_enex5 ) begin
      reg_is_start_enexo_60 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_60 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2590_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_60 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_11_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_144_cse | act_regs_data_and_2590_enex5 ) begin
      reg_act_regs_data_2_11_sva_8_30_26_enexo_1 <= act_regs_data_and_144_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_11_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2149_tmp | act_regs_data_and_2590_enex5 ) begin
      reg_act_regs_data_2_11_sva_dfm_2_30_26_enexo <= and_2149_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_60 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2590_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_60 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_12_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_204_cse | act_regs_data_and_2590_enex5 ) begin
      reg_act_regs_data_1_12_sva_8_30_26_enexo <= act_regs_data_and_204_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_61 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2591_enex5 ) begin
      reg_is_start_enexo_61 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_11_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_2021_cse | act_regs_data_and_2591_enex5 ) begin
      reg_act_regs_data_2_11_sva_dfm_2_25_22_enexo <= and_2021_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_61 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2591_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_61 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_11_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_144_cse | act_regs_data_and_2591_enex5 ) begin
      reg_act_regs_data_2_11_sva_8_25_22_enexo_1 <= act_regs_data_and_144_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_61 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2591_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_61 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_12_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_204_cse | act_regs_data_and_2591_enex5 ) begin
      reg_act_regs_data_1_12_sva_8_25_22_enexo <= act_regs_data_and_204_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_62 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2592_enex5 ) begin
      reg_is_start_enexo_62 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_62 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2592_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_62 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_11_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_144_cse | act_regs_data_and_2592_enex5 ) begin
      reg_act_regs_data_2_11_sva_8_21_0_enexo_1 <= act_regs_data_and_144_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_11_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_2021_cse | act_regs_data_and_2592_enex5 ) begin
      reg_act_regs_data_2_11_sva_dfm_2_21_0_enexo <= and_2021_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_62 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2592_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_62 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_12_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_204_cse | act_regs_data_and_2592_enex5 ) begin
      reg_act_regs_data_1_12_sva_8_21_0_enexo <= act_regs_data_and_204_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_63 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2593_enex5 ) begin
      reg_is_start_enexo_63 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_63 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2593_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_63 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_10_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_148_cse | act_regs_data_and_2593_enex5 ) begin
      reg_act_regs_data_2_10_sva_8_30_26_enexo_1 <= act_regs_data_and_148_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_10_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2147_tmp | act_regs_data_and_2593_enex5 ) begin
      reg_act_regs_data_2_10_sva_dfm_2_30_26_enexo <= and_2147_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_63 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2593_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_63 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_11_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_208_cse | act_regs_data_and_2593_enex5 ) begin
      reg_act_regs_data_1_11_sva_8_30_26_enexo <= act_regs_data_and_208_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_64 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2594_enex5 ) begin
      reg_is_start_enexo_64 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_10_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_2019_cse | act_regs_data_and_2594_enex5 ) begin
      reg_act_regs_data_2_10_sva_dfm_2_25_22_enexo <= and_2019_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_64 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2594_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_64 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_10_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_148_cse | act_regs_data_and_2594_enex5 ) begin
      reg_act_regs_data_2_10_sva_8_25_22_enexo_1 <= act_regs_data_and_148_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_64 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2594_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_64 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_11_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_208_cse | act_regs_data_and_2594_enex5 ) begin
      reg_act_regs_data_1_11_sva_8_25_22_enexo <= act_regs_data_and_208_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_65 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2595_enex5 ) begin
      reg_is_start_enexo_65 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_65 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2595_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_65 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_10_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_148_cse | act_regs_data_and_2595_enex5 ) begin
      reg_act_regs_data_2_10_sva_8_21_0_enexo_1 <= act_regs_data_and_148_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_10_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_2019_cse | act_regs_data_and_2595_enex5 ) begin
      reg_act_regs_data_2_10_sva_dfm_2_21_0_enexo <= and_2019_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_65 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2595_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_65 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_11_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_208_cse | act_regs_data_and_2595_enex5 ) begin
      reg_act_regs_data_1_11_sva_8_21_0_enexo <= act_regs_data_and_208_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_66 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2596_enex5 ) begin
      reg_is_start_enexo_66 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_66 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2596_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_66 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_9_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_152_cse | act_regs_data_and_2596_enex5 ) begin
      reg_act_regs_data_2_9_sva_8_30_26_enexo_1 <= act_regs_data_and_152_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_9_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2145_tmp | act_regs_data_and_2596_enex5 ) begin
      reg_act_regs_data_2_9_sva_dfm_2_30_26_enexo <= and_2145_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_66 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2596_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_66 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_0_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_188_cse | act_regs_data_and_2596_enex5 ) begin
      reg_act_regs_data_2_0_sva_8_30_26_enexo <= act_regs_data_and_188_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_67 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2597_enex5 ) begin
      reg_is_start_enexo_67 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_9_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_2017_cse | act_regs_data_and_2597_enex5 ) begin
      reg_act_regs_data_2_9_sva_dfm_2_25_22_enexo <= and_2017_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_67 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2597_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_67 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_9_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_152_cse | act_regs_data_and_2597_enex5 ) begin
      reg_act_regs_data_2_9_sva_8_25_22_enexo_1 <= act_regs_data_and_152_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_67 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2597_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_67 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_0_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_188_cse | act_regs_data_and_2597_enex5 ) begin
      reg_act_regs_data_2_0_sva_8_25_22_enexo <= act_regs_data_and_188_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_68 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2598_enex5 ) begin
      reg_is_start_enexo_68 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_68 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2598_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_68 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_9_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_152_cse | act_regs_data_and_2598_enex5 ) begin
      reg_act_regs_data_2_9_sva_8_21_0_enexo_1 <= act_regs_data_and_152_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_9_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_2017_cse | act_regs_data_and_2598_enex5 ) begin
      reg_act_regs_data_2_9_sva_dfm_2_21_0_enexo <= and_2017_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_68 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2598_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_68 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_0_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_188_cse | act_regs_data_and_2598_enex5 ) begin
      reg_act_regs_data_2_0_sva_8_21_0_enexo <= act_regs_data_and_188_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_69 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2599_enex5 ) begin
      reg_is_start_enexo_69 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_69 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2599_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_69 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_8_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_156_cse | act_regs_data_and_2599_enex5 ) begin
      reg_act_regs_data_2_8_sva_8_30_26_enexo_1 <= act_regs_data_and_156_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_8_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2143_tmp | act_regs_data_and_2599_enex5 ) begin
      reg_act_regs_data_2_8_sva_dfm_2_30_26_enexo <= and_2143_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_69 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2599_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_69 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_9_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_216_cse | act_regs_data_and_2599_enex5 ) begin
      reg_act_regs_data_1_9_sva_8_30_26_enexo <= act_regs_data_and_216_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_70 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2600_enex5 ) begin
      reg_is_start_enexo_70 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_8_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_2015_cse | act_regs_data_and_2600_enex5 ) begin
      reg_act_regs_data_2_8_sva_dfm_2_25_22_enexo <= and_2015_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_70 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2600_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_70 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_9_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_216_cse | act_regs_data_and_2600_enex5 ) begin
      reg_act_regs_data_1_9_sva_8_25_22_enexo <= act_regs_data_and_216_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_8_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_156_cse | act_regs_data_and_2600_enex5 ) begin
      reg_act_regs_data_2_8_sva_8_25_22_enexo_1 <= act_regs_data_and_156_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_70 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2600_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_70 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_71 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2601_enex5 ) begin
      reg_is_start_enexo_71 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_71 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2601_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_71 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_9_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_216_cse | act_regs_data_and_2601_enex5 ) begin
      reg_act_regs_data_1_9_sva_8_21_0_enexo <= act_regs_data_and_216_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_8_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_156_cse | act_regs_data_and_2601_enex5 ) begin
      reg_act_regs_data_2_8_sva_8_21_0_enexo_1 <= act_regs_data_and_156_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_8_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_2015_cse | act_regs_data_and_2601_enex5 ) begin
      reg_act_regs_data_2_8_sva_dfm_2_21_0_enexo <= and_2015_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_71 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2601_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_71 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_72 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2602_enex5 ) begin
      reg_is_start_enexo_72 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_72 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2602_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_72 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_8_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_220_cse | act_regs_data_and_2602_enex5 ) begin
      reg_act_regs_data_1_8_sva_8_30_26_enexo <= act_regs_data_and_220_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_7_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_160_cse | act_regs_data_and_2602_enex5 ) begin
      reg_act_regs_data_2_7_sva_8_30_26_enexo_1 <= act_regs_data_and_160_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_7_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2141_tmp | act_regs_data_and_2602_enex5 ) begin
      reg_act_regs_data_2_7_sva_dfm_2_30_26_enexo <= and_2141_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_72 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2602_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_72 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_73 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2603_enex5 ) begin
      reg_is_start_enexo_73 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_7_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_2013_cse | act_regs_data_and_2603_enex5 ) begin
      reg_act_regs_data_2_7_sva_dfm_2_25_22_enexo <= and_2013_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_73 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2603_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_73 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_8_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_220_cse | act_regs_data_and_2603_enex5 ) begin
      reg_act_regs_data_1_8_sva_8_25_22_enexo <= act_regs_data_and_220_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_7_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_160_cse | act_regs_data_and_2603_enex5 ) begin
      reg_act_regs_data_2_7_sva_8_25_22_enexo_1 <= act_regs_data_and_160_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_73 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2603_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_73 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_74 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2604_enex5 ) begin
      reg_is_start_enexo_74 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_74 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2604_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_74 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_8_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_220_cse | act_regs_data_and_2604_enex5 ) begin
      reg_act_regs_data_1_8_sva_8_21_0_enexo <= act_regs_data_and_220_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_7_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_160_cse | act_regs_data_and_2604_enex5 ) begin
      reg_act_regs_data_2_7_sva_8_21_0_enexo_1 <= act_regs_data_and_160_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_7_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_2013_cse | act_regs_data_and_2604_enex5 ) begin
      reg_act_regs_data_2_7_sva_dfm_2_21_0_enexo <= and_2013_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_74 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2604_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_74 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_75 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2605_enex5 ) begin
      reg_is_start_enexo_75 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_75 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2605_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_75 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_7_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_224_cse | act_regs_data_and_2605_enex5 ) begin
      reg_act_regs_data_1_7_sva_8_30_26_enexo <= act_regs_data_and_224_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_6_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_164_cse | act_regs_data_and_2605_enex5 ) begin
      reg_act_regs_data_2_6_sva_8_30_26_enexo_1 <= act_regs_data_and_164_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_6_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2139_tmp | act_regs_data_and_2605_enex5 ) begin
      reg_act_regs_data_2_6_sva_dfm_2_30_26_enexo <= and_2139_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_75 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2605_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_75 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_76 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2606_enex5 ) begin
      reg_is_start_enexo_76 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_6_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_2011_cse | act_regs_data_and_2606_enex5 ) begin
      reg_act_regs_data_2_6_sva_dfm_2_25_22_enexo <= and_2011_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_76 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2606_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_76 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_7_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_224_cse | act_regs_data_and_2606_enex5 ) begin
      reg_act_regs_data_1_7_sva_8_25_22_enexo <= act_regs_data_and_224_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_6_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_164_cse | act_regs_data_and_2606_enex5 ) begin
      reg_act_regs_data_2_6_sva_8_25_22_enexo_1 <= act_regs_data_and_164_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_76 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2606_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_76 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_77 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2607_enex5 ) begin
      reg_is_start_enexo_77 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_77 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2607_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_77 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_7_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_224_cse | act_regs_data_and_2607_enex5 ) begin
      reg_act_regs_data_1_7_sva_8_21_0_enexo <= act_regs_data_and_224_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_6_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_164_cse | act_regs_data_and_2607_enex5 ) begin
      reg_act_regs_data_2_6_sva_8_21_0_enexo_1 <= act_regs_data_and_164_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_6_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_2011_cse | act_regs_data_and_2607_enex5 ) begin
      reg_act_regs_data_2_6_sva_dfm_2_21_0_enexo <= and_2011_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_77 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2607_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_77 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_78 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2608_enex5 ) begin
      reg_is_start_enexo_78 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_78 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2608_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_78 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_6_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_228_cse | act_regs_data_and_2608_enex5 ) begin
      reg_act_regs_data_1_6_sva_8_30_26_enexo <= act_regs_data_and_228_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_5_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_168_cse | act_regs_data_and_2608_enex5 ) begin
      reg_act_regs_data_2_5_sva_8_30_26_enexo_1 <= act_regs_data_and_168_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_5_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2137_tmp | act_regs_data_and_2608_enex5 ) begin
      reg_act_regs_data_2_5_sva_dfm_2_30_26_enexo <= and_2137_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_78 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2608_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_78 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_79 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2609_enex5 ) begin
      reg_is_start_enexo_79 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_5_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_2009_cse | act_regs_data_and_2609_enex5 ) begin
      reg_act_regs_data_2_5_sva_dfm_2_25_22_enexo <= and_2009_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_79 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2609_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_79 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_6_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_228_cse | act_regs_data_and_2609_enex5 ) begin
      reg_act_regs_data_1_6_sva_8_25_22_enexo <= act_regs_data_and_228_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_5_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_168_cse | act_regs_data_and_2609_enex5 ) begin
      reg_act_regs_data_2_5_sva_8_25_22_enexo_1 <= act_regs_data_and_168_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_79 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2609_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_79 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_80 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2610_enex5 ) begin
      reg_is_start_enexo_80 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_80 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2610_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_80 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_6_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_228_cse | act_regs_data_and_2610_enex5 ) begin
      reg_act_regs_data_1_6_sva_8_21_0_enexo <= act_regs_data_and_228_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_5_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_2009_cse | act_regs_data_and_2610_enex5 ) begin
      reg_act_regs_data_2_5_sva_dfm_2_21_0_enexo <= and_2009_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_80 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2610_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_80 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_5_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_168_cse | act_regs_data_and_2610_enex5 ) begin
      reg_act_regs_data_2_5_sva_8_21_0_enexo_1 <= act_regs_data_and_168_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_81 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2611_enex5 ) begin
      reg_is_start_enexo_81 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_81 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2611_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_81 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_5_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_232_cse | act_regs_data_and_2611_enex5 ) begin
      reg_act_regs_data_1_5_sva_8_30_26_enexo <= act_regs_data_and_232_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_4_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2135_tmp | act_regs_data_and_2611_enex5 ) begin
      reg_act_regs_data_2_4_sva_dfm_2_30_26_enexo <= and_2135_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_81 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2611_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_81 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_4_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_172_cse | act_regs_data_and_2611_enex5 ) begin
      reg_act_regs_data_2_4_sva_8_30_26_enexo_1 <= act_regs_data_and_172_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_82 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2612_enex5 ) begin
      reg_is_start_enexo_82 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_4_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_2007_cse | act_regs_data_and_2612_enex5 ) begin
      reg_act_regs_data_2_4_sva_dfm_2_25_22_enexo <= and_2007_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_82 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2612_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_82 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_5_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_232_cse | act_regs_data_and_2612_enex5 ) begin
      reg_act_regs_data_1_5_sva_8_25_22_enexo <= act_regs_data_and_232_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_82 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2612_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_82 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_4_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_172_cse | act_regs_data_and_2612_enex5 ) begin
      reg_act_regs_data_2_4_sva_8_25_22_enexo_1 <= act_regs_data_and_172_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_83 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2613_enex5 ) begin
      reg_is_start_enexo_83 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_83 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2613_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_83 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_5_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_232_cse | act_regs_data_and_2613_enex5 ) begin
      reg_act_regs_data_1_5_sva_8_21_0_enexo <= act_regs_data_and_232_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_4_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_2007_cse | act_regs_data_and_2613_enex5 ) begin
      reg_act_regs_data_2_4_sva_dfm_2_21_0_enexo <= and_2007_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_83 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2613_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_83 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_4_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_172_cse | act_regs_data_and_2613_enex5 ) begin
      reg_act_regs_data_2_4_sva_8_21_0_enexo_1 <= act_regs_data_and_172_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_84 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2614_enex5 ) begin
      reg_is_start_enexo_84 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_84 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2614_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_84 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_4_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_236_cse | act_regs_data_and_2614_enex5 ) begin
      reg_act_regs_data_1_4_sva_8_30_26_enexo <= act_regs_data_and_236_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_3_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2133_tmp | act_regs_data_and_2614_enex5 ) begin
      reg_act_regs_data_2_3_sva_dfm_2_30_26_enexo <= and_2133_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_84 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2614_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_84 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_3_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_176_cse | act_regs_data_and_2614_enex5 ) begin
      reg_act_regs_data_2_3_sva_8_30_26_enexo_1 <= act_regs_data_and_176_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_85 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2615_enex5 ) begin
      reg_is_start_enexo_85 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_3_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_2005_cse | act_regs_data_and_2615_enex5 ) begin
      reg_act_regs_data_2_3_sva_dfm_2_25_22_enexo <= and_2005_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_85 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2615_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_85 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_4_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_236_cse | act_regs_data_and_2615_enex5 ) begin
      reg_act_regs_data_1_4_sva_8_25_22_enexo <= act_regs_data_and_236_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_85 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2615_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_85 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_3_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_176_cse | act_regs_data_and_2615_enex5 ) begin
      reg_act_regs_data_2_3_sva_8_25_22_enexo_1 <= act_regs_data_and_176_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_86 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2616_enex5 ) begin
      reg_is_start_enexo_86 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_86 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2616_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_86 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_4_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_236_cse | act_regs_data_and_2616_enex5 ) begin
      reg_act_regs_data_1_4_sva_8_21_0_enexo <= act_regs_data_and_236_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_3_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_2005_cse | act_regs_data_and_2616_enex5 ) begin
      reg_act_regs_data_2_3_sva_dfm_2_21_0_enexo <= and_2005_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_86 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2616_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_86 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_3_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_176_cse | act_regs_data_and_2616_enex5 ) begin
      reg_act_regs_data_2_3_sva_8_21_0_enexo_1 <= act_regs_data_and_176_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_87 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2617_enex5 ) begin
      reg_is_start_enexo_87 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_87 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2617_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_87 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_3_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_240_cse | act_regs_data_and_2617_enex5 ) begin
      reg_act_regs_data_1_3_sva_8_30_26_enexo <= act_regs_data_and_240_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_2_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2131_tmp | act_regs_data_and_2617_enex5 ) begin
      reg_act_regs_data_2_2_sva_dfm_2_30_26_enexo <= and_2131_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_87 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2617_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_87 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_2_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_180_cse | act_regs_data_and_2617_enex5 ) begin
      reg_act_regs_data_2_2_sva_8_30_26_enexo_1 <= act_regs_data_and_180_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_88 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2618_enex5 ) begin
      reg_is_start_enexo_88 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_2_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_2003_cse | act_regs_data_and_2618_enex5 ) begin
      reg_act_regs_data_2_2_sva_dfm_2_25_22_enexo <= and_2003_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_88 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2618_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_88 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_3_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_240_cse | act_regs_data_and_2618_enex5 ) begin
      reg_act_regs_data_1_3_sva_8_25_22_enexo <= act_regs_data_and_240_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_88 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2618_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_88 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_2_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_180_cse | act_regs_data_and_2618_enex5 ) begin
      reg_act_regs_data_2_2_sva_8_25_22_enexo_1 <= act_regs_data_and_180_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_89 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2619_enex5 ) begin
      reg_is_start_enexo_89 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_89 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2619_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_89 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_3_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_240_cse | act_regs_data_and_2619_enex5 ) begin
      reg_act_regs_data_1_3_sva_8_21_0_enexo <= act_regs_data_and_240_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_2_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_2003_cse | act_regs_data_and_2619_enex5 ) begin
      reg_act_regs_data_2_2_sva_dfm_2_21_0_enexo <= and_2003_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_89 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2619_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_89 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_2_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_180_cse | act_regs_data_and_2619_enex5 ) begin
      reg_act_regs_data_2_2_sva_8_21_0_enexo_1 <= act_regs_data_and_180_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_90 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2620_enex5 ) begin
      reg_is_start_enexo_90 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_90 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2620_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_90 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_1_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2129_tmp | act_regs_data_and_2620_enex5 ) begin
      reg_act_regs_data_2_1_sva_dfm_2_30_26_enexo <= and_2129_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_90 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2620_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_90 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_1_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_184_cse | act_regs_data_and_2620_enex5 ) begin
      reg_act_regs_data_2_1_sva_8_30_26_enexo_1 <= act_regs_data_and_184_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_10_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_212_cse | act_regs_data_and_2620_enex5 ) begin
      reg_act_regs_data_1_10_sva_8_30_26_enexo <= act_regs_data_and_212_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_91 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2621_enex5 ) begin
      reg_is_start_enexo_91 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_1_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_2001_cse | act_regs_data_and_2621_enex5 ) begin
      reg_act_regs_data_2_1_sva_dfm_2_25_22_enexo <= and_2001_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_91 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2621_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_91 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_91 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2621_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_91 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_1_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_184_cse | act_regs_data_and_2621_enex5 ) begin
      reg_act_regs_data_2_1_sva_8_25_22_enexo_1 <= act_regs_data_and_184_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_10_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_212_cse | act_regs_data_and_2621_enex5 ) begin
      reg_act_regs_data_1_10_sva_8_25_22_enexo <= act_regs_data_and_212_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_92 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2622_enex5 ) begin
      reg_is_start_enexo_92 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_92 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2622_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_92 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_1_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_2001_cse | act_regs_data_and_2622_enex5 ) begin
      reg_act_regs_data_2_1_sva_dfm_2_21_0_enexo <= and_2001_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_92 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2622_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_92 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_1_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_184_cse | act_regs_data_and_2622_enex5 ) begin
      reg_act_regs_data_2_1_sva_8_21_0_enexo_1 <= act_regs_data_and_184_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_10_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_212_cse | act_regs_data_and_2622_enex5 ) begin
      reg_act_regs_data_1_10_sva_8_21_0_enexo <= act_regs_data_and_212_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_93 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2623_enex5 ) begin
      reg_is_start_enexo_93 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_93 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2623_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_93 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_1_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_248_cse | act_regs_data_and_2623_enex5 ) begin
      reg_act_regs_data_1_1_sva_8_30_26_enexo <= act_regs_data_and_248_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_0_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2127_tmp | act_regs_data_and_2623_enex5 ) begin
      reg_act_regs_data_2_0_sva_dfm_2_30_26_enexo <= and_2127_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_93 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2623_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_93 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_0_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_188_cse | act_regs_data_and_2623_enex5 ) begin
      reg_act_regs_data_2_0_sva_8_30_26_enexo_1 <= act_regs_data_and_188_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_94 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2624_enex5 ) begin
      reg_is_start_enexo_94 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_0_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_1999_cse | act_regs_data_and_2624_enex5 ) begin
      reg_act_regs_data_2_0_sva_dfm_2_25_22_enexo <= and_1999_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_94 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2624_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_94 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_1_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_248_cse | act_regs_data_and_2624_enex5 ) begin
      reg_act_regs_data_1_1_sva_8_25_22_enexo <= act_regs_data_and_248_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_94 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2624_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_94 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_0_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_188_cse | act_regs_data_and_2624_enex5 ) begin
      reg_act_regs_data_2_0_sva_8_25_22_enexo_1 <= act_regs_data_and_188_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_95 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2625_enex5 ) begin
      reg_is_start_enexo_95 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_95 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2625_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_95 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_1_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_248_cse | act_regs_data_and_2625_enex5 ) begin
      reg_act_regs_data_1_1_sva_8_21_0_enexo <= act_regs_data_and_248_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_0_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_1999_cse | act_regs_data_and_2625_enex5 ) begin
      reg_act_regs_data_2_0_sva_dfm_2_21_0_enexo <= and_1999_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_95 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2625_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_95 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_0_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_188_cse | act_regs_data_and_2625_enex5 ) begin
      reg_act_regs_data_2_0_sva_8_21_0_enexo_1 <= act_regs_data_and_188_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_96 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2626_enex5 ) begin
      reg_is_start_enexo_96 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_2_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_308_cse | act_regs_data_and_2626_enex5 ) begin
      reg_act_regs_data_0_2_sva_8_30_26_enexo <= act_regs_data_and_308_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_96 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2626_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_96 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_15_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2125_tmp | act_regs_data_and_2626_enex5 ) begin
      reg_act_regs_data_1_15_sva_dfm_2_30_26_enexo <= and_2125_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_96 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2626_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_96 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_15_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_192_cse | act_regs_data_and_2626_enex5 ) begin
      reg_act_regs_data_1_15_sva_8_30_26_enexo_1 <= act_regs_data_and_192_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_97 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2627_enex5 ) begin
      reg_is_start_enexo_97 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_15_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_1997_cse | act_regs_data_and_2627_enex5 ) begin
      reg_act_regs_data_1_15_sva_dfm_2_25_22_enexo <= and_1997_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_2_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_308_cse | act_regs_data_and_2627_enex5 ) begin
      reg_act_regs_data_0_2_sva_8_25_22_enexo <= act_regs_data_and_308_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_97 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2627_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_97 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_97 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2627_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_97 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_15_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_192_cse | act_regs_data_and_2627_enex5 ) begin
      reg_act_regs_data_1_15_sva_8_25_22_enexo_1 <= act_regs_data_and_192_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_98 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2628_enex5 ) begin
      reg_is_start_enexo_98 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_2_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_308_cse | act_regs_data_and_2628_enex5 ) begin
      reg_act_regs_data_0_2_sva_8_21_0_enexo <= act_regs_data_and_308_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_98 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2628_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_98 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_15_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_1997_cse | act_regs_data_and_2628_enex5 ) begin
      reg_act_regs_data_1_15_sva_dfm_2_21_0_enexo <= and_1997_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_98 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2628_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_98 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_15_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_192_cse | act_regs_data_and_2628_enex5 ) begin
      reg_act_regs_data_1_15_sva_8_21_0_enexo_1 <= act_regs_data_and_192_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_99 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2629_enex5 ) begin
      reg_is_start_enexo_99 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_99 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2629_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_99 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_15_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_256_cse | act_regs_data_and_2629_enex5 ) begin
      reg_act_regs_data_0_15_sva_8_30_26_enexo <= act_regs_data_and_256_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_14_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2123_tmp | act_regs_data_and_2629_enex5 ) begin
      reg_act_regs_data_1_14_sva_dfm_2_30_26_enexo <= and_2123_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_99 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2629_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_99 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_14_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_196_cse | act_regs_data_and_2629_enex5 ) begin
      reg_act_regs_data_1_14_sva_8_30_26_enexo_1 <= act_regs_data_and_196_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_100 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2630_enex5 ) begin
      reg_is_start_enexo_100 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_14_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_1995_cse | act_regs_data_and_2630_enex5 ) begin
      reg_act_regs_data_1_14_sva_dfm_2_25_22_enexo <= and_1995_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_100 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2630_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_100 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_15_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_256_cse | act_regs_data_and_2630_enex5 ) begin
      reg_act_regs_data_0_15_sva_8_25_22_enexo <= act_regs_data_and_256_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_100 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2630_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_100 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_14_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_196_cse | act_regs_data_and_2630_enex5 ) begin
      reg_act_regs_data_1_14_sva_8_25_22_enexo_1 <= act_regs_data_and_196_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_101 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2631_enex5 ) begin
      reg_is_start_enexo_101 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_101 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2631_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_101 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_15_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_256_cse | act_regs_data_and_2631_enex5 ) begin
      reg_act_regs_data_0_15_sva_8_21_0_enexo <= act_regs_data_and_256_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_14_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_1995_cse | act_regs_data_and_2631_enex5 ) begin
      reg_act_regs_data_1_14_sva_dfm_2_21_0_enexo <= and_1995_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_101 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2631_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_101 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_14_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_196_cse | act_regs_data_and_2631_enex5 ) begin
      reg_act_regs_data_1_14_sva_8_21_0_enexo_1 <= act_regs_data_and_196_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_102 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2632_enex5 ) begin
      reg_is_start_enexo_102 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_102 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2632_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_102 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_14_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_260_cse | act_regs_data_and_2632_enex5 ) begin
      reg_act_regs_data_0_14_sva_8_30_26_enexo <= act_regs_data_and_260_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_13_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2121_tmp | act_regs_data_and_2632_enex5 ) begin
      reg_act_regs_data_1_13_sva_dfm_2_30_26_enexo <= and_2121_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_102 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2632_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_102 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_13_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_200_cse | act_regs_data_and_2632_enex5 ) begin
      reg_act_regs_data_1_13_sva_8_30_26_enexo_1 <= act_regs_data_and_200_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_103 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2633_enex5 ) begin
      reg_is_start_enexo_103 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_13_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_1993_cse | act_regs_data_and_2633_enex5 ) begin
      reg_act_regs_data_1_13_sva_dfm_2_25_22_enexo <= and_1993_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_103 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2633_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_103 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_14_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_260_cse | act_regs_data_and_2633_enex5 ) begin
      reg_act_regs_data_0_14_sva_8_25_22_enexo <= act_regs_data_and_260_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_103 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2633_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_103 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_13_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_200_cse | act_regs_data_and_2633_enex5 ) begin
      reg_act_regs_data_1_13_sva_8_25_22_enexo_1 <= act_regs_data_and_200_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_104 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2634_enex5 ) begin
      reg_is_start_enexo_104 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_104 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2634_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_104 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_14_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_260_cse | act_regs_data_and_2634_enex5 ) begin
      reg_act_regs_data_0_14_sva_8_21_0_enexo <= act_regs_data_and_260_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_13_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_1993_cse | act_regs_data_and_2634_enex5 ) begin
      reg_act_regs_data_1_13_sva_dfm_2_21_0_enexo <= and_1993_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_104 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2634_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_104 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_13_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_200_cse | act_regs_data_and_2634_enex5 ) begin
      reg_act_regs_data_1_13_sva_8_21_0_enexo_1 <= act_regs_data_and_200_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_105 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2635_enex5 ) begin
      reg_is_start_enexo_105 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_105 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2635_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_105 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_13_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_264_cse | act_regs_data_and_2635_enex5 ) begin
      reg_act_regs_data_0_13_sva_8_30_26_enexo <= act_regs_data_and_264_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_12_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2119_tmp | act_regs_data_and_2635_enex5 ) begin
      reg_act_regs_data_1_12_sva_dfm_2_30_26_enexo <= and_2119_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_105 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2635_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_105 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_12_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_204_cse | act_regs_data_and_2635_enex5 ) begin
      reg_act_regs_data_1_12_sva_8_30_26_enexo_1 <= act_regs_data_and_204_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_106 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2636_enex5 ) begin
      reg_is_start_enexo_106 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_12_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_1991_cse | act_regs_data_and_2636_enex5 ) begin
      reg_act_regs_data_1_12_sva_dfm_2_25_22_enexo <= and_1991_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_106 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2636_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_106 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_13_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_264_cse | act_regs_data_and_2636_enex5 ) begin
      reg_act_regs_data_0_13_sva_8_25_22_enexo <= act_regs_data_and_264_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_106 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2636_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_106 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_12_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_204_cse | act_regs_data_and_2636_enex5 ) begin
      reg_act_regs_data_1_12_sva_8_25_22_enexo_1 <= act_regs_data_and_204_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_107 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2637_enex5 ) begin
      reg_is_start_enexo_107 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_107 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2637_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_107 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_13_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_264_cse | act_regs_data_and_2637_enex5 ) begin
      reg_act_regs_data_0_13_sva_8_21_0_enexo <= act_regs_data_and_264_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_12_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_1991_cse | act_regs_data_and_2637_enex5 ) begin
      reg_act_regs_data_1_12_sva_dfm_2_21_0_enexo <= and_1991_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_107 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2637_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_107 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_12_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_204_cse | act_regs_data_and_2637_enex5 ) begin
      reg_act_regs_data_1_12_sva_8_21_0_enexo_1 <= act_regs_data_and_204_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_108 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2638_enex5 ) begin
      reg_is_start_enexo_108 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_108 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2638_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_108 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_12_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_268_cse | act_regs_data_and_2638_enex5 ) begin
      reg_act_regs_data_0_12_sva_8_30_26_enexo <= act_regs_data_and_268_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_11_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2117_tmp | act_regs_data_and_2638_enex5 ) begin
      reg_act_regs_data_1_11_sva_dfm_2_30_26_enexo <= and_2117_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_108 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2638_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_108 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_11_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_208_cse | act_regs_data_and_2638_enex5 ) begin
      reg_act_regs_data_1_11_sva_8_30_26_enexo_1 <= act_regs_data_and_208_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_109 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2639_enex5 ) begin
      reg_is_start_enexo_109 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_11_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_1989_cse | act_regs_data_and_2639_enex5 ) begin
      reg_act_regs_data_1_11_sva_dfm_2_25_22_enexo <= and_1989_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_109 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2639_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_109 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_12_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_268_cse | act_regs_data_and_2639_enex5 ) begin
      reg_act_regs_data_0_12_sva_8_25_22_enexo <= act_regs_data_and_268_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_109 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2639_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_109 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_11_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_208_cse | act_regs_data_and_2639_enex5 ) begin
      reg_act_regs_data_1_11_sva_8_25_22_enexo_1 <= act_regs_data_and_208_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_110 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2640_enex5 ) begin
      reg_is_start_enexo_110 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_110 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2640_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_110 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_12_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_268_cse | act_regs_data_and_2640_enex5 ) begin
      reg_act_regs_data_0_12_sva_8_21_0_enexo <= act_regs_data_and_268_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_11_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_1989_cse | act_regs_data_and_2640_enex5 ) begin
      reg_act_regs_data_1_11_sva_dfm_2_21_0_enexo <= and_1989_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_110 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2640_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_110 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_11_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_208_cse | act_regs_data_and_2640_enex5 ) begin
      reg_act_regs_data_1_11_sva_8_21_0_enexo_1 <= act_regs_data_and_208_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_111 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2641_enex5 ) begin
      reg_is_start_enexo_111 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_111 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2641_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_111 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_11_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_272_cse | act_regs_data_and_2641_enex5 ) begin
      reg_act_regs_data_0_11_sva_8_30_26_enexo <= act_regs_data_and_272_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_10_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2115_tmp | act_regs_data_and_2641_enex5 ) begin
      reg_act_regs_data_1_10_sva_dfm_2_30_26_enexo <= and_2115_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_111 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2641_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_111 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_10_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_212_cse | act_regs_data_and_2641_enex5 ) begin
      reg_act_regs_data_1_10_sva_8_30_26_enexo_1 <= act_regs_data_and_212_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_112 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2642_enex5 ) begin
      reg_is_start_enexo_112 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_10_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_1987_cse | act_regs_data_and_2642_enex5 ) begin
      reg_act_regs_data_1_10_sva_dfm_2_25_22_enexo <= and_1987_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_112 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2642_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_112 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_11_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_272_cse | act_regs_data_and_2642_enex5 ) begin
      reg_act_regs_data_0_11_sva_8_25_22_enexo <= act_regs_data_and_272_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_112 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2642_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_112 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_10_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_212_cse | act_regs_data_and_2642_enex5 ) begin
      reg_act_regs_data_1_10_sva_8_25_22_enexo_1 <= act_regs_data_and_212_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_113 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2643_enex5 ) begin
      reg_is_start_enexo_113 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_113 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2643_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_113 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_11_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_272_cse | act_regs_data_and_2643_enex5 ) begin
      reg_act_regs_data_0_11_sva_8_21_0_enexo <= act_regs_data_and_272_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_10_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_1987_cse | act_regs_data_and_2643_enex5 ) begin
      reg_act_regs_data_1_10_sva_dfm_2_21_0_enexo <= and_1987_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_113 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2643_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_113 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_10_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_212_cse | act_regs_data_and_2643_enex5 ) begin
      reg_act_regs_data_1_10_sva_8_21_0_enexo_1 <= act_regs_data_and_212_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_114 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2644_enex5 ) begin
      reg_is_start_enexo_114 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_114 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2644_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_114 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_0_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_252_cse | act_regs_data_and_2644_enex5 ) begin
      reg_act_regs_data_1_0_sva_8_30_26_enexo <= act_regs_data_and_252_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_9_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2113_tmp | act_regs_data_and_2644_enex5 ) begin
      reg_act_regs_data_1_9_sva_dfm_2_30_26_enexo <= and_2113_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_114 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2644_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_114 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_9_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_216_cse | act_regs_data_and_2644_enex5 ) begin
      reg_act_regs_data_1_9_sva_8_30_26_enexo_1 <= act_regs_data_and_216_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_115 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2645_enex5 ) begin
      reg_is_start_enexo_115 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_9_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_1985_cse | act_regs_data_and_2645_enex5 ) begin
      reg_act_regs_data_1_9_sva_dfm_2_25_22_enexo <= and_1985_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_115 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2645_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_115 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_9_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_216_cse | act_regs_data_and_2645_enex5 ) begin
      reg_act_regs_data_1_9_sva_8_25_22_enexo_1 <= act_regs_data_and_216_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_0_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_252_cse | act_regs_data_and_2645_enex5 ) begin
      reg_act_regs_data_1_0_sva_8_25_22_enexo <= act_regs_data_and_252_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_115 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2645_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_115 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_116 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2646_enex5 ) begin
      reg_is_start_enexo_116 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_116 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2646_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_116 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_9_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_216_cse | act_regs_data_and_2646_enex5 ) begin
      reg_act_regs_data_1_9_sva_8_21_0_enexo_1 <= act_regs_data_and_216_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_0_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_252_cse | act_regs_data_and_2646_enex5 ) begin
      reg_act_regs_data_1_0_sva_8_21_0_enexo <= act_regs_data_and_252_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_9_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_1985_cse | act_regs_data_and_2646_enex5 ) begin
      reg_act_regs_data_1_9_sva_dfm_2_21_0_enexo <= and_1985_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_116 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2646_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_116 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_117 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2647_enex5 ) begin
      reg_is_start_enexo_117 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_117 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2647_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_117 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_8_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_220_cse | act_regs_data_and_2647_enex5 ) begin
      reg_act_regs_data_1_8_sva_8_30_26_enexo_1 <= act_regs_data_and_220_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_9_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_280_cse | act_regs_data_and_2647_enex5 ) begin
      reg_act_regs_data_0_9_sva_8_30_26_enexo <= act_regs_data_and_280_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_8_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2111_tmp | act_regs_data_and_2647_enex5 ) begin
      reg_act_regs_data_1_8_sva_dfm_2_30_26_enexo <= and_2111_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_117 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2647_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_117 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_118 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2648_enex5 ) begin
      reg_is_start_enexo_118 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_118 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2648_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_118 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_8_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_220_cse | act_regs_data_and_2648_enex5 ) begin
      reg_act_regs_data_1_8_sva_8_25_22_enexo_1 <= act_regs_data_and_220_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_9_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_280_cse | act_regs_data_and_2648_enex5 ) begin
      reg_act_regs_data_0_9_sva_8_25_22_enexo <= act_regs_data_and_280_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_8_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_1983_cse | act_regs_data_and_2648_enex5 ) begin
      reg_act_regs_data_1_8_sva_dfm_2_25_22_enexo <= and_1983_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_118 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2648_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_118 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_119 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2649_enex5 ) begin
      reg_is_start_enexo_119 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_119 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2649_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_119 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_8_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_220_cse | act_regs_data_and_2649_enex5 ) begin
      reg_act_regs_data_1_8_sva_8_21_0_enexo_1 <= act_regs_data_and_220_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_9_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_280_cse | act_regs_data_and_2649_enex5 ) begin
      reg_act_regs_data_0_9_sva_8_21_0_enexo <= act_regs_data_and_280_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_8_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_1983_cse | act_regs_data_and_2649_enex5 ) begin
      reg_act_regs_data_1_8_sva_dfm_2_21_0_enexo <= and_1983_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_119 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2649_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_119 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_120 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2650_enex5 ) begin
      reg_is_start_enexo_120 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_120 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2650_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_120 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_7_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_224_cse | act_regs_data_and_2650_enex5 ) begin
      reg_act_regs_data_1_7_sva_8_30_26_enexo_1 <= act_regs_data_and_224_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_8_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_284_cse | act_regs_data_and_2650_enex5 ) begin
      reg_act_regs_data_0_8_sva_8_30_26_enexo <= act_regs_data_and_284_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_7_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2109_tmp | act_regs_data_and_2650_enex5 ) begin
      reg_act_regs_data_1_7_sva_dfm_2_30_26_enexo <= and_2109_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_120 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2650_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_120 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_121 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2651_enex5 ) begin
      reg_is_start_enexo_121 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_121 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2651_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_121 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_7_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_224_cse | act_regs_data_and_2651_enex5 ) begin
      reg_act_regs_data_1_7_sva_8_25_22_enexo_1 <= act_regs_data_and_224_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_8_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_284_cse | act_regs_data_and_2651_enex5 ) begin
      reg_act_regs_data_0_8_sva_8_25_22_enexo <= act_regs_data_and_284_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_7_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_1981_cse | act_regs_data_and_2651_enex5 ) begin
      reg_act_regs_data_1_7_sva_dfm_2_25_22_enexo <= and_1981_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_121 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2651_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_121 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_122 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2652_enex5 ) begin
      reg_is_start_enexo_122 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_122 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2652_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_122 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_7_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_224_cse | act_regs_data_and_2652_enex5 ) begin
      reg_act_regs_data_1_7_sva_8_21_0_enexo_1 <= act_regs_data_and_224_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_8_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_284_cse | act_regs_data_and_2652_enex5 ) begin
      reg_act_regs_data_0_8_sva_8_21_0_enexo <= act_regs_data_and_284_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_7_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_1981_cse | act_regs_data_and_2652_enex5 ) begin
      reg_act_regs_data_1_7_sva_dfm_2_21_0_enexo <= and_1981_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_122 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2652_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_122 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_123 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2653_enex5 ) begin
      reg_is_start_enexo_123 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_123 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2653_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_123 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_6_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_228_cse | act_regs_data_and_2653_enex5 ) begin
      reg_act_regs_data_1_6_sva_8_30_26_enexo_1 <= act_regs_data_and_228_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_7_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_288_cse | act_regs_data_and_2653_enex5 ) begin
      reg_act_regs_data_0_7_sva_8_30_26_enexo <= act_regs_data_and_288_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_6_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2107_tmp | act_regs_data_and_2653_enex5 ) begin
      reg_act_regs_data_1_6_sva_dfm_2_30_26_enexo <= and_2107_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_123 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2653_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_123 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_124 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2654_enex5 ) begin
      reg_is_start_enexo_124 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_124 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2654_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_124 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_6_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_228_cse | act_regs_data_and_2654_enex5 ) begin
      reg_act_regs_data_1_6_sva_8_25_22_enexo_1 <= act_regs_data_and_228_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_7_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_288_cse | act_regs_data_and_2654_enex5 ) begin
      reg_act_regs_data_0_7_sva_8_25_22_enexo <= act_regs_data_and_288_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_6_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_1979_cse | act_regs_data_and_2654_enex5 ) begin
      reg_act_regs_data_1_6_sva_dfm_2_25_22_enexo <= and_1979_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_124 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2654_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_124 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_125 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2655_enex5 ) begin
      reg_is_start_enexo_125 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_125 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2655_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_125 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_6_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_228_cse | act_regs_data_and_2655_enex5 ) begin
      reg_act_regs_data_1_6_sva_8_21_0_enexo_1 <= act_regs_data_and_228_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_7_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_288_cse | act_regs_data_and_2655_enex5 ) begin
      reg_act_regs_data_0_7_sva_8_21_0_enexo <= act_regs_data_and_288_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_6_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_1979_cse | act_regs_data_and_2655_enex5 ) begin
      reg_act_regs_data_1_6_sva_dfm_2_21_0_enexo <= and_1979_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_125 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2655_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_125 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_126 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2656_enex5 ) begin
      reg_is_start_enexo_126 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_126 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2656_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_126 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_5_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_232_cse | act_regs_data_and_2656_enex5 ) begin
      reg_act_regs_data_1_5_sva_8_30_26_enexo_1 <= act_regs_data_and_232_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_6_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_292_cse | act_regs_data_and_2656_enex5 ) begin
      reg_act_regs_data_0_6_sva_8_30_26_enexo <= act_regs_data_and_292_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_5_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2105_tmp | act_regs_data_and_2656_enex5 ) begin
      reg_act_regs_data_1_5_sva_dfm_2_30_26_enexo <= and_2105_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_126 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2656_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_126 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_127 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2657_enex5 ) begin
      reg_is_start_enexo_127 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_127 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2657_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_127 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_5_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_232_cse | act_regs_data_and_2657_enex5 ) begin
      reg_act_regs_data_1_5_sva_8_25_22_enexo_1 <= act_regs_data_and_232_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_6_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_292_cse | act_regs_data_and_2657_enex5 ) begin
      reg_act_regs_data_0_6_sva_8_25_22_enexo <= act_regs_data_and_292_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_5_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_1977_cse | act_regs_data_and_2657_enex5 ) begin
      reg_act_regs_data_1_5_sva_dfm_2_25_22_enexo <= and_1977_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_127 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2657_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_127 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_128 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2658_enex5 ) begin
      reg_is_start_enexo_128 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_128 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2658_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_128 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_5_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_232_cse | act_regs_data_and_2658_enex5 ) begin
      reg_act_regs_data_1_5_sva_8_21_0_enexo_1 <= act_regs_data_and_232_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_6_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_292_cse | act_regs_data_and_2658_enex5 ) begin
      reg_act_regs_data_0_6_sva_8_21_0_enexo <= act_regs_data_and_292_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_5_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_1977_cse | act_regs_data_and_2658_enex5 ) begin
      reg_act_regs_data_1_5_sva_dfm_2_21_0_enexo <= and_1977_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_128 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2658_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_128 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_129 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2659_enex5 ) begin
      reg_is_start_enexo_129 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_129 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2659_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_129 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_4_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_236_cse | act_regs_data_and_2659_enex5 ) begin
      reg_act_regs_data_1_4_sva_8_30_26_enexo_1 <= act_regs_data_and_236_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_5_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_296_cse | act_regs_data_and_2659_enex5 ) begin
      reg_act_regs_data_0_5_sva_8_30_26_enexo <= act_regs_data_and_296_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_4_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2103_tmp | act_regs_data_and_2659_enex5 ) begin
      reg_act_regs_data_1_4_sva_dfm_2_30_26_enexo <= and_2103_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_129 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2659_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_129 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_130 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2660_enex5 ) begin
      reg_is_start_enexo_130 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_130 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2660_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_130 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_4_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_236_cse | act_regs_data_and_2660_enex5 ) begin
      reg_act_regs_data_1_4_sva_8_25_22_enexo_1 <= act_regs_data_and_236_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_5_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_296_cse | act_regs_data_and_2660_enex5 ) begin
      reg_act_regs_data_0_5_sva_8_25_22_enexo <= act_regs_data_and_296_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_4_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_1975_cse | act_regs_data_and_2660_enex5 ) begin
      reg_act_regs_data_1_4_sva_dfm_2_25_22_enexo <= and_1975_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_130 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2660_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_130 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_131 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2661_enex5 ) begin
      reg_is_start_enexo_131 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_131 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2661_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_131 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_4_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_236_cse | act_regs_data_and_2661_enex5 ) begin
      reg_act_regs_data_1_4_sva_8_21_0_enexo_1 <= act_regs_data_and_236_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_5_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_296_cse | act_regs_data_and_2661_enex5 ) begin
      reg_act_regs_data_0_5_sva_8_21_0_enexo <= act_regs_data_and_296_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_4_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_1975_cse | act_regs_data_and_2661_enex5 ) begin
      reg_act_regs_data_1_4_sva_dfm_2_21_0_enexo <= and_1975_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_131 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2661_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_131 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_132 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2662_enex5 ) begin
      reg_is_start_enexo_132 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_132 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2662_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_132 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_3_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_240_cse | act_regs_data_and_2662_enex5 ) begin
      reg_act_regs_data_1_3_sva_8_30_26_enexo_1 <= act_regs_data_and_240_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_4_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_300_cse | act_regs_data_and_2662_enex5 ) begin
      reg_act_regs_data_0_4_sva_8_30_26_enexo <= act_regs_data_and_300_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_3_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2101_tmp | act_regs_data_and_2662_enex5 ) begin
      reg_act_regs_data_1_3_sva_dfm_2_30_26_enexo <= and_2101_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_132 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2662_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_132 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_133 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2663_enex5 ) begin
      reg_is_start_enexo_133 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_4_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_300_cse | act_regs_data_and_2663_enex5 ) begin
      reg_act_regs_data_0_4_sva_8_25_22_enexo <= act_regs_data_and_300_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_133 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2663_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_133 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_3_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_240_cse | act_regs_data_and_2663_enex5 ) begin
      reg_act_regs_data_1_3_sva_8_25_22_enexo_1 <= act_regs_data_and_240_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_3_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_1973_cse | act_regs_data_and_2663_enex5 ) begin
      reg_act_regs_data_1_3_sva_dfm_2_25_22_enexo <= and_1973_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_133 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2663_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_133 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_134 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2664_enex5 ) begin
      reg_is_start_enexo_134 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_4_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_300_cse | act_regs_data_and_2664_enex5 ) begin
      reg_act_regs_data_0_4_sva_8_21_0_enexo <= act_regs_data_and_300_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_134 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2664_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_134 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_3_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_240_cse | act_regs_data_and_2664_enex5 ) begin
      reg_act_regs_data_1_3_sva_8_21_0_enexo_1 <= act_regs_data_and_240_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_3_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_1973_cse | act_regs_data_and_2664_enex5 ) begin
      reg_act_regs_data_1_3_sva_dfm_2_21_0_enexo <= and_1973_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_134 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2664_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_134 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_135 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2665_enex5 ) begin
      reg_is_start_enexo_135 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_3_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_304_cse | act_regs_data_and_2665_enex5 ) begin
      reg_act_regs_data_0_3_sva_8_30_26_enexo <= act_regs_data_and_304_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_135 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2665_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_135 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_2_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_244_cse | act_regs_data_and_2665_enex5 ) begin
      reg_act_regs_data_1_2_sva_8_30_26_enexo_1 <= act_regs_data_and_244_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_2_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2099_tmp | act_regs_data_and_2665_enex5 ) begin
      reg_act_regs_data_1_2_sva_dfm_2_30_26_enexo <= and_2099_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_135 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2665_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_135 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_136 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2666_enex5 ) begin
      reg_is_start_enexo_136 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_3_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_304_cse | act_regs_data_and_2666_enex5 ) begin
      reg_act_regs_data_0_3_sva_8_25_22_enexo <= act_regs_data_and_304_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_136 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2666_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_136 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_2_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_244_cse | act_regs_data_and_2666_enex5 ) begin
      reg_act_regs_data_1_2_sva_8_25_22_enexo_1 <= act_regs_data_and_244_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_2_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_1971_cse | act_regs_data_and_2666_enex5 ) begin
      reg_act_regs_data_1_2_sva_dfm_2_25_22_enexo <= and_1971_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_136 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2666_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_136 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_137 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2667_enex5 ) begin
      reg_is_start_enexo_137 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_3_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_304_cse | act_regs_data_and_2667_enex5 ) begin
      reg_act_regs_data_0_3_sva_8_21_0_enexo <= act_regs_data_and_304_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_137 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2667_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_137 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_2_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_244_cse | act_regs_data_and_2667_enex5 ) begin
      reg_act_regs_data_1_2_sva_8_21_0_enexo_1 <= act_regs_data_and_244_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_2_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_1971_cse | act_regs_data_and_2667_enex5 ) begin
      reg_act_regs_data_1_2_sva_dfm_2_21_0_enexo <= and_1971_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_137 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2667_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_137 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_138 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2668_enex5 ) begin
      reg_is_start_enexo_138 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_138 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2668_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_138 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_1_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_248_cse | act_regs_data_and_2668_enex5 ) begin
      reg_act_regs_data_1_1_sva_8_30_26_enexo_1 <= act_regs_data_and_248_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_10_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_276_cse | act_regs_data_and_2668_enex5 ) begin
      reg_act_regs_data_0_10_sva_8_30_26_enexo <= act_regs_data_and_276_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_1_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2097_tmp | act_regs_data_and_2668_enex5 ) begin
      reg_act_regs_data_1_1_sva_dfm_2_30_26_enexo <= and_2097_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_138 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2668_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_138 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_139 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2669_enex5 ) begin
      reg_is_start_enexo_139 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_139 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2669_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_139 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_1_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_248_cse | act_regs_data_and_2669_enex5 ) begin
      reg_act_regs_data_1_1_sva_8_25_22_enexo_1 <= act_regs_data_and_248_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_10_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_276_cse | act_regs_data_and_2669_enex5 ) begin
      reg_act_regs_data_0_10_sva_8_25_22_enexo <= act_regs_data_and_276_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_1_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_1969_cse | act_regs_data_and_2669_enex5 ) begin
      reg_act_regs_data_1_1_sva_dfm_2_25_22_enexo <= and_1969_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_139 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2669_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_139 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_140 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2670_enex5 ) begin
      reg_is_start_enexo_140 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_140 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2670_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_140 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_1_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_248_cse | act_regs_data_and_2670_enex5 ) begin
      reg_act_regs_data_1_1_sva_8_21_0_enexo_1 <= act_regs_data_and_248_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_10_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_276_cse | act_regs_data_and_2670_enex5 ) begin
      reg_act_regs_data_0_10_sva_8_21_0_enexo <= act_regs_data_and_276_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_1_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_1969_cse | act_regs_data_and_2670_enex5 ) begin
      reg_act_regs_data_1_1_sva_dfm_2_21_0_enexo <= and_1969_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_140 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2670_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_140 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_141 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2671_enex5 ) begin
      reg_is_start_enexo_141 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_1_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_312_cse | act_regs_data_and_2671_enex5 ) begin
      reg_act_regs_data_0_1_sva_8_30_26_enexo <= act_regs_data_and_312_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_141 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2671_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_141 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_0_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_252_cse | act_regs_data_and_2671_enex5 ) begin
      reg_act_regs_data_1_0_sva_8_30_26_enexo_1 <= act_regs_data_and_252_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_0_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2095_tmp | act_regs_data_and_2671_enex5 ) begin
      reg_act_regs_data_1_0_sva_dfm_2_30_26_enexo <= and_2095_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_141 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2671_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_141 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_142 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2672_enex5 ) begin
      reg_is_start_enexo_142 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_1_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_312_cse | act_regs_data_and_2672_enex5 ) begin
      reg_act_regs_data_0_1_sva_8_25_22_enexo <= act_regs_data_and_312_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_142 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2672_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_142 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_0_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_252_cse | act_regs_data_and_2672_enex5 ) begin
      reg_act_regs_data_1_0_sva_8_25_22_enexo_1 <= act_regs_data_and_252_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_0_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_1967_cse | act_regs_data_and_2672_enex5 ) begin
      reg_act_regs_data_1_0_sva_dfm_2_25_22_enexo <= and_1967_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_142 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2672_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_142 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_143 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2673_enex5 ) begin
      reg_is_start_enexo_143 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_1_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_312_cse | act_regs_data_and_2673_enex5 ) begin
      reg_act_regs_data_0_1_sva_8_21_0_enexo <= act_regs_data_and_312_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_143 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2673_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_143 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_0_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_252_cse | act_regs_data_and_2673_enex5 ) begin
      reg_act_regs_data_1_0_sva_8_21_0_enexo_1 <= act_regs_data_and_252_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_0_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_1967_cse | act_regs_data_and_2673_enex5 ) begin
      reg_act_regs_data_1_0_sva_dfm_2_21_0_enexo <= and_1967_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_143 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2673_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_143 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_144 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2674_enex5 ) begin
      reg_is_start_enexo_144 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_144 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2674_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_144 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_15_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_256_cse | act_regs_data_and_2674_enex5 ) begin
      reg_act_regs_data_0_15_sva_8_30_26_enexo_1 <= act_regs_data_and_256_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_1_30_26_enexo <=
          1'b1;
    end
    else if ( ActUnit_PushOutput_if_output_port_reg_data_data_and_22_cse | act_regs_data_and_2674_enex5
        ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_1_30_26_enexo <=
          ActUnit_PushOutput_if_output_port_reg_data_data_and_22_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_15_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2093_tmp | act_regs_data_and_2674_enex5 ) begin
      reg_act_regs_data_0_15_sva_dfm_2_30_26_enexo <= and_2093_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_144 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2674_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_144 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_145 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2675_enex5 ) begin
      reg_is_start_enexo_145 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_145 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2675_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_145 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_1_25_22_enexo <=
          1'b1;
    end
    else if ( and_1891_tmp | act_regs_data_and_2675_enex5 ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_1_25_22_enexo <=
          and_1891_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_15_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_256_cse | act_regs_data_and_2675_enex5 ) begin
      reg_act_regs_data_0_15_sva_8_25_22_enexo_1 <= act_regs_data_and_256_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_15_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_1965_cse | act_regs_data_and_2675_enex5 ) begin
      reg_act_regs_data_0_15_sva_dfm_2_25_22_enexo <= and_1965_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_145 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2675_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_145 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_146 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2676_enex5 ) begin
      reg_is_start_enexo_146 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_146 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2676_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_146 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_15_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_256_cse | act_regs_data_and_2676_enex5 ) begin
      reg_act_regs_data_0_15_sva_8_21_0_enexo_1 <= act_regs_data_and_256_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_15_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_1965_cse | act_regs_data_and_2676_enex5 ) begin
      reg_act_regs_data_0_15_sva_dfm_2_21_0_enexo <= and_1965_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Silu_for_3_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo
          <= 1'b1;
    end
    else if ( and_1867_tmp | act_regs_data_and_2676_enex5 ) begin
      reg_Silu_for_3_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo
          <= and_1867_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_146 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2676_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_146 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_147 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2677_enex5 ) begin
      reg_is_start_enexo_147 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_147 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2677_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_147 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_14_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_260_cse | act_regs_data_and_2677_enex5 ) begin
      reg_act_regs_data_0_14_sva_8_30_26_enexo_1 <= act_regs_data_and_260_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_1_30_26_enexo <=
          1'b1;
    end
    else if ( and_1933_tmp | act_regs_data_and_2677_enex5 ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_1_30_26_enexo <=
          and_1933_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_14_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2091_tmp | act_regs_data_and_2677_enex5 ) begin
      reg_act_regs_data_0_14_sva_dfm_2_30_26_enexo <= and_2091_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_147 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2677_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_147 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_148 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2678_enex5 ) begin
      reg_is_start_enexo_148 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_148 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2678_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_148 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_1_25_22_enexo <=
          1'b1;
    end
    else if ( and_1889_tmp | act_regs_data_and_2678_enex5 ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_1_25_22_enexo <=
          and_1889_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_14_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_260_cse | act_regs_data_and_2678_enex5 ) begin
      reg_act_regs_data_0_14_sva_8_25_22_enexo_1 <= act_regs_data_and_260_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_14_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_1963_cse | act_regs_data_and_2678_enex5 ) begin
      reg_act_regs_data_0_14_sva_dfm_2_25_22_enexo <= and_1963_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_148 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2678_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_148 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_149 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2679_enex5 ) begin
      reg_is_start_enexo_149 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Silu_for_2_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo
          <= 1'b1;
    end
    else if ( and_1865_tmp | act_regs_data_and_2679_enex5 ) begin
      reg_Silu_for_2_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo
          <= and_1865_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_149 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2679_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_149 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_14_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_260_cse | act_regs_data_and_2679_enex5 ) begin
      reg_act_regs_data_0_14_sva_8_21_0_enexo_1 <= act_regs_data_and_260_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_14_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_1963_cse | act_regs_data_and_2679_enex5 ) begin
      reg_act_regs_data_0_14_sva_dfm_2_21_0_enexo <= and_1963_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_149 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2679_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_149 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_150 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2680_enex5 ) begin
      reg_is_start_enexo_150 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_150 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2680_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_150 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_9_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_280_cse | act_regs_data_and_2680_enex5 ) begin
      reg_act_regs_data_0_9_sva_8_30_26_enexo_1 <= act_regs_data_and_280_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_0_sva_8_30_26_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_316_cse | act_regs_data_and_2680_enex5 ) begin
      reg_act_regs_data_0_0_sva_8_30_26_enexo <= act_regs_data_and_316_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_9_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2081_tmp | act_regs_data_and_2680_enex5 ) begin
      reg_act_regs_data_0_9_sva_dfm_2_30_26_enexo <= and_2081_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_150 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2680_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_150 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_151 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2681_enex5 ) begin
      reg_is_start_enexo_151 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_151 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2681_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_151 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_9_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_280_cse | act_regs_data_and_2681_enex5 ) begin
      reg_act_regs_data_0_9_sva_8_25_22_enexo_1 <= act_regs_data_and_280_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_0_sva_8_25_22_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_316_cse | act_regs_data_and_2681_enex5 ) begin
      reg_act_regs_data_0_0_sva_8_25_22_enexo <= act_regs_data_and_316_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_9_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_1953_cse | act_regs_data_and_2681_enex5 ) begin
      reg_act_regs_data_0_9_sva_dfm_2_25_22_enexo <= and_1953_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_151 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2681_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_151 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_152 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2682_enex5 ) begin
      reg_is_start_enexo_152 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_152 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2682_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_152 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_9_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_280_cse | act_regs_data_and_2682_enex5 ) begin
      reg_act_regs_data_0_9_sva_8_21_0_enexo_1 <= act_regs_data_and_280_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_0_sva_8_21_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_316_cse | act_regs_data_and_2682_enex5 ) begin
      reg_act_regs_data_0_0_sva_8_21_0_enexo <= act_regs_data_and_316_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_9_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_1953_cse | act_regs_data_and_2682_enex5 ) begin
      reg_act_regs_data_0_9_sva_dfm_2_21_0_enexo <= and_1953_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_152 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2682_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_152 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_153 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2683_enex5 ) begin
      reg_is_start_enexo_153 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_153 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2683_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_153 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_8_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_284_cse | act_regs_data_and_2683_enex5 ) begin
      reg_act_regs_data_0_8_sva_8_30_26_enexo_1 <= act_regs_data_and_284_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_8_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2079_tmp | act_regs_data_and_2683_enex5 ) begin
      reg_act_regs_data_0_8_sva_dfm_2_30_26_enexo <= and_2079_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_1_30_26_enexo <=
          1'b1;
    end
    else if ( ActUnit_PushOutput_if_output_port_reg_data_data_and_33_cse | act_regs_data_and_2683_enex5
        ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_1_30_26_enexo <=
          ActUnit_PushOutput_if_output_port_reg_data_data_and_33_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_153 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2683_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_153 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_154 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2684_enex5 ) begin
      reg_is_start_enexo_154 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_154 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2684_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_154 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_8_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_284_cse | act_regs_data_and_2684_enex5 ) begin
      reg_act_regs_data_0_8_sva_8_25_22_enexo_1 <= act_regs_data_and_284_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_8_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_1951_cse | act_regs_data_and_2684_enex5 ) begin
      reg_act_regs_data_0_8_sva_dfm_2_25_22_enexo <= and_1951_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_1_25_22_enexo <=
          1'b1;
    end
    else if ( ActUnit_PushOutput_if_output_port_reg_data_data_and_33_cse | act_regs_data_and_2684_enex5
        ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_1_25_22_enexo <=
          ActUnit_PushOutput_if_output_port_reg_data_data_and_33_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_154 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2684_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_154 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_155 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2685_enex5 ) begin
      reg_is_start_enexo_155 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_155 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2685_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_155 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Silu_for_y_8_sva_3_24_0_1_enexo <= 1'b1;
    end
    else if ( and_1877_tmp | act_regs_data_and_2685_enex5 ) begin
      reg_Silu_for_y_8_sva_3_24_0_1_enexo <= and_1877_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_8_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_284_cse | act_regs_data_and_2685_enex5 ) begin
      reg_act_regs_data_0_8_sva_8_21_0_enexo_1 <= act_regs_data_and_284_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_8_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_1951_cse | act_regs_data_and_2685_enex5 ) begin
      reg_act_regs_data_0_8_sva_dfm_2_21_0_enexo <= and_1951_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_155 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2685_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_155 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_156 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2686_enex5 ) begin
      reg_is_start_enexo_156 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_156 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2686_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_156 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_7_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_288_cse | act_regs_data_and_2686_enex5 ) begin
      reg_act_regs_data_0_7_sva_8_30_26_enexo_1 <= act_regs_data_and_288_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_7_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2077_tmp | act_regs_data_and_2686_enex5 ) begin
      reg_act_regs_data_0_7_sva_dfm_2_30_26_enexo <= and_2077_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_1_30_26_enexo <=
          1'b1;
    end
    else if ( ActUnit_PushOutput_if_output_port_reg_data_data_and_38_cse | act_regs_data_and_2686_enex5
        ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_1_30_26_enexo <=
          ActUnit_PushOutput_if_output_port_reg_data_data_and_38_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_156 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2686_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_156 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_157 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2687_enex5 ) begin
      reg_is_start_enexo_157 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_157 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2687_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_157 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_7_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_288_cse | act_regs_data_and_2687_enex5 ) begin
      reg_act_regs_data_0_7_sva_8_25_22_enexo_1 <= act_regs_data_and_288_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_7_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_1949_cse | act_regs_data_and_2687_enex5 ) begin
      reg_act_regs_data_0_7_sva_dfm_2_25_22_enexo <= and_1949_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_1_25_22_enexo <=
          1'b1;
    end
    else if ( and_1903_tmp | act_regs_data_and_2687_enex5 ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_1_25_22_enexo <=
          and_1903_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_157 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2687_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_157 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_158 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2688_enex5 ) begin
      reg_is_start_enexo_158 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Silu_for_y_1_sva_3_24_0_1_enexo <= 1'b1;
    end
    else if ( and_1864_tmp | act_regs_data_and_2688_enex5 ) begin
      reg_Silu_for_y_1_sva_3_24_0_1_enexo <= and_1864_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_158 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2688_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_158 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_7_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_288_cse | act_regs_data_and_2688_enex5 ) begin
      reg_act_regs_data_0_7_sva_8_21_0_enexo_1 <= act_regs_data_and_288_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_7_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_1949_cse | act_regs_data_and_2688_enex5 ) begin
      reg_act_regs_data_0_7_sva_dfm_2_21_0_enexo <= and_1949_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_158 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2688_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_158 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_159 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2689_enex5 ) begin
      reg_is_start_enexo_159 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_159 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2689_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_159 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_6_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_292_cse | act_regs_data_and_2689_enex5 ) begin
      reg_act_regs_data_0_6_sva_8_30_26_enexo_1 <= act_regs_data_and_292_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_6_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2075_tmp | act_regs_data_and_2689_enex5 ) begin
      reg_act_regs_data_0_6_sva_dfm_2_30_26_enexo <= and_2075_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_1_30_26_enexo <=
          1'b1;
    end
    else if ( ActUnit_PushOutput_if_output_port_reg_data_data_and_40_cse | act_regs_data_and_2689_enex5
        ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_1_30_26_enexo <=
          ActUnit_PushOutput_if_output_port_reg_data_data_and_40_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_159 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2689_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_159 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_160 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2690_enex5 ) begin
      reg_is_start_enexo_160 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_160 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2690_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_160 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_6_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_292_cse | act_regs_data_and_2690_enex5 ) begin
      reg_act_regs_data_0_6_sva_8_25_22_enexo_1 <= act_regs_data_and_292_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_6_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_1947_cse | act_regs_data_and_2690_enex5 ) begin
      reg_act_regs_data_0_6_sva_dfm_2_25_22_enexo <= and_1947_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_1_25_22_enexo <=
          1'b1;
    end
    else if ( and_1901_tmp | act_regs_data_and_2690_enex5 ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_1_25_22_enexo <=
          and_1901_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_160 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2690_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_160 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_161 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2691_enex5 ) begin
      reg_is_start_enexo_161 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_161 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2691_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_161 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Silu_for_9_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo
          <= 1'b1;
    end
    else if ( and_1879_tmp | act_regs_data_and_2691_enex5 ) begin
      reg_Silu_for_9_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo
          <= and_1879_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_6_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_292_cse | act_regs_data_and_2691_enex5 ) begin
      reg_act_regs_data_0_6_sva_8_21_0_enexo_1 <= act_regs_data_and_292_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_6_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_1947_cse | act_regs_data_and_2691_enex5 ) begin
      reg_act_regs_data_0_6_sva_dfm_2_21_0_enexo <= and_1947_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_161 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2691_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_161 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_162 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2692_enex5 ) begin
      reg_is_start_enexo_162 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_162 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2692_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_162 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_5_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_296_cse | act_regs_data_and_2692_enex5 ) begin
      reg_act_regs_data_0_5_sva_8_30_26_enexo_1 <= act_regs_data_and_296_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_5_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2073_tmp | act_regs_data_and_2692_enex5 ) begin
      reg_act_regs_data_0_5_sva_dfm_2_30_26_enexo <= and_2073_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_1_30_26_enexo <=
          1'b1;
    end
    else if ( ActUnit_PushOutput_if_output_port_reg_data_data_and_36_cse | act_regs_data_and_2692_enex5
        ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_1_30_26_enexo <=
          ActUnit_PushOutput_if_output_port_reg_data_data_and_36_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_162 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2692_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_162 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_163 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2693_enex5 ) begin
      reg_is_start_enexo_163 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_163 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2693_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_163 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_5_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_296_cse | act_regs_data_and_2693_enex5 ) begin
      reg_act_regs_data_0_5_sva_8_25_22_enexo_1 <= act_regs_data_and_296_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_5_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_1945_cse | act_regs_data_and_2693_enex5 ) begin
      reg_act_regs_data_0_5_sva_dfm_2_25_22_enexo <= and_1945_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_1_25_22_enexo <=
          1'b1;
    end
    else if ( and_1899_tmp | act_regs_data_and_2693_enex5 ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_1_25_22_enexo <=
          and_1899_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_163 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2693_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_163 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_164 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2694_enex5 ) begin
      reg_is_start_enexo_164 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_164 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2694_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_164 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Silu_for_7_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo
          <= 1'b1;
    end
    else if ( and_1875_tmp | act_regs_data_and_2694_enex5 ) begin
      reg_Silu_for_7_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo
          <= and_1875_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_5_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_296_cse | act_regs_data_and_2694_enex5 ) begin
      reg_act_regs_data_0_5_sva_8_21_0_enexo_1 <= act_regs_data_and_296_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_5_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_1945_cse | act_regs_data_and_2694_enex5 ) begin
      reg_act_regs_data_0_5_sva_dfm_2_21_0_enexo <= and_1945_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_164 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2694_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_164 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_165 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2695_enex5 ) begin
      reg_is_start_enexo_165 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_165 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2695_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_165 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_4_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_300_cse | act_regs_data_and_2695_enex5 ) begin
      reg_act_regs_data_0_4_sva_8_30_26_enexo_1 <= act_regs_data_and_300_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_4_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2071_tmp | act_regs_data_and_2695_enex5 ) begin
      reg_act_regs_data_0_4_sva_dfm_2_30_26_enexo <= and_2071_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_1_30_26_enexo <=
          1'b1;
    end
    else if ( ActUnit_PushOutput_if_output_port_reg_data_data_and_31_cse | act_regs_data_and_2695_enex5
        ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_1_30_26_enexo <=
          ActUnit_PushOutput_if_output_port_reg_data_data_and_31_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_165 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2695_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_165 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_166 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2696_enex5 ) begin
      reg_is_start_enexo_166 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_4_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_300_cse | act_regs_data_and_2696_enex5 ) begin
      reg_act_regs_data_0_4_sva_8_25_22_enexo_1 <= act_regs_data_and_300_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_166 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2696_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_166 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_1_25_22_enexo <=
          1'b1;
    end
    else if ( and_1897_tmp | act_regs_data_and_2696_enex5 ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_1_25_22_enexo <=
          and_1897_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_4_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_1943_cse | act_regs_data_and_2696_enex5 ) begin
      reg_act_regs_data_0_4_sva_dfm_2_25_22_enexo <= and_1943_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_166 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2696_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_166 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_167 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2697_enex5 ) begin
      reg_is_start_enexo_167 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_4_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_300_cse | act_regs_data_and_2697_enex5 ) begin
      reg_act_regs_data_0_4_sva_8_21_0_enexo_1 <= act_regs_data_and_300_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_167 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2697_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_167 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_4_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_1943_cse | act_regs_data_and_2697_enex5 ) begin
      reg_act_regs_data_0_4_sva_dfm_2_21_0_enexo <= and_1943_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Silu_for_6_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo
          <= 1'b1;
    end
    else if ( and_1873_tmp | act_regs_data_and_2697_enex5 ) begin
      reg_Silu_for_6_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo
          <= and_1873_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_167 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2697_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_167 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_168 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2698_enex5 ) begin
      reg_is_start_enexo_168 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_3_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_304_cse | act_regs_data_and_2698_enex5 ) begin
      reg_act_regs_data_0_3_sva_8_30_26_enexo_1 <= act_regs_data_and_304_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_168 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2698_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_168 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_3_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2069_tmp | act_regs_data_and_2698_enex5 ) begin
      reg_act_regs_data_0_3_sva_dfm_2_30_26_enexo <= and_2069_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_1_30_26_enexo <=
          1'b1;
    end
    else if ( ActUnit_PushOutput_if_output_port_reg_data_data_and_28_cse | act_regs_data_and_2698_enex5
        ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_1_30_26_enexo <=
          ActUnit_PushOutput_if_output_port_reg_data_data_and_28_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_168 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2698_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_168 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_169 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2699_enex5 ) begin
      reg_is_start_enexo_169 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_3_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_304_cse | act_regs_data_and_2699_enex5 ) begin
      reg_act_regs_data_0_3_sva_8_25_22_enexo_1 <= act_regs_data_and_304_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_169 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2699_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_169 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_1_25_22_enexo <=
          1'b1;
    end
    else if ( and_1895_tmp | act_regs_data_and_2699_enex5 ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_1_25_22_enexo <=
          and_1895_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_3_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_1941_cse | act_regs_data_and_2699_enex5 ) begin
      reg_act_regs_data_0_3_sva_dfm_2_25_22_enexo <= and_1941_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_169 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2699_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_169 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_170 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2700_enex5 ) begin
      reg_is_start_enexo_170 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_3_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_304_cse | act_regs_data_and_2700_enex5 ) begin
      reg_act_regs_data_0_3_sva_8_21_0_enexo_1 <= act_regs_data_and_304_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_170 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2700_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_170 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_3_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_1941_cse | act_regs_data_and_2700_enex5 ) begin
      reg_act_regs_data_0_3_sva_dfm_2_21_0_enexo <= and_1941_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Silu_for_5_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo
          <= 1'b1;
    end
    else if ( and_1871_tmp | act_regs_data_and_2700_enex5 ) begin
      reg_Silu_for_5_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo
          <= and_1871_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_170 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2700_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_170 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_171 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2701_enex5 ) begin
      reg_is_start_enexo_171 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_2_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_308_cse | act_regs_data_and_2701_enex5 ) begin
      reg_act_regs_data_0_2_sva_8_30_26_enexo_1 <= act_regs_data_and_308_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_171 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2701_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_171 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_1_30_26_enexo <=
          1'b1;
    end
    else if ( ActUnit_PushOutput_if_output_port_reg_data_data_and_25_cse | act_regs_data_and_2701_enex5
        ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_1_30_26_enexo <=
          ActUnit_PushOutput_if_output_port_reg_data_data_and_25_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_2_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2067_tmp | act_regs_data_and_2701_enex5 ) begin
      reg_act_regs_data_0_2_sva_dfm_2_30_26_enexo <= and_2067_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_171 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2701_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_171 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_172 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2702_enex5 ) begin
      reg_is_start_enexo_172 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_2_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_308_cse | act_regs_data_and_2702_enex5 ) begin
      reg_act_regs_data_0_2_sva_8_25_22_enexo_1 <= act_regs_data_and_308_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_172 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2702_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_172 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_1_25_22_enexo <=
          1'b1;
    end
    else if ( and_1893_tmp | act_regs_data_and_2702_enex5 ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_1_25_22_enexo <=
          and_1893_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_2_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_1939_cse | act_regs_data_and_2702_enex5 ) begin
      reg_act_regs_data_0_2_sva_dfm_2_25_22_enexo <= and_1939_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_172 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2702_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_172 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_173 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2703_enex5 ) begin
      reg_is_start_enexo_173 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_2_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_308_cse | act_regs_data_and_2703_enex5 ) begin
      reg_act_regs_data_0_2_sva_8_21_0_enexo_1 <= act_regs_data_and_308_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_173 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2703_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_173 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_2_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_1939_cse | act_regs_data_and_2703_enex5 ) begin
      reg_act_regs_data_0_2_sva_dfm_2_21_0_enexo <= and_1939_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Silu_for_4_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo
          <= 1'b1;
    end
    else if ( and_1869_tmp | act_regs_data_and_2703_enex5 ) begin
      reg_Silu_for_4_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo
          <= and_1869_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_173 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2703_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_173 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_15_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_mem_banks_read_read_data_and_16_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_15_enexo <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_14_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_mem_banks_read_read_data_and_17_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_14_enexo <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_13_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_mem_banks_read_read_data_and_18_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_13_enexo <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_12_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_mem_banks_read_read_data_and_19_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_12_enexo <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_11_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_mem_banks_read_read_data_and_20_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_11_enexo <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_10_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_mem_banks_read_read_data_and_21_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_10_enexo <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_9_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_mem_banks_read_read_data_and_22_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_9_enexo <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_8_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_mem_banks_read_read_data_and_23_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_8_enexo <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_7_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_mem_banks_read_read_data_and_24_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_7_enexo <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_6_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_mem_banks_read_read_data_and_25_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_6_enexo <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_5_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_mem_banks_read_read_data_and_26_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_5_enexo <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_4_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_mem_banks_read_read_data_and_27_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_4_enexo <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_3_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_mem_banks_read_read_data_and_28_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_3_enexo <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_2_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_mem_banks_read_read_data_and_29_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_2_enexo <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_1_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_mem_banks_read_read_data_and_30_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_1_enexo <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_mem_banks_read_read_data_and_31_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_enexo <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_15_enexo_1 <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_port_read_out_data_and_16_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_15_enexo_1 <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_write_req_valid_lpi_1_dfm_5_enexo <= 1'b1;
    end
    else if ( ActUnitRun_wen | act_port_read_out_data_and_16_enex5 ) begin
      reg_act_write_req_valid_lpi_1_dfm_5_enexo <= ActUnitRun_wen;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_31_0_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_read_data_and_16_enex5 | act_port_read_out_data_and_16_enex5
        ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_31_0_enexo <= act_mem_banks_read_read_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_63_32_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_read_data_and_17_enex5 | act_port_read_out_data_and_17_enex5
        ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_63_32_enexo <= act_mem_banks_read_read_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_write_req_valid_lpi_1_dfm_5_enexo_1 <= 1'b1;
    end
    else if ( ActUnitRun_wen | act_port_read_out_data_and_17_enex5 ) begin
      reg_act_write_req_valid_lpi_1_dfm_5_enexo_1 <= ActUnitRun_wen;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_14_enexo_1 <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_port_read_out_data_and_17_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_14_enexo_1 <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_write_req_valid_lpi_1_dfm_5_enexo_2 <= 1'b1;
    end
    else if ( ActUnitRun_wen | act_port_read_out_data_and_18_enex5 ) begin
      reg_act_write_req_valid_lpi_1_dfm_5_enexo_2 <= ActUnitRun_wen;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_13_enexo_1 <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_port_read_out_data_and_18_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_13_enexo_1 <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_95_64_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_read_data_and_18_enex5 | act_port_read_out_data_and_18_enex5
        ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_95_64_enexo <= act_mem_banks_read_read_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_write_req_valid_lpi_1_dfm_5_enexo_3 <= 1'b1;
    end
    else if ( ActUnitRun_wen | act_port_read_out_data_and_19_enex5 ) begin
      reg_act_write_req_valid_lpi_1_dfm_5_enexo_3 <= ActUnitRun_wen;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_12_enexo_1 <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_port_read_out_data_and_19_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_12_enexo_1 <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_127_96_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_read_data_and_19_enex5 | act_port_read_out_data_and_19_enex5
        ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_127_96_enexo <= act_mem_banks_read_read_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_11_enexo_1 <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_port_read_out_data_and_20_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_11_enexo_1 <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_write_req_valid_lpi_1_dfm_5_enexo_4 <= 1'b1;
    end
    else if ( ActUnitRun_wen | act_port_read_out_data_and_20_enex5 ) begin
      reg_act_write_req_valid_lpi_1_dfm_5_enexo_4 <= ActUnitRun_wen;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_159_128_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_read_data_and_20_enex5 | act_port_read_out_data_and_20_enex5
        ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_159_128_enexo <= act_mem_banks_read_read_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_191_160_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_read_data_and_21_enex5 | act_port_read_out_data_and_21_enex5
        ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_191_160_enexo <= act_mem_banks_read_read_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_10_enexo_1 <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_port_read_out_data_and_21_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_10_enexo_1 <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_write_req_valid_lpi_1_dfm_5_enexo_5 <= 1'b1;
    end
    else if ( ActUnitRun_wen | act_port_read_out_data_and_21_enex5 ) begin
      reg_act_write_req_valid_lpi_1_dfm_5_enexo_5 <= ActUnitRun_wen;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_9_enexo_1 <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_port_read_out_data_and_22_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_9_enexo_1 <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_write_req_valid_lpi_1_dfm_5_enexo_6 <= 1'b1;
    end
    else if ( ActUnitRun_wen | act_port_read_out_data_and_22_enex5 ) begin
      reg_act_write_req_valid_lpi_1_dfm_5_enexo_6 <= ActUnitRun_wen;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_223_192_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_read_data_and_22_enex5 | act_port_read_out_data_and_22_enex5
        ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_223_192_enexo <= act_mem_banks_read_read_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_255_224_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_read_data_and_23_enex5 | act_port_read_out_data_and_23_enex5
        ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_255_224_enexo <= act_mem_banks_read_read_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_8_enexo_1 <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_port_read_out_data_and_23_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_8_enexo_1 <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_write_req_valid_lpi_1_dfm_5_enexo_7 <= 1'b1;
    end
    else if ( ActUnitRun_wen | act_port_read_out_data_and_23_enex5 ) begin
      reg_act_write_req_valid_lpi_1_dfm_5_enexo_7 <= ActUnitRun_wen;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_287_256_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_read_data_and_24_enex5 | act_port_read_out_data_and_24_enex5
        ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_287_256_enexo <= act_mem_banks_read_read_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_7_enexo_1 <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_port_read_out_data_and_24_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_7_enexo_1 <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_write_req_valid_lpi_1_dfm_5_enexo_8 <= 1'b1;
    end
    else if ( ActUnitRun_wen | act_port_read_out_data_and_24_enex5 ) begin
      reg_act_write_req_valid_lpi_1_dfm_5_enexo_8 <= ActUnitRun_wen;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_319_288_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_read_data_and_25_enex5 | act_port_read_out_data_and_25_enex5
        ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_319_288_enexo <= act_mem_banks_read_read_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_6_enexo_1 <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_port_read_out_data_and_25_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_6_enexo_1 <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_write_req_valid_lpi_1_dfm_5_enexo_9 <= 1'b1;
    end
    else if ( ActUnitRun_wen | act_port_read_out_data_and_25_enex5 ) begin
      reg_act_write_req_valid_lpi_1_dfm_5_enexo_9 <= ActUnitRun_wen;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_351_320_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_read_data_and_26_enex5 | act_port_read_out_data_and_26_enex5
        ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_351_320_enexo <= act_mem_banks_read_read_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_write_req_valid_lpi_1_dfm_5_enexo_10 <= 1'b1;
    end
    else if ( ActUnitRun_wen | act_port_read_out_data_and_26_enex5 ) begin
      reg_act_write_req_valid_lpi_1_dfm_5_enexo_10 <= ActUnitRun_wen;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_5_enexo_1 <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_port_read_out_data_and_26_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_5_enexo_1 <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_383_352_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_read_data_and_27_enex5 | act_port_read_out_data_and_27_enex5
        ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_383_352_enexo <= act_mem_banks_read_read_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_write_req_valid_lpi_1_dfm_5_enexo_11 <= 1'b1;
    end
    else if ( ActUnitRun_wen | act_port_read_out_data_and_27_enex5 ) begin
      reg_act_write_req_valid_lpi_1_dfm_5_enexo_11 <= ActUnitRun_wen;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_4_enexo_1 <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_port_read_out_data_and_27_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_4_enexo_1 <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_415_384_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_read_data_and_28_enex5 | act_port_read_out_data_and_28_enex5
        ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_415_384_enexo <= act_mem_banks_read_read_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_write_req_valid_lpi_1_dfm_5_enexo_12 <= 1'b1;
    end
    else if ( ActUnitRun_wen | act_port_read_out_data_and_28_enex5 ) begin
      reg_act_write_req_valid_lpi_1_dfm_5_enexo_12 <= ActUnitRun_wen;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_3_enexo_1 <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_port_read_out_data_and_28_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_3_enexo_1 <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_2_enexo_1 <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_port_read_out_data_and_29_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_2_enexo_1 <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_write_req_valid_lpi_1_dfm_5_enexo_13 <= 1'b1;
    end
    else if ( ActUnitRun_wen | act_port_read_out_data_and_29_enex5 ) begin
      reg_act_write_req_valid_lpi_1_dfm_5_enexo_13 <= ActUnitRun_wen;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_447_416_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_read_data_and_29_enex5 | act_port_read_out_data_and_29_enex5
        ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_447_416_enexo <= act_mem_banks_read_read_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_1_enexo_1 <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_port_read_out_data_and_30_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_1_enexo_1 <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_479_448_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_read_data_and_30_enex5 | act_port_read_out_data_and_30_enex5
        ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_479_448_enexo <= act_mem_banks_read_read_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_write_req_valid_lpi_1_dfm_5_enexo_14 <= 1'b1;
    end
    else if ( ActUnitRun_wen | act_port_read_out_data_and_30_enex5 ) begin
      reg_act_write_req_valid_lpi_1_dfm_5_enexo_14 <= ActUnitRun_wen;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_for_mux_enexo_1 <= 1'b1;
    end
    else if ( act_mem_banks_read_for_and_cse | act_port_read_out_data_and_31_enex5
        ) begin
      reg_act_mem_banks_read_for_mux_enexo_1 <= act_mem_banks_read_for_and_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_511_480_enexo <= 1'b1;
    end
    else if ( act_mem_banks_read_read_data_and_31_enex5 | act_port_read_out_data_and_31_enex5
        ) begin
      reg_act_mem_banks_read_read_data_lpi_1_dfm_1_511_480_enexo <= act_mem_banks_read_read_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_write_req_valid_lpi_1_dfm_5_enexo_15 <= 1'b1;
    end
    else if ( ActUnitRun_wen | act_port_read_out_data_and_31_enex5 ) begin
      reg_act_write_req_valid_lpi_1_dfm_5_enexo_15 <= ActUnitRun_wen;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_37_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_37_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_37_enex5
        ) begin
      reg_act_config_inst_counter_enexo <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_15_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2674_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_37_enex5
        ) begin
      reg_act_regs_data_0_15_1_enexo <= act_regs_data_and_2674_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_15_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2626_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_37_enex5
        ) begin
      reg_act_regs_data_1_15_1_enexo <= act_regs_data_and_2626_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_15_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2578_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_37_enex5
        ) begin
      reg_act_regs_data_2_15_1_enexo <= act_regs_data_and_2578_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_15_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2530_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_37_enex5
        ) begin
      reg_act_regs_data_3_15_1_enexo <= act_regs_data_and_2530_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_1 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_38_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_1 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_1 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_38_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_1 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_1 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_38_enex5
        ) begin
      reg_act_config_inst_counter_enexo_1 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_15_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2531_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_38_enex5
        ) begin
      reg_act_regs_data_3_15_2_enexo <= act_regs_data_and_2531_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_15_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2579_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_38_enex5
        ) begin
      reg_act_regs_data_2_15_2_enexo <= act_regs_data_and_2579_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_15_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2675_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_38_enex5
        ) begin
      reg_act_regs_data_0_15_2_enexo <= act_regs_data_and_2675_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_15_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2627_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_38_enex5
        ) begin
      reg_act_regs_data_1_15_2_enexo <= act_regs_data_and_2627_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_2 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_39_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_2 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_2 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_39_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_2 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_15_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2580_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_39_enex5
        ) begin
      reg_act_regs_data_2_15_3_enexo <= act_regs_data_and_2580_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_2 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_39_enex5
        ) begin
      reg_act_config_inst_counter_enexo_2 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_15_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2676_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_39_enex5
        ) begin
      reg_act_regs_data_0_15_3_enexo <= act_regs_data_and_2676_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_15_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2628_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_39_enex5
        ) begin
      reg_act_regs_data_1_15_3_enexo <= act_regs_data_and_2628_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_15_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2532_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_39_enex5
        ) begin
      reg_act_regs_data_3_15_3_enexo <= act_regs_data_and_2532_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_3 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_40_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_3 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_14_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2629_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_40_enex5
        ) begin
      reg_act_regs_data_1_14_1_enexo <= act_regs_data_and_2629_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_3 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_40_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_3 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_3 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_40_enex5
        ) begin
      reg_act_config_inst_counter_enexo_3 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_14_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2581_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_40_enex5
        ) begin
      reg_act_regs_data_2_14_1_enexo <= act_regs_data_and_2581_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_14_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2533_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_40_enex5
        ) begin
      reg_act_regs_data_3_14_1_enexo <= act_regs_data_and_2533_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_14_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2677_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_40_enex5
        ) begin
      reg_act_regs_data_0_14_1_enexo <= act_regs_data_and_2677_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_4 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_41_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_4 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_14_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2678_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_41_enex5
        ) begin
      reg_act_regs_data_0_14_2_enexo <= act_regs_data_and_2678_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_4 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_41_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_4 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_4 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_41_enex5
        ) begin
      reg_act_config_inst_counter_enexo_4 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_14_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2582_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_41_enex5
        ) begin
      reg_act_regs_data_2_14_2_enexo <= act_regs_data_and_2582_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_14_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2534_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_41_enex5
        ) begin
      reg_act_regs_data_3_14_2_enexo <= act_regs_data_and_2534_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_14_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2630_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_41_enex5
        ) begin
      reg_act_regs_data_1_14_2_enexo <= act_regs_data_and_2630_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_5 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_42_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_5 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_5 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_42_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_5 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_5 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_42_enex5
        ) begin
      reg_act_config_inst_counter_enexo_5 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_14_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2679_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_42_enex5
        ) begin
      reg_act_regs_data_0_14_3_enexo <= act_regs_data_and_2679_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_14_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2583_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_42_enex5
        ) begin
      reg_act_regs_data_2_14_3_enexo <= act_regs_data_and_2583_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_14_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2535_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_42_enex5
        ) begin
      reg_act_regs_data_3_14_3_enexo <= act_regs_data_and_2535_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_14_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2631_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_42_enex5
        ) begin
      reg_act_regs_data_1_14_3_enexo <= act_regs_data_and_2631_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_6 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_43_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_6 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_13_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2632_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_43_enex5
        ) begin
      reg_act_regs_data_1_13_1_enexo <= act_regs_data_and_2632_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_13_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2584_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_43_enex5
        ) begin
      reg_act_regs_data_2_13_1_enexo <= act_regs_data_and_2584_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_6 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_43_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_6 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_6 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_43_enex5
        ) begin
      reg_act_config_inst_counter_enexo_6 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_13_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2749_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_43_enex5
        ) begin
      reg_act_regs_data_0_13_1_enexo <= act_regs_data_and_2749_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_13_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2536_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_43_enex5
        ) begin
      reg_act_regs_data_3_13_1_enexo <= act_regs_data_and_2536_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_13_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2537_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_44_enex5
        ) begin
      reg_act_regs_data_3_13_2_enexo <= act_regs_data_and_2537_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_7 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_44_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_7 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_7 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_44_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_7 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_13_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2750_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_44_enex5
        ) begin
      reg_act_regs_data_0_13_2_enexo <= act_regs_data_and_2750_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_7 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_44_enex5
        ) begin
      reg_act_config_inst_counter_enexo_7 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_13_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2633_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_44_enex5
        ) begin
      reg_act_regs_data_1_13_2_enexo <= act_regs_data_and_2633_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_13_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2585_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_44_enex5
        ) begin
      reg_act_regs_data_2_13_2_enexo <= act_regs_data_and_2585_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_8 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_45_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_8 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_8 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_45_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_8 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_8 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_45_enex5
        ) begin
      reg_act_config_inst_counter_enexo_8 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_13_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2586_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_45_enex5
        ) begin
      reg_act_regs_data_2_13_3_enexo <= act_regs_data_and_2586_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_13_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2538_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_45_enex5
        ) begin
      reg_act_regs_data_3_13_3_enexo <= act_regs_data_and_2538_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_13_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2634_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_45_enex5
        ) begin
      reg_act_regs_data_1_13_3_enexo <= act_regs_data_and_2634_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_13_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2751_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_45_enex5
        ) begin
      reg_act_regs_data_0_13_3_enexo <= act_regs_data_and_2751_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_9 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_46_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_9 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_9 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_46_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_9 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_9 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_46_enex5
        ) begin
      reg_act_config_inst_counter_enexo_9 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_12_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2587_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_46_enex5
        ) begin
      reg_act_regs_data_2_12_1_enexo <= act_regs_data_and_2587_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_12_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2752_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_46_enex5
        ) begin
      reg_act_regs_data_0_12_1_enexo <= act_regs_data_and_2752_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_12_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2635_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_46_enex5
        ) begin
      reg_act_regs_data_1_12_1_enexo <= act_regs_data_and_2635_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_12_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2539_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_46_enex5
        ) begin
      reg_act_regs_data_3_12_1_enexo <= act_regs_data_and_2539_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_10 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_47_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_10 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_10 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_47_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_10 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_12_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2588_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_47_enex5
        ) begin
      reg_act_regs_data_2_12_2_enexo <= act_regs_data_and_2588_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_10 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_47_enex5
        ) begin
      reg_act_config_inst_counter_enexo_10 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_12_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2753_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_47_enex5
        ) begin
      reg_act_regs_data_0_12_2_enexo <= act_regs_data_and_2753_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_12_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2540_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_47_enex5
        ) begin
      reg_act_regs_data_3_12_2_enexo <= act_regs_data_and_2540_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_12_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2636_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_47_enex5
        ) begin
      reg_act_regs_data_1_12_2_enexo <= act_regs_data_and_2636_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_11 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_48_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_11 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_11 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_48_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_11 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_11 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_48_enex5
        ) begin
      reg_act_config_inst_counter_enexo_11 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_12_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2754_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_48_enex5
        ) begin
      reg_act_regs_data_0_12_3_enexo <= act_regs_data_and_2754_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_12_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2589_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_48_enex5
        ) begin
      reg_act_regs_data_2_12_3_enexo <= act_regs_data_and_2589_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_12_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2541_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_48_enex5
        ) begin
      reg_act_regs_data_3_12_3_enexo <= act_regs_data_and_2541_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_12_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2637_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_48_enex5
        ) begin
      reg_act_regs_data_1_12_3_enexo <= act_regs_data_and_2637_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_12 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_49_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_12 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_12 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_49_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_12 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_12 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_49_enex5
        ) begin
      reg_act_config_inst_counter_enexo_12 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_11_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2590_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_49_enex5
        ) begin
      reg_act_regs_data_2_11_1_enexo <= act_regs_data_and_2590_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_11_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2542_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_49_enex5
        ) begin
      reg_act_regs_data_3_11_1_enexo <= act_regs_data_and_2542_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_11_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2755_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_49_enex5
        ) begin
      reg_act_regs_data_0_11_1_enexo <= act_regs_data_and_2755_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_11_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2638_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_49_enex5
        ) begin
      reg_act_regs_data_1_11_1_enexo <= act_regs_data_and_2638_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_13 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_50_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_13 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_13 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_50_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_13 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_13 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_50_enex5
        ) begin
      reg_act_config_inst_counter_enexo_13 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_11_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2591_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_50_enex5
        ) begin
      reg_act_regs_data_2_11_2_enexo <= act_regs_data_and_2591_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_11_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2756_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_50_enex5
        ) begin
      reg_act_regs_data_0_11_2_enexo <= act_regs_data_and_2756_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_11_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2543_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_50_enex5
        ) begin
      reg_act_regs_data_3_11_2_enexo <= act_regs_data_and_2543_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_11_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2639_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_50_enex5
        ) begin
      reg_act_regs_data_1_11_2_enexo <= act_regs_data_and_2639_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_14 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_51_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_14 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_14 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_51_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_14 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_14 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_51_enex5
        ) begin
      reg_act_config_inst_counter_enexo_14 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_11_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2757_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_51_enex5
        ) begin
      reg_act_regs_data_0_11_3_enexo <= act_regs_data_and_2757_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_11_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2640_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_51_enex5
        ) begin
      reg_act_regs_data_1_11_3_enexo <= act_regs_data_and_2640_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_11_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2592_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_51_enex5
        ) begin
      reg_act_regs_data_2_11_3_enexo <= act_regs_data_and_2592_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_11_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2544_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_51_enex5
        ) begin
      reg_act_regs_data_3_11_3_enexo <= act_regs_data_and_2544_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_15 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_52_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_15 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_15 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_52_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_15 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_15 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_52_enex5
        ) begin
      reg_act_config_inst_counter_enexo_15 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_10_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2641_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_52_enex5
        ) begin
      reg_act_regs_data_1_10_1_enexo <= act_regs_data_and_2641_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_10_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2593_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_52_enex5
        ) begin
      reg_act_regs_data_2_10_1_enexo <= act_regs_data_and_2593_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_10_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2545_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_52_enex5
        ) begin
      reg_act_regs_data_3_10_1_enexo <= act_regs_data_and_2545_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_10_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2758_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_52_enex5
        ) begin
      reg_act_regs_data_0_10_1_enexo <= act_regs_data_and_2758_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_16 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_53_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_16 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_16 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_53_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_16 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_16 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_53_enex5
        ) begin
      reg_act_config_inst_counter_enexo_16 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_10_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2642_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_53_enex5
        ) begin
      reg_act_regs_data_1_10_2_enexo <= act_regs_data_and_2642_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_10_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2759_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_53_enex5
        ) begin
      reg_act_regs_data_0_10_2_enexo <= act_regs_data_and_2759_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_10_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2546_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_53_enex5
        ) begin
      reg_act_regs_data_3_10_2_enexo <= act_regs_data_and_2546_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_10_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2594_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_53_enex5
        ) begin
      reg_act_regs_data_2_10_2_enexo <= act_regs_data_and_2594_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_17 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_54_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_17 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_17 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_54_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_17 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_17 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_54_enex5
        ) begin
      reg_act_config_inst_counter_enexo_17 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_10_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2547_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_54_enex5
        ) begin
      reg_act_regs_data_3_10_3_enexo <= act_regs_data_and_2547_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_10_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2760_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_54_enex5
        ) begin
      reg_act_regs_data_0_10_3_enexo <= act_regs_data_and_2760_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_10_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2595_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_54_enex5
        ) begin
      reg_act_regs_data_2_10_3_enexo <= act_regs_data_and_2595_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_10_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2643_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_54_enex5
        ) begin
      reg_act_regs_data_1_10_3_enexo <= act_regs_data_and_2643_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_18 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_55_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_18 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_18 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_55_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_18 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_18 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_55_enex5
        ) begin
      reg_act_config_inst_counter_enexo_18 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_9_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2644_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_55_enex5
        ) begin
      reg_act_regs_data_1_9_1_enexo <= act_regs_data_and_2644_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_9_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2548_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_55_enex5
        ) begin
      reg_act_regs_data_3_9_1_enexo <= act_regs_data_and_2548_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_9_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2680_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_55_enex5
        ) begin
      reg_act_regs_data_0_9_1_enexo <= act_regs_data_and_2680_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_9_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2596_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_55_enex5
        ) begin
      reg_act_regs_data_2_9_1_enexo <= act_regs_data_and_2596_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_19 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_56_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_19 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_19 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_56_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_19 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_19 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_56_enex5
        ) begin
      reg_act_config_inst_counter_enexo_19 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_9_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2681_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_56_enex5
        ) begin
      reg_act_regs_data_0_9_2_enexo <= act_regs_data_and_2681_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_9_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2597_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_56_enex5
        ) begin
      reg_act_regs_data_2_9_2_enexo <= act_regs_data_and_2597_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_9_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2645_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_56_enex5
        ) begin
      reg_act_regs_data_1_9_2_enexo <= act_regs_data_and_2645_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_9_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2549_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_56_enex5
        ) begin
      reg_act_regs_data_3_9_2_enexo <= act_regs_data_and_2549_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_20 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_57_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_20 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_20 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_57_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_20 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_20 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_57_enex5
        ) begin
      reg_act_config_inst_counter_enexo_20 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_9_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2646_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_57_enex5
        ) begin
      reg_act_regs_data_1_9_3_enexo <= act_regs_data_and_2646_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_9_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2682_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_57_enex5
        ) begin
      reg_act_regs_data_0_9_3_enexo <= act_regs_data_and_2682_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_9_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2598_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_57_enex5
        ) begin
      reg_act_regs_data_2_9_3_enexo <= act_regs_data_and_2598_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_9_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2550_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_57_enex5
        ) begin
      reg_act_regs_data_3_9_3_enexo <= act_regs_data_and_2550_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_21 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_58_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_21 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_21 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_58_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_21 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_21 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_58_enex5
        ) begin
      reg_act_config_inst_counter_enexo_21 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_8_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2599_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_58_enex5
        ) begin
      reg_act_regs_data_2_8_1_enexo <= act_regs_data_and_2599_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_8_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2683_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_58_enex5
        ) begin
      reg_act_regs_data_0_8_1_enexo <= act_regs_data_and_2683_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_8_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2551_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_58_enex5
        ) begin
      reg_act_regs_data_3_8_1_enexo <= act_regs_data_and_2551_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_8_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2647_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_58_enex5
        ) begin
      reg_act_regs_data_1_8_1_enexo <= act_regs_data_and_2647_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_22 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_59_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_22 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_22 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_59_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_22 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_22 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_59_enex5
        ) begin
      reg_act_config_inst_counter_enexo_22 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_8_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2684_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_59_enex5
        ) begin
      reg_act_regs_data_0_8_2_enexo <= act_regs_data_and_2684_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_8_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2648_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_59_enex5
        ) begin
      reg_act_regs_data_1_8_2_enexo <= act_regs_data_and_2648_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_8_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2600_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_59_enex5
        ) begin
      reg_act_regs_data_2_8_2_enexo <= act_regs_data_and_2600_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_8_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2552_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_59_enex5
        ) begin
      reg_act_regs_data_3_8_2_enexo <= act_regs_data_and_2552_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_23 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_60_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_23 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_23 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_60_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_23 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_23 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_60_enex5
        ) begin
      reg_act_config_inst_counter_enexo_23 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_8_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2685_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_60_enex5
        ) begin
      reg_act_regs_data_0_8_3_enexo <= act_regs_data_and_2685_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_8_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2601_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_60_enex5
        ) begin
      reg_act_regs_data_2_8_3_enexo <= act_regs_data_and_2601_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_8_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2649_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_60_enex5
        ) begin
      reg_act_regs_data_1_8_3_enexo <= act_regs_data_and_2649_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_8_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2553_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_60_enex5
        ) begin
      reg_act_regs_data_3_8_3_enexo <= act_regs_data_and_2553_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_24 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_61_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_24 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_24 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_61_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_24 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_24 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_61_enex5
        ) begin
      reg_act_config_inst_counter_enexo_24 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_7_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2554_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_61_enex5
        ) begin
      reg_act_regs_data_3_7_1_enexo <= act_regs_data_and_2554_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_7_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2650_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_61_enex5
        ) begin
      reg_act_regs_data_1_7_1_enexo <= act_regs_data_and_2650_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_7_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2686_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_61_enex5
        ) begin
      reg_act_regs_data_0_7_1_enexo <= act_regs_data_and_2686_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_7_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2602_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_61_enex5
        ) begin
      reg_act_regs_data_2_7_1_enexo <= act_regs_data_and_2602_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_25 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_62_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_25 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_25 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_62_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_25 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_25 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_62_enex5
        ) begin
      reg_act_config_inst_counter_enexo_25 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_7_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2687_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_62_enex5
        ) begin
      reg_act_regs_data_0_7_2_enexo <= act_regs_data_and_2687_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_7_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2603_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_62_enex5
        ) begin
      reg_act_regs_data_2_7_2_enexo <= act_regs_data_and_2603_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_7_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2555_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_62_enex5
        ) begin
      reg_act_regs_data_3_7_2_enexo <= act_regs_data_and_2555_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_7_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2651_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_62_enex5
        ) begin
      reg_act_regs_data_1_7_2_enexo <= act_regs_data_and_2651_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_26 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_63_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_26 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_26 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_63_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_26 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_26 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_63_enex5
        ) begin
      reg_act_config_inst_counter_enexo_26 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_7_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2688_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_63_enex5
        ) begin
      reg_act_regs_data_0_7_3_enexo <= act_regs_data_and_2688_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_7_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2652_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_63_enex5
        ) begin
      reg_act_regs_data_1_7_3_enexo <= act_regs_data_and_2652_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_7_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2556_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_63_enex5
        ) begin
      reg_act_regs_data_3_7_3_enexo <= act_regs_data_and_2556_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_7_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2604_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_63_enex5
        ) begin
      reg_act_regs_data_2_7_3_enexo <= act_regs_data_and_2604_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_27 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_64_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_27 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_27 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_64_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_27 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_27 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_64_enex5
        ) begin
      reg_act_config_inst_counter_enexo_27 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_6_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2557_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_64_enex5
        ) begin
      reg_act_regs_data_3_6_1_enexo <= act_regs_data_and_2557_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_6_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2653_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_64_enex5
        ) begin
      reg_act_regs_data_1_6_1_enexo <= act_regs_data_and_2653_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_6_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2605_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_64_enex5
        ) begin
      reg_act_regs_data_2_6_1_enexo <= act_regs_data_and_2605_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_6_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2689_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_64_enex5
        ) begin
      reg_act_regs_data_0_6_1_enexo <= act_regs_data_and_2689_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_28 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_65_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_28 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_28 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_65_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_28 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_28 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_65_enex5
        ) begin
      reg_act_config_inst_counter_enexo_28 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_6_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2606_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_65_enex5
        ) begin
      reg_act_regs_data_2_6_2_enexo <= act_regs_data_and_2606_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_6_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2654_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_65_enex5
        ) begin
      reg_act_regs_data_1_6_2_enexo <= act_regs_data_and_2654_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_6_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2558_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_65_enex5
        ) begin
      reg_act_regs_data_3_6_2_enexo <= act_regs_data_and_2558_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_6_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2690_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_65_enex5
        ) begin
      reg_act_regs_data_0_6_2_enexo <= act_regs_data_and_2690_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_29 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_66_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_29 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_29 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_66_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_29 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_29 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_66_enex5
        ) begin
      reg_act_config_inst_counter_enexo_29 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_6_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2607_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_66_enex5
        ) begin
      reg_act_regs_data_2_6_3_enexo <= act_regs_data_and_2607_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_6_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2559_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_66_enex5
        ) begin
      reg_act_regs_data_3_6_3_enexo <= act_regs_data_and_2559_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_6_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2691_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_66_enex5
        ) begin
      reg_act_regs_data_0_6_3_enexo <= act_regs_data_and_2691_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_6_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2655_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_66_enex5
        ) begin
      reg_act_regs_data_1_6_3_enexo <= act_regs_data_and_2655_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_30 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_67_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_30 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_30 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_67_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_30 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_30 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_67_enex5
        ) begin
      reg_act_config_inst_counter_enexo_30 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_5_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2560_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_67_enex5
        ) begin
      reg_act_regs_data_3_5_1_enexo <= act_regs_data_and_2560_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_5_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2692_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_67_enex5
        ) begin
      reg_act_regs_data_0_5_1_enexo <= act_regs_data_and_2692_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_5_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2656_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_67_enex5
        ) begin
      reg_act_regs_data_1_5_1_enexo <= act_regs_data_and_2656_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_5_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2608_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_67_enex5
        ) begin
      reg_act_regs_data_2_5_1_enexo <= act_regs_data_and_2608_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_31 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_68_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_31 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_31 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_68_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_31 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_31 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_68_enex5
        ) begin
      reg_act_config_inst_counter_enexo_31 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_5_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2609_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_68_enex5
        ) begin
      reg_act_regs_data_2_5_2_enexo <= act_regs_data_and_2609_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_5_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2657_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_68_enex5
        ) begin
      reg_act_regs_data_1_5_2_enexo <= act_regs_data_and_2657_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_5_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2561_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_68_enex5
        ) begin
      reg_act_regs_data_3_5_2_enexo <= act_regs_data_and_2561_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_5_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2693_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_68_enex5
        ) begin
      reg_act_regs_data_0_5_2_enexo <= act_regs_data_and_2693_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_32 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_69_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_32 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_32 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_69_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_32 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_5_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2694_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_69_enex5
        ) begin
      reg_act_regs_data_0_5_3_enexo <= act_regs_data_and_2694_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_32 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_69_enex5
        ) begin
      reg_act_config_inst_counter_enexo_32 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_5_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2658_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_69_enex5
        ) begin
      reg_act_regs_data_1_5_3_enexo <= act_regs_data_and_2658_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_5_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2562_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_69_enex5
        ) begin
      reg_act_regs_data_3_5_3_enexo <= act_regs_data_and_2562_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_5_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2610_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_69_enex5
        ) begin
      reg_act_regs_data_2_5_3_enexo <= act_regs_data_and_2610_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_33 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_70_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_33 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_33 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_70_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_33 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_33 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_70_enex5
        ) begin
      reg_act_config_inst_counter_enexo_33 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_4_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2563_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_70_enex5
        ) begin
      reg_act_regs_data_3_4_1_enexo <= act_regs_data_and_2563_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_4_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2695_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_70_enex5
        ) begin
      reg_act_regs_data_0_4_1_enexo <= act_regs_data_and_2695_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_4_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2611_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_70_enex5
        ) begin
      reg_act_regs_data_2_4_1_enexo <= act_regs_data_and_2611_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_4_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2659_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_70_enex5
        ) begin
      reg_act_regs_data_1_4_1_enexo <= act_regs_data_and_2659_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_34 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_71_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_34 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_34 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_71_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_34 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_34 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_71_enex5
        ) begin
      reg_act_config_inst_counter_enexo_34 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_4_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2564_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_71_enex5
        ) begin
      reg_act_regs_data_3_4_2_enexo <= act_regs_data_and_2564_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_4_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2660_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_71_enex5
        ) begin
      reg_act_regs_data_1_4_2_enexo <= act_regs_data_and_2660_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_4_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2696_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_71_enex5
        ) begin
      reg_act_regs_data_0_4_2_enexo <= act_regs_data_and_2696_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_4_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2612_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_71_enex5
        ) begin
      reg_act_regs_data_2_4_2_enexo <= act_regs_data_and_2612_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_35 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_72_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_35 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_35 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_72_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_35 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_35 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_72_enex5
        ) begin
      reg_act_config_inst_counter_enexo_35 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_4_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2697_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_72_enex5
        ) begin
      reg_act_regs_data_0_4_3_enexo <= act_regs_data_and_2697_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_4_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2661_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_72_enex5
        ) begin
      reg_act_regs_data_1_4_3_enexo <= act_regs_data_and_2661_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_4_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2565_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_72_enex5
        ) begin
      reg_act_regs_data_3_4_3_enexo <= act_regs_data_and_2565_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_4_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2613_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_72_enex5
        ) begin
      reg_act_regs_data_2_4_3_enexo <= act_regs_data_and_2613_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_36 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_73_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_36 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_36 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_73_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_36 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_36 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_73_enex5
        ) begin
      reg_act_config_inst_counter_enexo_36 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_3_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2698_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_73_enex5
        ) begin
      reg_act_regs_data_0_3_1_enexo <= act_regs_data_and_2698_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_3_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2566_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_73_enex5
        ) begin
      reg_act_regs_data_3_3_1_enexo <= act_regs_data_and_2566_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_3_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2662_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_73_enex5
        ) begin
      reg_act_regs_data_1_3_1_enexo <= act_regs_data_and_2662_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_3_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2614_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_73_enex5
        ) begin
      reg_act_regs_data_2_3_1_enexo <= act_regs_data_and_2614_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_37 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_74_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_37 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_37 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_74_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_37 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_37 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_74_enex5
        ) begin
      reg_act_config_inst_counter_enexo_37 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_3_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2699_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_74_enex5
        ) begin
      reg_act_regs_data_0_3_2_enexo <= act_regs_data_and_2699_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_3_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2663_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_74_enex5
        ) begin
      reg_act_regs_data_1_3_2_enexo <= act_regs_data_and_2663_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_3_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2567_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_74_enex5
        ) begin
      reg_act_regs_data_3_3_2_enexo <= act_regs_data_and_2567_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_3_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2615_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_74_enex5
        ) begin
      reg_act_regs_data_2_3_2_enexo <= act_regs_data_and_2615_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_38 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_75_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_38 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_38 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_75_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_38 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_38 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_75_enex5
        ) begin
      reg_act_config_inst_counter_enexo_38 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_3_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2700_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_75_enex5
        ) begin
      reg_act_regs_data_0_3_3_enexo <= act_regs_data_and_2700_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_3_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2568_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_75_enex5
        ) begin
      reg_act_regs_data_3_3_3_enexo <= act_regs_data_and_2568_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_3_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2664_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_75_enex5
        ) begin
      reg_act_regs_data_1_3_3_enexo <= act_regs_data_and_2664_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_3_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2616_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_75_enex5
        ) begin
      reg_act_regs_data_2_3_3_enexo <= act_regs_data_and_2616_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_2_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2617_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_76_enex5
        ) begin
      reg_act_regs_data_2_2_1_enexo <= act_regs_data_and_2617_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_39 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_76_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_39 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_39 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_76_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_39 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_39 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_76_enex5
        ) begin
      reg_act_config_inst_counter_enexo_39 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_2_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2569_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_76_enex5
        ) begin
      reg_act_regs_data_3_2_1_enexo <= act_regs_data_and_2569_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_2_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2665_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_76_enex5
        ) begin
      reg_act_regs_data_1_2_1_enexo <= act_regs_data_and_2665_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_2_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2701_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_76_enex5
        ) begin
      reg_act_regs_data_0_2_1_enexo <= act_regs_data_and_2701_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_40 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_77_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_40 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_40 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_77_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_40 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_40 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_77_enex5
        ) begin
      reg_act_config_inst_counter_enexo_40 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_2_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2702_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_77_enex5
        ) begin
      reg_act_regs_data_0_2_2_enexo <= act_regs_data_and_2702_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_2_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2666_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_77_enex5
        ) begin
      reg_act_regs_data_1_2_2_enexo <= act_regs_data_and_2666_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_2_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2570_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_77_enex5
        ) begin
      reg_act_regs_data_3_2_2_enexo <= act_regs_data_and_2570_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_2_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2618_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_77_enex5
        ) begin
      reg_act_regs_data_2_2_2_enexo <= act_regs_data_and_2618_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_41 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_78_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_41 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_41 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_78_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_41 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_41 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_78_enex5
        ) begin
      reg_act_config_inst_counter_enexo_41 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_2_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2571_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_78_enex5
        ) begin
      reg_act_regs_data_3_2_3_enexo <= act_regs_data_and_2571_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_2_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2619_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_78_enex5
        ) begin
      reg_act_regs_data_2_2_3_enexo <= act_regs_data_and_2619_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_2_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2703_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_78_enex5
        ) begin
      reg_act_regs_data_0_2_3_enexo <= act_regs_data_and_2703_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_2_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2667_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_78_enex5
        ) begin
      reg_act_regs_data_1_2_3_enexo <= act_regs_data_and_2667_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_42 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_79_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_42 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_42 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_79_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_42 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_1_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2620_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_79_enex5
        ) begin
      reg_act_regs_data_2_1_1_enexo <= act_regs_data_and_2620_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_42 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_79_enex5
        ) begin
      reg_act_config_inst_counter_enexo_42 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_1_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2572_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_79_enex5
        ) begin
      reg_act_regs_data_3_1_1_enexo <= act_regs_data_and_2572_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_1_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2761_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_79_enex5
        ) begin
      reg_act_regs_data_0_1_1_enexo <= act_regs_data_and_2761_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_1_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2668_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_79_enex5
        ) begin
      reg_act_regs_data_1_1_1_enexo <= act_regs_data_and_2668_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_43 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_80_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_43 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_43 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_80_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_43 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_43 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_80_enex5
        ) begin
      reg_act_config_inst_counter_enexo_43 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_1_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2669_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_80_enex5
        ) begin
      reg_act_regs_data_1_1_2_enexo <= act_regs_data_and_2669_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_1_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2573_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_80_enex5
        ) begin
      reg_act_regs_data_3_1_2_enexo <= act_regs_data_and_2573_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_1_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2762_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_80_enex5
        ) begin
      reg_act_regs_data_0_1_2_enexo <= act_regs_data_and_2762_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_1_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2621_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_80_enex5
        ) begin
      reg_act_regs_data_2_1_2_enexo <= act_regs_data_and_2621_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_44 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_81_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_44 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_44 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_81_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_44 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_44 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_81_enex5
        ) begin
      reg_act_config_inst_counter_enexo_44 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_1_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2763_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_81_enex5
        ) begin
      reg_act_regs_data_0_1_3_enexo <= act_regs_data_and_2763_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_1_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2574_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_81_enex5
        ) begin
      reg_act_regs_data_3_1_3_enexo <= act_regs_data_and_2574_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_1_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2670_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_81_enex5
        ) begin
      reg_act_regs_data_1_1_3_enexo <= act_regs_data_and_2670_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_1_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2622_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_81_enex5
        ) begin
      reg_act_regs_data_2_1_3_enexo <= act_regs_data_and_2622_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_45 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_82_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_45 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_0_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2575_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_82_enex5
        ) begin
      reg_act_regs_data_3_0_1_enexo <= act_regs_data_and_2575_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_45 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_82_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_45 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_45 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_82_enex5
        ) begin
      reg_act_config_inst_counter_enexo_45 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_0_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2764_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_82_enex5
        ) begin
      reg_act_regs_data_0_0_1_enexo <= act_regs_data_and_2764_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_0_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2623_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_82_enex5
        ) begin
      reg_act_regs_data_2_0_1_enexo <= act_regs_data_and_2623_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_0_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2671_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_82_enex5
        ) begin
      reg_act_regs_data_1_0_1_enexo <= act_regs_data_and_2671_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_46 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_83_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_46 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_46 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_83_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_46 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_46 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_83_enex5
        ) begin
      reg_act_config_inst_counter_enexo_46 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_0_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2576_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_83_enex5
        ) begin
      reg_act_regs_data_3_0_2_enexo <= act_regs_data_and_2576_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_0_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2765_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_83_enex5
        ) begin
      reg_act_regs_data_0_0_2_enexo <= act_regs_data_and_2765_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_0_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2672_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_83_enex5
        ) begin
      reg_act_regs_data_1_0_2_enexo <= act_regs_data_and_2672_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_0_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2624_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_83_enex5
        ) begin
      reg_act_regs_data_2_0_2_enexo <= act_regs_data_and_2624_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_47 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_84_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_47 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_47 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_84_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_47 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_47 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_84_enex5
        ) begin
      reg_act_config_inst_counter_enexo_47 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_0_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2577_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_84_enex5
        ) begin
      reg_act_regs_data_3_0_3_enexo <= act_regs_data_and_2577_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_0_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2766_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_84_enex5
        ) begin
      reg_act_regs_data_0_0_3_enexo <= act_regs_data_and_2766_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_0_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2625_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_84_enex5
        ) begin
      reg_act_regs_data_2_0_3_enexo <= act_regs_data_and_2625_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_0_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_2673_enex5 | nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_84_enex5
        ) begin
      reg_act_regs_data_1_0_3_enexo <= act_regs_data_and_2673_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_48 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Tanh_for_y_and_31_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_48 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_48 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Tanh_for_y_and_31_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_48 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_15_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2580_enex5 | Tanh_for_y_and_31_enex5 ) begin
      reg_act_regs_data_2_15_3_enexo_1 <= act_regs_data_and_2580_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_48 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Tanh_for_y_and_31_enex5 ) begin
      reg_act_config_inst_counter_enexo_48 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_15_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Tanh_for_y_and_31_enex5 ) begin
      reg_act_regs_data_1_15_enexo <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_15_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2674_enex5 | Tanh_for_y_and_31_enex5 ) begin
      reg_act_regs_data_0_15_1_enexo_1 <= act_regs_data_and_2674_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_15_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2626_enex5 | Tanh_for_y_and_31_enex5 ) begin
      reg_act_regs_data_1_15_1_enexo_1 <= act_regs_data_and_2626_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_15_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2676_enex5 | Tanh_for_y_and_31_enex5 ) begin
      reg_act_regs_data_0_15_3_enexo_1 <= act_regs_data_and_2676_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_15_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2628_enex5 | Tanh_for_y_and_31_enex5 ) begin
      reg_act_regs_data_1_15_3_enexo_1 <= act_regs_data_and_2628_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_15_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2531_enex5 | Tanh_for_y_and_31_enex5 ) begin
      reg_act_regs_data_3_15_2_enexo_1 <= act_regs_data_and_2531_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_15_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2532_enex5 | Tanh_for_y_and_31_enex5 ) begin
      reg_act_regs_data_3_15_3_enexo_1 <= act_regs_data_and_2532_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_15_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2579_enex5 | Tanh_for_y_and_31_enex5 ) begin
      reg_act_regs_data_2_15_2_enexo_1 <= act_regs_data_and_2579_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_15_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2675_enex5 | Tanh_for_y_and_31_enex5 ) begin
      reg_act_regs_data_0_15_2_enexo_1 <= act_regs_data_and_2675_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_15_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2578_enex5 | Tanh_for_y_and_31_enex5 ) begin
      reg_act_regs_data_2_15_1_enexo_1 <= act_regs_data_and_2578_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_15_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2530_enex5 | Tanh_for_y_and_31_enex5 ) begin
      reg_act_regs_data_3_15_1_enexo_1 <= act_regs_data_and_2530_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_15_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2627_enex5 | Tanh_for_y_and_31_enex5 ) begin
      reg_act_regs_data_1_15_2_enexo_1 <= act_regs_data_and_2627_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_49 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Tanh_for_y_and_32_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_49 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_49 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Tanh_for_y_and_32_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_49 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_15_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2580_enex5 | Tanh_for_y_and_32_enex5 ) begin
      reg_act_regs_data_2_15_3_enexo_2 <= act_regs_data_and_2580_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_49 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Tanh_for_y_and_32_enex5 ) begin
      reg_act_config_inst_counter_enexo_49 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_15_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Tanh_for_y_and_32_enex5 ) begin
      reg_act_regs_data_1_15_enexo_1 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_15_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2674_enex5 | Tanh_for_y_and_32_enex5 ) begin
      reg_act_regs_data_0_15_1_enexo_2 <= act_regs_data_and_2674_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_15_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2626_enex5 | Tanh_for_y_and_32_enex5 ) begin
      reg_act_regs_data_1_15_1_enexo_2 <= act_regs_data_and_2626_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_15_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2676_enex5 | Tanh_for_y_and_32_enex5 ) begin
      reg_act_regs_data_0_15_3_enexo_2 <= act_regs_data_and_2676_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_15_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2628_enex5 | Tanh_for_y_and_32_enex5 ) begin
      reg_act_regs_data_1_15_3_enexo_2 <= act_regs_data_and_2628_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_15_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2531_enex5 | Tanh_for_y_and_32_enex5 ) begin
      reg_act_regs_data_3_15_2_enexo_2 <= act_regs_data_and_2531_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_15_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2532_enex5 | Tanh_for_y_and_32_enex5 ) begin
      reg_act_regs_data_3_15_3_enexo_2 <= act_regs_data_and_2532_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_15_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2579_enex5 | Tanh_for_y_and_32_enex5 ) begin
      reg_act_regs_data_2_15_2_enexo_2 <= act_regs_data_and_2579_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_15_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2675_enex5 | Tanh_for_y_and_32_enex5 ) begin
      reg_act_regs_data_0_15_2_enexo_2 <= act_regs_data_and_2675_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_15_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2578_enex5 | Tanh_for_y_and_32_enex5 ) begin
      reg_act_regs_data_2_15_1_enexo_2 <= act_regs_data_and_2578_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_15_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2530_enex5 | Tanh_for_y_and_32_enex5 ) begin
      reg_act_regs_data_3_15_1_enexo_2 <= act_regs_data_and_2530_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_15_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2627_enex5 | Tanh_for_y_and_32_enex5 ) begin
      reg_act_regs_data_1_15_2_enexo_2 <= act_regs_data_and_2627_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_50 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Tanh_for_y_and_33_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_50 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_14_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2678_enex5 | Tanh_for_y_and_33_enex5 ) begin
      reg_act_regs_data_0_14_2_enexo_1 <= act_regs_data_and_2678_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_14_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2629_enex5 | Tanh_for_y_and_33_enex5 ) begin
      reg_act_regs_data_1_14_1_enexo_1 <= act_regs_data_and_2629_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_50 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Tanh_for_y_and_33_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_50 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_50 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Tanh_for_y_and_33_enex5 ) begin
      reg_act_config_inst_counter_enexo_50 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_14_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Tanh_for_y_and_33_enex5 ) begin
      reg_act_regs_data_0_14_enexo <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_14_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2582_enex5 | Tanh_for_y_and_33_enex5 ) begin
      reg_act_regs_data_2_14_2_enexo_1 <= act_regs_data_and_2582_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_14_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2679_enex5 | Tanh_for_y_and_33_enex5 ) begin
      reg_act_regs_data_0_14_3_enexo_1 <= act_regs_data_and_2679_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_14_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2534_enex5 | Tanh_for_y_and_33_enex5 ) begin
      reg_act_regs_data_3_14_2_enexo_1 <= act_regs_data_and_2534_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_14_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2581_enex5 | Tanh_for_y_and_33_enex5 ) begin
      reg_act_regs_data_2_14_1_enexo_1 <= act_regs_data_and_2581_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_14_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2630_enex5 | Tanh_for_y_and_33_enex5 ) begin
      reg_act_regs_data_1_14_2_enexo_1 <= act_regs_data_and_2630_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_14_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2533_enex5 | Tanh_for_y_and_33_enex5 ) begin
      reg_act_regs_data_3_14_1_enexo_1 <= act_regs_data_and_2533_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_14_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2583_enex5 | Tanh_for_y_and_33_enex5 ) begin
      reg_act_regs_data_2_14_3_enexo_1 <= act_regs_data_and_2583_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_14_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2677_enex5 | Tanh_for_y_and_33_enex5 ) begin
      reg_act_regs_data_0_14_1_enexo_1 <= act_regs_data_and_2677_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_14_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2535_enex5 | Tanh_for_y_and_33_enex5 ) begin
      reg_act_regs_data_3_14_3_enexo_1 <= act_regs_data_and_2535_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_14_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2631_enex5 | Tanh_for_y_and_33_enex5 ) begin
      reg_act_regs_data_1_14_3_enexo_1 <= act_regs_data_and_2631_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_51 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Tanh_for_y_and_34_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_51 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_14_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2678_enex5 | Tanh_for_y_and_34_enex5 ) begin
      reg_act_regs_data_0_14_2_enexo_2 <= act_regs_data_and_2678_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_14_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2629_enex5 | Tanh_for_y_and_34_enex5 ) begin
      reg_act_regs_data_1_14_1_enexo_2 <= act_regs_data_and_2629_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_51 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Tanh_for_y_and_34_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_51 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_51 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Tanh_for_y_and_34_enex5 ) begin
      reg_act_config_inst_counter_enexo_51 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_14_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Tanh_for_y_and_34_enex5 ) begin
      reg_act_regs_data_0_14_enexo_1 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_14_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2582_enex5 | Tanh_for_y_and_34_enex5 ) begin
      reg_act_regs_data_2_14_2_enexo_2 <= act_regs_data_and_2582_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_14_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2679_enex5 | Tanh_for_y_and_34_enex5 ) begin
      reg_act_regs_data_0_14_3_enexo_2 <= act_regs_data_and_2679_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_14_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2534_enex5 | Tanh_for_y_and_34_enex5 ) begin
      reg_act_regs_data_3_14_2_enexo_2 <= act_regs_data_and_2534_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_14_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2581_enex5 | Tanh_for_y_and_34_enex5 ) begin
      reg_act_regs_data_2_14_1_enexo_2 <= act_regs_data_and_2581_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_14_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2630_enex5 | Tanh_for_y_and_34_enex5 ) begin
      reg_act_regs_data_1_14_2_enexo_2 <= act_regs_data_and_2630_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_14_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2533_enex5 | Tanh_for_y_and_34_enex5 ) begin
      reg_act_regs_data_3_14_1_enexo_2 <= act_regs_data_and_2533_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_14_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2583_enex5 | Tanh_for_y_and_34_enex5 ) begin
      reg_act_regs_data_2_14_3_enexo_2 <= act_regs_data_and_2583_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_14_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2677_enex5 | Tanh_for_y_and_34_enex5 ) begin
      reg_act_regs_data_0_14_1_enexo_2 <= act_regs_data_and_2677_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_14_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2535_enex5 | Tanh_for_y_and_34_enex5 ) begin
      reg_act_regs_data_3_14_3_enexo_2 <= act_regs_data_and_2535_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_14_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2631_enex5 | Tanh_for_y_and_34_enex5 ) begin
      reg_act_regs_data_1_14_3_enexo_2 <= act_regs_data_and_2631_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_13_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2537_enex5 | Tanh_for_y_and_35_enex5 ) begin
      reg_act_regs_data_3_13_2_enexo_1 <= act_regs_data_and_2537_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_52 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Tanh_for_y_and_35_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_52 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_13_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2632_enex5 | Tanh_for_y_and_35_enex5 ) begin
      reg_act_regs_data_1_13_1_enexo_1 <= act_regs_data_and_2632_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_13_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2584_enex5 | Tanh_for_y_and_35_enex5 ) begin
      reg_act_regs_data_2_13_1_enexo_1 <= act_regs_data_and_2584_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_52 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Tanh_for_y_and_35_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_52 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_13_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2750_enex5 | Tanh_for_y_and_35_enex5 ) begin
      reg_act_regs_data_0_13_2_enexo_1 <= act_regs_data_and_2750_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_52 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Tanh_for_y_and_35_enex5 ) begin
      reg_act_config_inst_counter_enexo_52 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_13_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2749_enex5 | Tanh_for_y_and_35_enex5 ) begin
      reg_act_regs_data_0_13_1_enexo_1 <= act_regs_data_and_2749_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_13_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2633_enex5 | Tanh_for_y_and_35_enex5 ) begin
      reg_act_regs_data_1_13_2_enexo_1 <= act_regs_data_and_2633_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_13_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Tanh_for_y_and_35_enex5 ) begin
      reg_act_regs_data_3_13_enexo <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_13_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2586_enex5 | Tanh_for_y_and_35_enex5 ) begin
      reg_act_regs_data_2_13_3_enexo_1 <= act_regs_data_and_2586_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_13_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2585_enex5 | Tanh_for_y_and_35_enex5 ) begin
      reg_act_regs_data_2_13_2_enexo_1 <= act_regs_data_and_2585_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_13_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2538_enex5 | Tanh_for_y_and_35_enex5 ) begin
      reg_act_regs_data_3_13_3_enexo_1 <= act_regs_data_and_2538_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_13_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2536_enex5 | Tanh_for_y_and_35_enex5 ) begin
      reg_act_regs_data_3_13_1_enexo_1 <= act_regs_data_and_2536_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_13_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2634_enex5 | Tanh_for_y_and_35_enex5 ) begin
      reg_act_regs_data_1_13_3_enexo_1 <= act_regs_data_and_2634_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_13_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2751_enex5 | Tanh_for_y_and_35_enex5 ) begin
      reg_act_regs_data_0_13_3_enexo_1 <= act_regs_data_and_2751_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_13_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2537_enex5 | Tanh_for_y_and_36_enex5 ) begin
      reg_act_regs_data_3_13_2_enexo_2 <= act_regs_data_and_2537_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_53 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Tanh_for_y_and_36_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_53 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_13_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2632_enex5 | Tanh_for_y_and_36_enex5 ) begin
      reg_act_regs_data_1_13_1_enexo_2 <= act_regs_data_and_2632_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_13_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2584_enex5 | Tanh_for_y_and_36_enex5 ) begin
      reg_act_regs_data_2_13_1_enexo_2 <= act_regs_data_and_2584_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_53 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Tanh_for_y_and_36_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_53 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_13_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2750_enex5 | Tanh_for_y_and_36_enex5 ) begin
      reg_act_regs_data_0_13_2_enexo_2 <= act_regs_data_and_2750_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_53 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Tanh_for_y_and_36_enex5 ) begin
      reg_act_config_inst_counter_enexo_53 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_13_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2749_enex5 | Tanh_for_y_and_36_enex5 ) begin
      reg_act_regs_data_0_13_1_enexo_2 <= act_regs_data_and_2749_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_13_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2633_enex5 | Tanh_for_y_and_36_enex5 ) begin
      reg_act_regs_data_1_13_2_enexo_2 <= act_regs_data_and_2633_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_13_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Tanh_for_y_and_36_enex5 ) begin
      reg_act_regs_data_3_13_enexo_1 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_13_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2586_enex5 | Tanh_for_y_and_36_enex5 ) begin
      reg_act_regs_data_2_13_3_enexo_2 <= act_regs_data_and_2586_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_13_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2585_enex5 | Tanh_for_y_and_36_enex5 ) begin
      reg_act_regs_data_2_13_2_enexo_2 <= act_regs_data_and_2585_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_13_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2538_enex5 | Tanh_for_y_and_36_enex5 ) begin
      reg_act_regs_data_3_13_3_enexo_2 <= act_regs_data_and_2538_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_13_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2536_enex5 | Tanh_for_y_and_36_enex5 ) begin
      reg_act_regs_data_3_13_1_enexo_2 <= act_regs_data_and_2536_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_13_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2634_enex5 | Tanh_for_y_and_36_enex5 ) begin
      reg_act_regs_data_1_13_3_enexo_2 <= act_regs_data_and_2634_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_13_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2751_enex5 | Tanh_for_y_and_36_enex5 ) begin
      reg_act_regs_data_0_13_3_enexo_2 <= act_regs_data_and_2751_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_54 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Tanh_for_y_and_37_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_54 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_54 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Tanh_for_y_and_37_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_54 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_12_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2588_enex5 | Tanh_for_y_and_37_enex5 ) begin
      reg_act_regs_data_2_12_2_enexo_1 <= act_regs_data_and_2588_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_54 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Tanh_for_y_and_37_enex5 ) begin
      reg_act_config_inst_counter_enexo_54 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_12_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2587_enex5 | Tanh_for_y_and_37_enex5 ) begin
      reg_act_regs_data_2_12_1_enexo_1 <= act_regs_data_and_2587_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_12_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Tanh_for_y_and_37_enex5 ) begin
      reg_act_regs_data_0_12_enexo <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_12_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2752_enex5 | Tanh_for_y_and_37_enex5 ) begin
      reg_act_regs_data_0_12_1_enexo_1 <= act_regs_data_and_2752_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_12_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2635_enex5 | Tanh_for_y_and_37_enex5 ) begin
      reg_act_regs_data_1_12_1_enexo_1 <= act_regs_data_and_2635_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_12_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2753_enex5 | Tanh_for_y_and_37_enex5 ) begin
      reg_act_regs_data_0_12_2_enexo_1 <= act_regs_data_and_2753_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_12_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2754_enex5 | Tanh_for_y_and_37_enex5 ) begin
      reg_act_regs_data_0_12_3_enexo_1 <= act_regs_data_and_2754_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_12_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2540_enex5 | Tanh_for_y_and_37_enex5 ) begin
      reg_act_regs_data_3_12_2_enexo_1 <= act_regs_data_and_2540_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_12_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2589_enex5 | Tanh_for_y_and_37_enex5 ) begin
      reg_act_regs_data_2_12_3_enexo_1 <= act_regs_data_and_2589_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_12_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2541_enex5 | Tanh_for_y_and_37_enex5 ) begin
      reg_act_regs_data_3_12_3_enexo_1 <= act_regs_data_and_2541_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_12_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2636_enex5 | Tanh_for_y_and_37_enex5 ) begin
      reg_act_regs_data_1_12_2_enexo_1 <= act_regs_data_and_2636_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_12_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2637_enex5 | Tanh_for_y_and_37_enex5 ) begin
      reg_act_regs_data_1_12_3_enexo_1 <= act_regs_data_and_2637_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_12_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2539_enex5 | Tanh_for_y_and_37_enex5 ) begin
      reg_act_regs_data_3_12_1_enexo_1 <= act_regs_data_and_2539_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_55 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Tanh_for_y_and_38_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_55 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_55 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Tanh_for_y_and_38_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_55 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_12_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2588_enex5 | Tanh_for_y_and_38_enex5 ) begin
      reg_act_regs_data_2_12_2_enexo_2 <= act_regs_data_and_2588_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_55 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Tanh_for_y_and_38_enex5 ) begin
      reg_act_config_inst_counter_enexo_55 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_12_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2587_enex5 | Tanh_for_y_and_38_enex5 ) begin
      reg_act_regs_data_2_12_1_enexo_2 <= act_regs_data_and_2587_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_12_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Tanh_for_y_and_38_enex5 ) begin
      reg_act_regs_data_0_12_enexo_1 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_12_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2752_enex5 | Tanh_for_y_and_38_enex5 ) begin
      reg_act_regs_data_0_12_1_enexo_2 <= act_regs_data_and_2752_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_12_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2635_enex5 | Tanh_for_y_and_38_enex5 ) begin
      reg_act_regs_data_1_12_1_enexo_2 <= act_regs_data_and_2635_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_12_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2753_enex5 | Tanh_for_y_and_38_enex5 ) begin
      reg_act_regs_data_0_12_2_enexo_2 <= act_regs_data_and_2753_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_12_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2754_enex5 | Tanh_for_y_and_38_enex5 ) begin
      reg_act_regs_data_0_12_3_enexo_2 <= act_regs_data_and_2754_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_12_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2540_enex5 | Tanh_for_y_and_38_enex5 ) begin
      reg_act_regs_data_3_12_2_enexo_2 <= act_regs_data_and_2540_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_12_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2589_enex5 | Tanh_for_y_and_38_enex5 ) begin
      reg_act_regs_data_2_12_3_enexo_2 <= act_regs_data_and_2589_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_12_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2541_enex5 | Tanh_for_y_and_38_enex5 ) begin
      reg_act_regs_data_3_12_3_enexo_2 <= act_regs_data_and_2541_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_12_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2636_enex5 | Tanh_for_y_and_38_enex5 ) begin
      reg_act_regs_data_1_12_2_enexo_2 <= act_regs_data_and_2636_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_12_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2637_enex5 | Tanh_for_y_and_38_enex5 ) begin
      reg_act_regs_data_1_12_3_enexo_2 <= act_regs_data_and_2637_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_12_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2539_enex5 | Tanh_for_y_and_38_enex5 ) begin
      reg_act_regs_data_3_12_1_enexo_2 <= act_regs_data_and_2539_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_56 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Tanh_for_y_and_39_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_56 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_11_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Tanh_for_y_and_39_enex5 ) begin
      reg_act_regs_data_2_11_enexo <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_56 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Tanh_for_y_and_39_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_56 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_56 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Tanh_for_y_and_39_enex5 ) begin
      reg_act_config_inst_counter_enexo_56 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_11_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2757_enex5 | Tanh_for_y_and_39_enex5 ) begin
      reg_act_regs_data_0_11_3_enexo_1 <= act_regs_data_and_2757_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_11_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2590_enex5 | Tanh_for_y_and_39_enex5 ) begin
      reg_act_regs_data_2_11_1_enexo_1 <= act_regs_data_and_2590_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_11_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2640_enex5 | Tanh_for_y_and_39_enex5 ) begin
      reg_act_regs_data_1_11_3_enexo_1 <= act_regs_data_and_2640_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_11_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2591_enex5 | Tanh_for_y_and_39_enex5 ) begin
      reg_act_regs_data_2_11_2_enexo_1 <= act_regs_data_and_2591_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_11_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2756_enex5 | Tanh_for_y_and_39_enex5 ) begin
      reg_act_regs_data_0_11_2_enexo_1 <= act_regs_data_and_2756_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_11_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2592_enex5 | Tanh_for_y_and_39_enex5 ) begin
      reg_act_regs_data_2_11_3_enexo_1 <= act_regs_data_and_2592_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_11_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2542_enex5 | Tanh_for_y_and_39_enex5 ) begin
      reg_act_regs_data_3_11_1_enexo_1 <= act_regs_data_and_2542_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_11_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2755_enex5 | Tanh_for_y_and_39_enex5 ) begin
      reg_act_regs_data_0_11_1_enexo_1 <= act_regs_data_and_2755_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_11_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2544_enex5 | Tanh_for_y_and_39_enex5 ) begin
      reg_act_regs_data_3_11_3_enexo_1 <= act_regs_data_and_2544_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_11_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2543_enex5 | Tanh_for_y_and_39_enex5 ) begin
      reg_act_regs_data_3_11_2_enexo_1 <= act_regs_data_and_2543_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_11_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2638_enex5 | Tanh_for_y_and_39_enex5 ) begin
      reg_act_regs_data_1_11_1_enexo_1 <= act_regs_data_and_2638_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_11_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2639_enex5 | Tanh_for_y_and_39_enex5 ) begin
      reg_act_regs_data_1_11_2_enexo_1 <= act_regs_data_and_2639_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_57 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Tanh_for_y_and_40_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_57 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_11_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Tanh_for_y_and_40_enex5 ) begin
      reg_act_regs_data_2_11_enexo_1 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_57 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Tanh_for_y_and_40_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_57 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_57 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Tanh_for_y_and_40_enex5 ) begin
      reg_act_config_inst_counter_enexo_57 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_11_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2757_enex5 | Tanh_for_y_and_40_enex5 ) begin
      reg_act_regs_data_0_11_3_enexo_2 <= act_regs_data_and_2757_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_11_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2590_enex5 | Tanh_for_y_and_40_enex5 ) begin
      reg_act_regs_data_2_11_1_enexo_2 <= act_regs_data_and_2590_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_11_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2640_enex5 | Tanh_for_y_and_40_enex5 ) begin
      reg_act_regs_data_1_11_3_enexo_2 <= act_regs_data_and_2640_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_11_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2591_enex5 | Tanh_for_y_and_40_enex5 ) begin
      reg_act_regs_data_2_11_2_enexo_2 <= act_regs_data_and_2591_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_11_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2756_enex5 | Tanh_for_y_and_40_enex5 ) begin
      reg_act_regs_data_0_11_2_enexo_2 <= act_regs_data_and_2756_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_11_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2592_enex5 | Tanh_for_y_and_40_enex5 ) begin
      reg_act_regs_data_2_11_3_enexo_2 <= act_regs_data_and_2592_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_11_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2542_enex5 | Tanh_for_y_and_40_enex5 ) begin
      reg_act_regs_data_3_11_1_enexo_2 <= act_regs_data_and_2542_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_11_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2755_enex5 | Tanh_for_y_and_40_enex5 ) begin
      reg_act_regs_data_0_11_1_enexo_2 <= act_regs_data_and_2755_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_11_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2544_enex5 | Tanh_for_y_and_40_enex5 ) begin
      reg_act_regs_data_3_11_3_enexo_2 <= act_regs_data_and_2544_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_11_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2543_enex5 | Tanh_for_y_and_40_enex5 ) begin
      reg_act_regs_data_3_11_2_enexo_2 <= act_regs_data_and_2543_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_11_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2638_enex5 | Tanh_for_y_and_40_enex5 ) begin
      reg_act_regs_data_1_11_1_enexo_2 <= act_regs_data_and_2638_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_11_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2639_enex5 | Tanh_for_y_and_40_enex5 ) begin
      reg_act_regs_data_1_11_2_enexo_2 <= act_regs_data_and_2639_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_58 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Tanh_for_y_and_41_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_58 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_58 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Tanh_for_y_and_41_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_58 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_58 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Tanh_for_y_and_41_enex5 ) begin
      reg_act_config_inst_counter_enexo_58 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_10_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2641_enex5 | Tanh_for_y_and_41_enex5 ) begin
      reg_act_regs_data_1_10_1_enexo_1 <= act_regs_data_and_2641_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_10_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2642_enex5 | Tanh_for_y_and_41_enex5 ) begin
      reg_act_regs_data_1_10_2_enexo_1 <= act_regs_data_and_2642_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_10_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2547_enex5 | Tanh_for_y_and_41_enex5 ) begin
      reg_act_regs_data_3_10_3_enexo_1 <= act_regs_data_and_2547_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_10_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2593_enex5 | Tanh_for_y_and_41_enex5 ) begin
      reg_act_regs_data_2_10_1_enexo_1 <= act_regs_data_and_2593_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_10_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Tanh_for_y_and_41_enex5 ) begin
      reg_act_regs_data_0_10_enexo <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_10_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2759_enex5 | Tanh_for_y_and_41_enex5 ) begin
      reg_act_regs_data_0_10_2_enexo_1 <= act_regs_data_and_2759_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_10_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2760_enex5 | Tanh_for_y_and_41_enex5 ) begin
      reg_act_regs_data_0_10_3_enexo_1 <= act_regs_data_and_2760_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_10_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2545_enex5 | Tanh_for_y_and_41_enex5 ) begin
      reg_act_regs_data_3_10_1_enexo_1 <= act_regs_data_and_2545_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_10_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2595_enex5 | Tanh_for_y_and_41_enex5 ) begin
      reg_act_regs_data_2_10_3_enexo_1 <= act_regs_data_and_2595_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_10_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2643_enex5 | Tanh_for_y_and_41_enex5 ) begin
      reg_act_regs_data_1_10_3_enexo_1 <= act_regs_data_and_2643_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_10_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2758_enex5 | Tanh_for_y_and_41_enex5 ) begin
      reg_act_regs_data_0_10_1_enexo_1 <= act_regs_data_and_2758_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_10_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2546_enex5 | Tanh_for_y_and_41_enex5 ) begin
      reg_act_regs_data_3_10_2_enexo_1 <= act_regs_data_and_2546_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_10_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2594_enex5 | Tanh_for_y_and_41_enex5 ) begin
      reg_act_regs_data_2_10_2_enexo_1 <= act_regs_data_and_2594_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_59 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Tanh_for_y_and_42_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_59 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_59 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Tanh_for_y_and_42_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_59 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_59 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Tanh_for_y_and_42_enex5 ) begin
      reg_act_config_inst_counter_enexo_59 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_10_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2641_enex5 | Tanh_for_y_and_42_enex5 ) begin
      reg_act_regs_data_1_10_1_enexo_2 <= act_regs_data_and_2641_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_10_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2642_enex5 | Tanh_for_y_and_42_enex5 ) begin
      reg_act_regs_data_1_10_2_enexo_2 <= act_regs_data_and_2642_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_10_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2547_enex5 | Tanh_for_y_and_42_enex5 ) begin
      reg_act_regs_data_3_10_3_enexo_2 <= act_regs_data_and_2547_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_10_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2593_enex5 | Tanh_for_y_and_42_enex5 ) begin
      reg_act_regs_data_2_10_1_enexo_2 <= act_regs_data_and_2593_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_10_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Tanh_for_y_and_42_enex5 ) begin
      reg_act_regs_data_0_10_enexo_1 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_10_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2759_enex5 | Tanh_for_y_and_42_enex5 ) begin
      reg_act_regs_data_0_10_2_enexo_2 <= act_regs_data_and_2759_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_10_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2760_enex5 | Tanh_for_y_and_42_enex5 ) begin
      reg_act_regs_data_0_10_3_enexo_2 <= act_regs_data_and_2760_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_10_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2545_enex5 | Tanh_for_y_and_42_enex5 ) begin
      reg_act_regs_data_3_10_1_enexo_2 <= act_regs_data_and_2545_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_10_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2595_enex5 | Tanh_for_y_and_42_enex5 ) begin
      reg_act_regs_data_2_10_3_enexo_2 <= act_regs_data_and_2595_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_10_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2643_enex5 | Tanh_for_y_and_42_enex5 ) begin
      reg_act_regs_data_1_10_3_enexo_2 <= act_regs_data_and_2643_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_10_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2758_enex5 | Tanh_for_y_and_42_enex5 ) begin
      reg_act_regs_data_0_10_1_enexo_2 <= act_regs_data_and_2758_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_10_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2546_enex5 | Tanh_for_y_and_42_enex5 ) begin
      reg_act_regs_data_3_10_2_enexo_2 <= act_regs_data_and_2546_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_10_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2594_enex5 | Tanh_for_y_and_42_enex5 ) begin
      reg_act_regs_data_2_10_2_enexo_2 <= act_regs_data_and_2594_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_60 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Tanh_for_y_and_43_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_60 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_60 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Tanh_for_y_and_43_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_60 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_60 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Tanh_for_y_and_43_enex5 ) begin
      reg_act_config_inst_counter_enexo_60 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_9_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2646_enex5 | Tanh_for_y_and_43_enex5 ) begin
      reg_act_regs_data_1_9_3_enexo_1 <= act_regs_data_and_2646_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_9_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2681_enex5 | Tanh_for_y_and_43_enex5 ) begin
      reg_act_regs_data_0_9_2_enexo_1 <= act_regs_data_and_2681_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_9_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2644_enex5 | Tanh_for_y_and_43_enex5 ) begin
      reg_act_regs_data_1_9_1_enexo_1 <= act_regs_data_and_2644_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_9_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Tanh_for_y_and_43_enex5 ) begin
      reg_act_regs_data_1_9_enexo <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_9_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2682_enex5 | Tanh_for_y_and_43_enex5 ) begin
      reg_act_regs_data_0_9_3_enexo_1 <= act_regs_data_and_2682_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_9_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2598_enex5 | Tanh_for_y_and_43_enex5 ) begin
      reg_act_regs_data_2_9_3_enexo_1 <= act_regs_data_and_2598_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_9_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2597_enex5 | Tanh_for_y_and_43_enex5 ) begin
      reg_act_regs_data_2_9_2_enexo_1 <= act_regs_data_and_2597_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_9_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2548_enex5 | Tanh_for_y_and_43_enex5 ) begin
      reg_act_regs_data_3_9_1_enexo_1 <= act_regs_data_and_2548_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_9_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2645_enex5 | Tanh_for_y_and_43_enex5 ) begin
      reg_act_regs_data_1_9_2_enexo_1 <= act_regs_data_and_2645_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_9_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2549_enex5 | Tanh_for_y_and_43_enex5 ) begin
      reg_act_regs_data_3_9_2_enexo_1 <= act_regs_data_and_2549_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_9_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2680_enex5 | Tanh_for_y_and_43_enex5 ) begin
      reg_act_regs_data_0_9_1_enexo_1 <= act_regs_data_and_2680_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_9_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2550_enex5 | Tanh_for_y_and_43_enex5 ) begin
      reg_act_regs_data_3_9_3_enexo_1 <= act_regs_data_and_2550_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_9_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2596_enex5 | Tanh_for_y_and_43_enex5 ) begin
      reg_act_regs_data_2_9_1_enexo_1 <= act_regs_data_and_2596_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_61 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Tanh_for_y_and_44_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_61 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_61 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Tanh_for_y_and_44_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_61 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_61 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Tanh_for_y_and_44_enex5 ) begin
      reg_act_config_inst_counter_enexo_61 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_9_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2646_enex5 | Tanh_for_y_and_44_enex5 ) begin
      reg_act_regs_data_1_9_3_enexo_2 <= act_regs_data_and_2646_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_9_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2681_enex5 | Tanh_for_y_and_44_enex5 ) begin
      reg_act_regs_data_0_9_2_enexo_2 <= act_regs_data_and_2681_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_9_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2644_enex5 | Tanh_for_y_and_44_enex5 ) begin
      reg_act_regs_data_1_9_1_enexo_2 <= act_regs_data_and_2644_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_9_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Tanh_for_y_and_44_enex5 ) begin
      reg_act_regs_data_1_9_enexo_1 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_9_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2682_enex5 | Tanh_for_y_and_44_enex5 ) begin
      reg_act_regs_data_0_9_3_enexo_2 <= act_regs_data_and_2682_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_9_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2598_enex5 | Tanh_for_y_and_44_enex5 ) begin
      reg_act_regs_data_2_9_3_enexo_2 <= act_regs_data_and_2598_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_9_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2597_enex5 | Tanh_for_y_and_44_enex5 ) begin
      reg_act_regs_data_2_9_2_enexo_2 <= act_regs_data_and_2597_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_9_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2548_enex5 | Tanh_for_y_and_44_enex5 ) begin
      reg_act_regs_data_3_9_1_enexo_2 <= act_regs_data_and_2548_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_9_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2645_enex5 | Tanh_for_y_and_44_enex5 ) begin
      reg_act_regs_data_1_9_2_enexo_2 <= act_regs_data_and_2645_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_9_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2549_enex5 | Tanh_for_y_and_44_enex5 ) begin
      reg_act_regs_data_3_9_2_enexo_2 <= act_regs_data_and_2549_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_9_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2680_enex5 | Tanh_for_y_and_44_enex5 ) begin
      reg_act_regs_data_0_9_1_enexo_2 <= act_regs_data_and_2680_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_9_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2550_enex5 | Tanh_for_y_and_44_enex5 ) begin
      reg_act_regs_data_3_9_3_enexo_2 <= act_regs_data_and_2550_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_9_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2596_enex5 | Tanh_for_y_and_44_enex5 ) begin
      reg_act_regs_data_2_9_1_enexo_2 <= act_regs_data_and_2596_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_62 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Tanh_for_y_and_45_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_62 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_62 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Tanh_for_y_and_45_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_62 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_62 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Tanh_for_y_and_45_enex5 ) begin
      reg_act_config_inst_counter_enexo_62 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_8_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Tanh_for_y_and_45_enex5 ) begin
      reg_act_regs_data_2_8_enexo <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_8_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2684_enex5 | Tanh_for_y_and_45_enex5 ) begin
      reg_act_regs_data_0_8_2_enexo_1 <= act_regs_data_and_2684_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_8_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2648_enex5 | Tanh_for_y_and_45_enex5 ) begin
      reg_act_regs_data_1_8_2_enexo_1 <= act_regs_data_and_2648_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_8_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2599_enex5 | Tanh_for_y_and_45_enex5 ) begin
      reg_act_regs_data_2_8_1_enexo_1 <= act_regs_data_and_2599_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_8_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2683_enex5 | Tanh_for_y_and_45_enex5 ) begin
      reg_act_regs_data_0_8_1_enexo_1 <= act_regs_data_and_2683_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_8_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2685_enex5 | Tanh_for_y_and_45_enex5 ) begin
      reg_act_regs_data_0_8_3_enexo_1 <= act_regs_data_and_2685_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_8_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2600_enex5 | Tanh_for_y_and_45_enex5 ) begin
      reg_act_regs_data_2_8_2_enexo_1 <= act_regs_data_and_2600_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_8_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2551_enex5 | Tanh_for_y_and_45_enex5 ) begin
      reg_act_regs_data_3_8_1_enexo_1 <= act_regs_data_and_2551_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_8_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2601_enex5 | Tanh_for_y_and_45_enex5 ) begin
      reg_act_regs_data_2_8_3_enexo_1 <= act_regs_data_and_2601_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_8_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2552_enex5 | Tanh_for_y_and_45_enex5 ) begin
      reg_act_regs_data_3_8_2_enexo_1 <= act_regs_data_and_2552_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_8_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2647_enex5 | Tanh_for_y_and_45_enex5 ) begin
      reg_act_regs_data_1_8_1_enexo_1 <= act_regs_data_and_2647_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_8_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2649_enex5 | Tanh_for_y_and_45_enex5 ) begin
      reg_act_regs_data_1_8_3_enexo_1 <= act_regs_data_and_2649_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_8_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2553_enex5 | Tanh_for_y_and_45_enex5 ) begin
      reg_act_regs_data_3_8_3_enexo_1 <= act_regs_data_and_2553_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_63 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Tanh_for_y_and_46_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_63 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_63 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Tanh_for_y_and_46_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_63 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_63 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Tanh_for_y_and_46_enex5 ) begin
      reg_act_config_inst_counter_enexo_63 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_8_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Tanh_for_y_and_46_enex5 ) begin
      reg_act_regs_data_2_8_enexo_1 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_8_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2684_enex5 | Tanh_for_y_and_46_enex5 ) begin
      reg_act_regs_data_0_8_2_enexo_2 <= act_regs_data_and_2684_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_8_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2648_enex5 | Tanh_for_y_and_46_enex5 ) begin
      reg_act_regs_data_1_8_2_enexo_2 <= act_regs_data_and_2648_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_8_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2599_enex5 | Tanh_for_y_and_46_enex5 ) begin
      reg_act_regs_data_2_8_1_enexo_2 <= act_regs_data_and_2599_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_8_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2683_enex5 | Tanh_for_y_and_46_enex5 ) begin
      reg_act_regs_data_0_8_1_enexo_2 <= act_regs_data_and_2683_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_8_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2685_enex5 | Tanh_for_y_and_46_enex5 ) begin
      reg_act_regs_data_0_8_3_enexo_2 <= act_regs_data_and_2685_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_8_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2600_enex5 | Tanh_for_y_and_46_enex5 ) begin
      reg_act_regs_data_2_8_2_enexo_2 <= act_regs_data_and_2600_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_8_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2551_enex5 | Tanh_for_y_and_46_enex5 ) begin
      reg_act_regs_data_3_8_1_enexo_2 <= act_regs_data_and_2551_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_8_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2601_enex5 | Tanh_for_y_and_46_enex5 ) begin
      reg_act_regs_data_2_8_3_enexo_2 <= act_regs_data_and_2601_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_8_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2552_enex5 | Tanh_for_y_and_46_enex5 ) begin
      reg_act_regs_data_3_8_2_enexo_2 <= act_regs_data_and_2552_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_8_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2647_enex5 | Tanh_for_y_and_46_enex5 ) begin
      reg_act_regs_data_1_8_1_enexo_2 <= act_regs_data_and_2647_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_8_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2649_enex5 | Tanh_for_y_and_46_enex5 ) begin
      reg_act_regs_data_1_8_3_enexo_2 <= act_regs_data_and_2649_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_8_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2553_enex5 | Tanh_for_y_and_46_enex5 ) begin
      reg_act_regs_data_3_8_3_enexo_2 <= act_regs_data_and_2553_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_64 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Tanh_for_y_and_47_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_64 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_64 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Tanh_for_y_and_47_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_64 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_64 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Tanh_for_y_and_47_enex5 ) begin
      reg_act_config_inst_counter_enexo_64 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_7_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2688_enex5 | Tanh_for_y_and_47_enex5 ) begin
      reg_act_regs_data_0_7_3_enexo_1 <= act_regs_data_and_2688_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_7_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2652_enex5 | Tanh_for_y_and_47_enex5 ) begin
      reg_act_regs_data_1_7_3_enexo_1 <= act_regs_data_and_2652_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_7_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2556_enex5 | Tanh_for_y_and_47_enex5 ) begin
      reg_act_regs_data_3_7_3_enexo_1 <= act_regs_data_and_2556_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_7_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Tanh_for_y_and_47_enex5 ) begin
      reg_act_regs_data_1_7_enexo <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_7_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2687_enex5 | Tanh_for_y_and_47_enex5 ) begin
      reg_act_regs_data_0_7_2_enexo_1 <= act_regs_data_and_2687_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_7_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2603_enex5 | Tanh_for_y_and_47_enex5 ) begin
      reg_act_regs_data_2_7_2_enexo_1 <= act_regs_data_and_2603_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_7_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2604_enex5 | Tanh_for_y_and_47_enex5 ) begin
      reg_act_regs_data_2_7_3_enexo_1 <= act_regs_data_and_2604_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_7_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2555_enex5 | Tanh_for_y_and_47_enex5 ) begin
      reg_act_regs_data_3_7_2_enexo_1 <= act_regs_data_and_2555_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_7_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2554_enex5 | Tanh_for_y_and_47_enex5 ) begin
      reg_act_regs_data_3_7_1_enexo_1 <= act_regs_data_and_2554_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_7_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2650_enex5 | Tanh_for_y_and_47_enex5 ) begin
      reg_act_regs_data_1_7_1_enexo_1 <= act_regs_data_and_2650_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_7_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2651_enex5 | Tanh_for_y_and_47_enex5 ) begin
      reg_act_regs_data_1_7_2_enexo_1 <= act_regs_data_and_2651_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_7_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2686_enex5 | Tanh_for_y_and_47_enex5 ) begin
      reg_act_regs_data_0_7_1_enexo_1 <= act_regs_data_and_2686_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_7_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2602_enex5 | Tanh_for_y_and_47_enex5 ) begin
      reg_act_regs_data_2_7_1_enexo_1 <= act_regs_data_and_2602_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_65 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Tanh_for_y_and_48_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_65 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_65 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Tanh_for_y_and_48_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_65 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_65 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Tanh_for_y_and_48_enex5 ) begin
      reg_act_config_inst_counter_enexo_65 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_7_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2688_enex5 | Tanh_for_y_and_48_enex5 ) begin
      reg_act_regs_data_0_7_3_enexo_2 <= act_regs_data_and_2688_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_7_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2652_enex5 | Tanh_for_y_and_48_enex5 ) begin
      reg_act_regs_data_1_7_3_enexo_2 <= act_regs_data_and_2652_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_7_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2556_enex5 | Tanh_for_y_and_48_enex5 ) begin
      reg_act_regs_data_3_7_3_enexo_2 <= act_regs_data_and_2556_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_7_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Tanh_for_y_and_48_enex5 ) begin
      reg_act_regs_data_1_7_enexo_1 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_7_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2687_enex5 | Tanh_for_y_and_48_enex5 ) begin
      reg_act_regs_data_0_7_2_enexo_2 <= act_regs_data_and_2687_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_7_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2603_enex5 | Tanh_for_y_and_48_enex5 ) begin
      reg_act_regs_data_2_7_2_enexo_2 <= act_regs_data_and_2603_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_7_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2604_enex5 | Tanh_for_y_and_48_enex5 ) begin
      reg_act_regs_data_2_7_3_enexo_2 <= act_regs_data_and_2604_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_7_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2555_enex5 | Tanh_for_y_and_48_enex5 ) begin
      reg_act_regs_data_3_7_2_enexo_2 <= act_regs_data_and_2555_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_7_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2554_enex5 | Tanh_for_y_and_48_enex5 ) begin
      reg_act_regs_data_3_7_1_enexo_2 <= act_regs_data_and_2554_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_7_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2650_enex5 | Tanh_for_y_and_48_enex5 ) begin
      reg_act_regs_data_1_7_1_enexo_2 <= act_regs_data_and_2650_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_7_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2651_enex5 | Tanh_for_y_and_48_enex5 ) begin
      reg_act_regs_data_1_7_2_enexo_2 <= act_regs_data_and_2651_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_7_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2686_enex5 | Tanh_for_y_and_48_enex5 ) begin
      reg_act_regs_data_0_7_1_enexo_2 <= act_regs_data_and_2686_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_7_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2602_enex5 | Tanh_for_y_and_48_enex5 ) begin
      reg_act_regs_data_2_7_1_enexo_2 <= act_regs_data_and_2602_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_66 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Tanh_for_y_and_49_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_66 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_66 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Tanh_for_y_and_49_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_66 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_66 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Tanh_for_y_and_49_enex5 ) begin
      reg_act_config_inst_counter_enexo_66 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_6_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2557_enex5 | Tanh_for_y_and_49_enex5 ) begin
      reg_act_regs_data_3_6_1_enexo_1 <= act_regs_data_and_2557_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_6_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2653_enex5 | Tanh_for_y_and_49_enex5 ) begin
      reg_act_regs_data_1_6_1_enexo_1 <= act_regs_data_and_2653_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_6_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2607_enex5 | Tanh_for_y_and_49_enex5 ) begin
      reg_act_regs_data_2_6_3_enexo_1 <= act_regs_data_and_2607_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_6_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2559_enex5 | Tanh_for_y_and_49_enex5 ) begin
      reg_act_regs_data_3_6_3_enexo_1 <= act_regs_data_and_2559_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_6_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Tanh_for_y_and_49_enex5 ) begin
      reg_act_regs_data_3_6_enexo <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_6_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2605_enex5 | Tanh_for_y_and_49_enex5 ) begin
      reg_act_regs_data_2_6_1_enexo_1 <= act_regs_data_and_2605_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_6_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2606_enex5 | Tanh_for_y_and_49_enex5 ) begin
      reg_act_regs_data_2_6_2_enexo_1 <= act_regs_data_and_2606_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_6_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2691_enex5 | Tanh_for_y_and_49_enex5 ) begin
      reg_act_regs_data_0_6_3_enexo_1 <= act_regs_data_and_2691_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_6_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2655_enex5 | Tanh_for_y_and_49_enex5 ) begin
      reg_act_regs_data_1_6_3_enexo_1 <= act_regs_data_and_2655_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_6_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2654_enex5 | Tanh_for_y_and_49_enex5 ) begin
      reg_act_regs_data_1_6_2_enexo_1 <= act_regs_data_and_2654_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_6_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2689_enex5 | Tanh_for_y_and_49_enex5 ) begin
      reg_act_regs_data_0_6_1_enexo_1 <= act_regs_data_and_2689_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_6_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2558_enex5 | Tanh_for_y_and_49_enex5 ) begin
      reg_act_regs_data_3_6_2_enexo_1 <= act_regs_data_and_2558_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_6_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2690_enex5 | Tanh_for_y_and_49_enex5 ) begin
      reg_act_regs_data_0_6_2_enexo_1 <= act_regs_data_and_2690_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_67 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Tanh_for_y_and_50_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_67 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_67 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Tanh_for_y_and_50_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_67 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_67 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Tanh_for_y_and_50_enex5 ) begin
      reg_act_config_inst_counter_enexo_67 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_6_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2557_enex5 | Tanh_for_y_and_50_enex5 ) begin
      reg_act_regs_data_3_6_1_enexo_2 <= act_regs_data_and_2557_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_6_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2653_enex5 | Tanh_for_y_and_50_enex5 ) begin
      reg_act_regs_data_1_6_1_enexo_2 <= act_regs_data_and_2653_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_6_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2607_enex5 | Tanh_for_y_and_50_enex5 ) begin
      reg_act_regs_data_2_6_3_enexo_2 <= act_regs_data_and_2607_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_6_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2559_enex5 | Tanh_for_y_and_50_enex5 ) begin
      reg_act_regs_data_3_6_3_enexo_2 <= act_regs_data_and_2559_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_6_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Tanh_for_y_and_50_enex5 ) begin
      reg_act_regs_data_3_6_enexo_1 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_6_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2605_enex5 | Tanh_for_y_and_50_enex5 ) begin
      reg_act_regs_data_2_6_1_enexo_2 <= act_regs_data_and_2605_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_6_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2606_enex5 | Tanh_for_y_and_50_enex5 ) begin
      reg_act_regs_data_2_6_2_enexo_2 <= act_regs_data_and_2606_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_6_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2691_enex5 | Tanh_for_y_and_50_enex5 ) begin
      reg_act_regs_data_0_6_3_enexo_2 <= act_regs_data_and_2691_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_6_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2655_enex5 | Tanh_for_y_and_50_enex5 ) begin
      reg_act_regs_data_1_6_3_enexo_2 <= act_regs_data_and_2655_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_6_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2654_enex5 | Tanh_for_y_and_50_enex5 ) begin
      reg_act_regs_data_1_6_2_enexo_2 <= act_regs_data_and_2654_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_6_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2689_enex5 | Tanh_for_y_and_50_enex5 ) begin
      reg_act_regs_data_0_6_1_enexo_2 <= act_regs_data_and_2689_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_6_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2558_enex5 | Tanh_for_y_and_50_enex5 ) begin
      reg_act_regs_data_3_6_2_enexo_2 <= act_regs_data_and_2558_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_6_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2690_enex5 | Tanh_for_y_and_50_enex5 ) begin
      reg_act_regs_data_0_6_2_enexo_2 <= act_regs_data_and_2690_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_68 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Tanh_for_y_and_51_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_68 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_68 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Tanh_for_y_and_51_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_68 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_5_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2694_enex5 | Tanh_for_y_and_51_enex5 ) begin
      reg_act_regs_data_0_5_3_enexo_1 <= act_regs_data_and_2694_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_68 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Tanh_for_y_and_51_enex5 ) begin
      reg_act_config_inst_counter_enexo_68 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_5_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2609_enex5 | Tanh_for_y_and_51_enex5 ) begin
      reg_act_regs_data_2_5_2_enexo_1 <= act_regs_data_and_2609_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_5_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2560_enex5 | Tanh_for_y_and_51_enex5 ) begin
      reg_act_regs_data_3_5_1_enexo_1 <= act_regs_data_and_2560_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_5_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2692_enex5 | Tanh_for_y_and_51_enex5 ) begin
      reg_act_regs_data_0_5_1_enexo_1 <= act_regs_data_and_2692_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_5_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Tanh_for_y_and_51_enex5 ) begin
      reg_act_regs_data_1_5_enexo <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_5_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2656_enex5 | Tanh_for_y_and_51_enex5 ) begin
      reg_act_regs_data_1_5_1_enexo_1 <= act_regs_data_and_2656_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_5_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2657_enex5 | Tanh_for_y_and_51_enex5 ) begin
      reg_act_regs_data_1_5_2_enexo_1 <= act_regs_data_and_2657_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_5_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2561_enex5 | Tanh_for_y_and_51_enex5 ) begin
      reg_act_regs_data_3_5_2_enexo_1 <= act_regs_data_and_2561_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_5_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2693_enex5 | Tanh_for_y_and_51_enex5 ) begin
      reg_act_regs_data_0_5_2_enexo_1 <= act_regs_data_and_2693_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_5_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2658_enex5 | Tanh_for_y_and_51_enex5 ) begin
      reg_act_regs_data_1_5_3_enexo_1 <= act_regs_data_and_2658_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_5_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2562_enex5 | Tanh_for_y_and_51_enex5 ) begin
      reg_act_regs_data_3_5_3_enexo_1 <= act_regs_data_and_2562_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_5_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2608_enex5 | Tanh_for_y_and_51_enex5 ) begin
      reg_act_regs_data_2_5_1_enexo_1 <= act_regs_data_and_2608_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_5_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2610_enex5 | Tanh_for_y_and_51_enex5 ) begin
      reg_act_regs_data_2_5_3_enexo_1 <= act_regs_data_and_2610_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_69 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Tanh_for_y_and_52_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_69 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_69 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Tanh_for_y_and_52_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_69 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_5_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2694_enex5 | Tanh_for_y_and_52_enex5 ) begin
      reg_act_regs_data_0_5_3_enexo_2 <= act_regs_data_and_2694_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_69 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Tanh_for_y_and_52_enex5 ) begin
      reg_act_config_inst_counter_enexo_69 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_5_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2609_enex5 | Tanh_for_y_and_52_enex5 ) begin
      reg_act_regs_data_2_5_2_enexo_2 <= act_regs_data_and_2609_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_5_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2560_enex5 | Tanh_for_y_and_52_enex5 ) begin
      reg_act_regs_data_3_5_1_enexo_2 <= act_regs_data_and_2560_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_5_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2692_enex5 | Tanh_for_y_and_52_enex5 ) begin
      reg_act_regs_data_0_5_1_enexo_2 <= act_regs_data_and_2692_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_5_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Tanh_for_y_and_52_enex5 ) begin
      reg_act_regs_data_1_5_enexo_1 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_5_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2656_enex5 | Tanh_for_y_and_52_enex5 ) begin
      reg_act_regs_data_1_5_1_enexo_2 <= act_regs_data_and_2656_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_5_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2657_enex5 | Tanh_for_y_and_52_enex5 ) begin
      reg_act_regs_data_1_5_2_enexo_2 <= act_regs_data_and_2657_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_5_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2561_enex5 | Tanh_for_y_and_52_enex5 ) begin
      reg_act_regs_data_3_5_2_enexo_2 <= act_regs_data_and_2561_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_5_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2693_enex5 | Tanh_for_y_and_52_enex5 ) begin
      reg_act_regs_data_0_5_2_enexo_2 <= act_regs_data_and_2693_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_5_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2658_enex5 | Tanh_for_y_and_52_enex5 ) begin
      reg_act_regs_data_1_5_3_enexo_2 <= act_regs_data_and_2658_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_5_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2562_enex5 | Tanh_for_y_and_52_enex5 ) begin
      reg_act_regs_data_3_5_3_enexo_2 <= act_regs_data_and_2562_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_5_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2608_enex5 | Tanh_for_y_and_52_enex5 ) begin
      reg_act_regs_data_2_5_1_enexo_2 <= act_regs_data_and_2608_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_5_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2610_enex5 | Tanh_for_y_and_52_enex5 ) begin
      reg_act_regs_data_2_5_3_enexo_2 <= act_regs_data_and_2610_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_70 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Tanh_for_y_and_53_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_70 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_70 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Tanh_for_y_and_53_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_70 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_70 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Tanh_for_y_and_53_enex5 ) begin
      reg_act_config_inst_counter_enexo_70 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_4_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2697_enex5 | Tanh_for_y_and_53_enex5 ) begin
      reg_act_regs_data_0_4_3_enexo_1 <= act_regs_data_and_2697_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_4_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2563_enex5 | Tanh_for_y_and_53_enex5 ) begin
      reg_act_regs_data_3_4_1_enexo_1 <= act_regs_data_and_2563_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_4_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2564_enex5 | Tanh_for_y_and_53_enex5 ) begin
      reg_act_regs_data_3_4_2_enexo_1 <= act_regs_data_and_2564_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_4_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2661_enex5 | Tanh_for_y_and_53_enex5 ) begin
      reg_act_regs_data_1_4_3_enexo_1 <= act_regs_data_and_2661_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_4_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2695_enex5 | Tanh_for_y_and_53_enex5 ) begin
      reg_act_regs_data_0_4_1_enexo_1 <= act_regs_data_and_2695_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_4_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2611_enex5 | Tanh_for_y_and_53_enex5 ) begin
      reg_act_regs_data_2_4_1_enexo_1 <= act_regs_data_and_2611_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_4_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2565_enex5 | Tanh_for_y_and_53_enex5 ) begin
      reg_act_regs_data_3_4_3_enexo_1 <= act_regs_data_and_2565_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_4_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2660_enex5 | Tanh_for_y_and_53_enex5 ) begin
      reg_act_regs_data_1_4_2_enexo_1 <= act_regs_data_and_2660_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_4_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Tanh_for_y_and_53_enex5 ) begin
      reg_act_regs_data_3_4_enexo <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_4_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2613_enex5 | Tanh_for_y_and_53_enex5 ) begin
      reg_act_regs_data_2_4_3_enexo_1 <= act_regs_data_and_2613_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_4_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2659_enex5 | Tanh_for_y_and_53_enex5 ) begin
      reg_act_regs_data_1_4_1_enexo_1 <= act_regs_data_and_2659_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_4_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2696_enex5 | Tanh_for_y_and_53_enex5 ) begin
      reg_act_regs_data_0_4_2_enexo_1 <= act_regs_data_and_2696_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_4_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2612_enex5 | Tanh_for_y_and_53_enex5 ) begin
      reg_act_regs_data_2_4_2_enexo_1 <= act_regs_data_and_2612_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_71 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Tanh_for_y_and_54_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_71 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_71 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Tanh_for_y_and_54_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_71 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_71 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Tanh_for_y_and_54_enex5 ) begin
      reg_act_config_inst_counter_enexo_71 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_4_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2697_enex5 | Tanh_for_y_and_54_enex5 ) begin
      reg_act_regs_data_0_4_3_enexo_2 <= act_regs_data_and_2697_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_4_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2563_enex5 | Tanh_for_y_and_54_enex5 ) begin
      reg_act_regs_data_3_4_1_enexo_2 <= act_regs_data_and_2563_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_4_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2564_enex5 | Tanh_for_y_and_54_enex5 ) begin
      reg_act_regs_data_3_4_2_enexo_2 <= act_regs_data_and_2564_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_4_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2661_enex5 | Tanh_for_y_and_54_enex5 ) begin
      reg_act_regs_data_1_4_3_enexo_2 <= act_regs_data_and_2661_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_4_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2695_enex5 | Tanh_for_y_and_54_enex5 ) begin
      reg_act_regs_data_0_4_1_enexo_2 <= act_regs_data_and_2695_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_4_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2611_enex5 | Tanh_for_y_and_54_enex5 ) begin
      reg_act_regs_data_2_4_1_enexo_2 <= act_regs_data_and_2611_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_4_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2565_enex5 | Tanh_for_y_and_54_enex5 ) begin
      reg_act_regs_data_3_4_3_enexo_2 <= act_regs_data_and_2565_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_4_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2660_enex5 | Tanh_for_y_and_54_enex5 ) begin
      reg_act_regs_data_1_4_2_enexo_2 <= act_regs_data_and_2660_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_4_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Tanh_for_y_and_54_enex5 ) begin
      reg_act_regs_data_3_4_enexo_1 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_4_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2613_enex5 | Tanh_for_y_and_54_enex5 ) begin
      reg_act_regs_data_2_4_3_enexo_2 <= act_regs_data_and_2613_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_4_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2659_enex5 | Tanh_for_y_and_54_enex5 ) begin
      reg_act_regs_data_1_4_1_enexo_2 <= act_regs_data_and_2659_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_4_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2696_enex5 | Tanh_for_y_and_54_enex5 ) begin
      reg_act_regs_data_0_4_2_enexo_2 <= act_regs_data_and_2696_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_4_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2612_enex5 | Tanh_for_y_and_54_enex5 ) begin
      reg_act_regs_data_2_4_2_enexo_2 <= act_regs_data_and_2612_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_72 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Tanh_for_y_and_55_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_72 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_72 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Tanh_for_y_and_55_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_72 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_72 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Tanh_for_y_and_55_enex5 ) begin
      reg_act_config_inst_counter_enexo_72 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_3_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2700_enex5 | Tanh_for_y_and_55_enex5 ) begin
      reg_act_regs_data_0_3_3_enexo_1 <= act_regs_data_and_2700_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_3_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2568_enex5 | Tanh_for_y_and_55_enex5 ) begin
      reg_act_regs_data_3_3_3_enexo_1 <= act_regs_data_and_2568_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_3_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2698_enex5 | Tanh_for_y_and_55_enex5 ) begin
      reg_act_regs_data_0_3_1_enexo_1 <= act_regs_data_and_2698_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_3_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Tanh_for_y_and_55_enex5 ) begin
      reg_act_regs_data_3_3_enexo <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_3_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2566_enex5 | Tanh_for_y_and_55_enex5 ) begin
      reg_act_regs_data_3_3_1_enexo_1 <= act_regs_data_and_2566_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_3_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2662_enex5 | Tanh_for_y_and_55_enex5 ) begin
      reg_act_regs_data_1_3_1_enexo_1 <= act_regs_data_and_2662_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_3_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2699_enex5 | Tanh_for_y_and_55_enex5 ) begin
      reg_act_regs_data_0_3_2_enexo_1 <= act_regs_data_and_2699_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_3_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2664_enex5 | Tanh_for_y_and_55_enex5 ) begin
      reg_act_regs_data_1_3_3_enexo_1 <= act_regs_data_and_2664_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_3_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2663_enex5 | Tanh_for_y_and_55_enex5 ) begin
      reg_act_regs_data_1_3_2_enexo_1 <= act_regs_data_and_2663_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_3_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2567_enex5 | Tanh_for_y_and_55_enex5 ) begin
      reg_act_regs_data_3_3_2_enexo_1 <= act_regs_data_and_2567_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_3_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2614_enex5 | Tanh_for_y_and_55_enex5 ) begin
      reg_act_regs_data_2_3_1_enexo_1 <= act_regs_data_and_2614_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_3_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2616_enex5 | Tanh_for_y_and_55_enex5 ) begin
      reg_act_regs_data_2_3_3_enexo_1 <= act_regs_data_and_2616_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_3_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2615_enex5 | Tanh_for_y_and_55_enex5 ) begin
      reg_act_regs_data_2_3_2_enexo_1 <= act_regs_data_and_2615_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_73 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Tanh_for_y_and_56_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_73 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_73 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Tanh_for_y_and_56_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_73 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_73 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Tanh_for_y_and_56_enex5 ) begin
      reg_act_config_inst_counter_enexo_73 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_3_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2700_enex5 | Tanh_for_y_and_56_enex5 ) begin
      reg_act_regs_data_0_3_3_enexo_2 <= act_regs_data_and_2700_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_3_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2568_enex5 | Tanh_for_y_and_56_enex5 ) begin
      reg_act_regs_data_3_3_3_enexo_2 <= act_regs_data_and_2568_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_3_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2698_enex5 | Tanh_for_y_and_56_enex5 ) begin
      reg_act_regs_data_0_3_1_enexo_2 <= act_regs_data_and_2698_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Tanh_for_y_and_56_enex5 ) begin
      reg_act_regs_data_3_3_enexo_1 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_3_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2566_enex5 | Tanh_for_y_and_56_enex5 ) begin
      reg_act_regs_data_3_3_1_enexo_2 <= act_regs_data_and_2566_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_3_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2662_enex5 | Tanh_for_y_and_56_enex5 ) begin
      reg_act_regs_data_1_3_1_enexo_2 <= act_regs_data_and_2662_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_3_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2699_enex5 | Tanh_for_y_and_56_enex5 ) begin
      reg_act_regs_data_0_3_2_enexo_2 <= act_regs_data_and_2699_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_3_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2664_enex5 | Tanh_for_y_and_56_enex5 ) begin
      reg_act_regs_data_1_3_3_enexo_2 <= act_regs_data_and_2664_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_3_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2663_enex5 | Tanh_for_y_and_56_enex5 ) begin
      reg_act_regs_data_1_3_2_enexo_2 <= act_regs_data_and_2663_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_3_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2567_enex5 | Tanh_for_y_and_56_enex5 ) begin
      reg_act_regs_data_3_3_2_enexo_2 <= act_regs_data_and_2567_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_3_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2614_enex5 | Tanh_for_y_and_56_enex5 ) begin
      reg_act_regs_data_2_3_1_enexo_2 <= act_regs_data_and_2614_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_3_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2616_enex5 | Tanh_for_y_and_56_enex5 ) begin
      reg_act_regs_data_2_3_3_enexo_2 <= act_regs_data_and_2616_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_3_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2615_enex5 | Tanh_for_y_and_56_enex5 ) begin
      reg_act_regs_data_2_3_2_enexo_2 <= act_regs_data_and_2615_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_2_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2617_enex5 | Tanh_for_y_and_57_enex5 ) begin
      reg_act_regs_data_2_2_1_enexo_1 <= act_regs_data_and_2617_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_74 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Tanh_for_y_and_57_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_74 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_74 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Tanh_for_y_and_57_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_74 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_74 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Tanh_for_y_and_57_enex5 ) begin
      reg_act_config_inst_counter_enexo_74 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_2_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Tanh_for_y_and_57_enex5 ) begin
      reg_act_regs_data_3_2_enexo <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_2_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2702_enex5 | Tanh_for_y_and_57_enex5 ) begin
      reg_act_regs_data_0_2_2_enexo_1 <= act_regs_data_and_2702_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_2_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2569_enex5 | Tanh_for_y_and_57_enex5 ) begin
      reg_act_regs_data_3_2_1_enexo_1 <= act_regs_data_and_2569_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_2_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2571_enex5 | Tanh_for_y_and_57_enex5 ) begin
      reg_act_regs_data_3_2_3_enexo_1 <= act_regs_data_and_2571_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_2_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2619_enex5 | Tanh_for_y_and_57_enex5 ) begin
      reg_act_regs_data_2_2_3_enexo_1 <= act_regs_data_and_2619_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_2_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2665_enex5 | Tanh_for_y_and_57_enex5 ) begin
      reg_act_regs_data_1_2_1_enexo_1 <= act_regs_data_and_2665_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_2_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2666_enex5 | Tanh_for_y_and_57_enex5 ) begin
      reg_act_regs_data_1_2_2_enexo_1 <= act_regs_data_and_2666_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_2_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2570_enex5 | Tanh_for_y_and_57_enex5 ) begin
      reg_act_regs_data_3_2_2_enexo_1 <= act_regs_data_and_2570_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_2_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2618_enex5 | Tanh_for_y_and_57_enex5 ) begin
      reg_act_regs_data_2_2_2_enexo_1 <= act_regs_data_and_2618_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_2_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2703_enex5 | Tanh_for_y_and_57_enex5 ) begin
      reg_act_regs_data_0_2_3_enexo_1 <= act_regs_data_and_2703_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_2_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2701_enex5 | Tanh_for_y_and_57_enex5 ) begin
      reg_act_regs_data_0_2_1_enexo_1 <= act_regs_data_and_2701_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_2_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2667_enex5 | Tanh_for_y_and_57_enex5 ) begin
      reg_act_regs_data_1_2_3_enexo_1 <= act_regs_data_and_2667_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_2_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2617_enex5 | Tanh_for_y_and_58_enex5 ) begin
      reg_act_regs_data_2_2_1_enexo_2 <= act_regs_data_and_2617_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_75 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Tanh_for_y_and_58_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_75 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_75 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Tanh_for_y_and_58_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_75 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_75 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Tanh_for_y_and_58_enex5 ) begin
      reg_act_config_inst_counter_enexo_75 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Tanh_for_y_and_58_enex5 ) begin
      reg_act_regs_data_3_2_enexo_1 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_2_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2702_enex5 | Tanh_for_y_and_58_enex5 ) begin
      reg_act_regs_data_0_2_2_enexo_2 <= act_regs_data_and_2702_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_2_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2569_enex5 | Tanh_for_y_and_58_enex5 ) begin
      reg_act_regs_data_3_2_1_enexo_2 <= act_regs_data_and_2569_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_2_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2571_enex5 | Tanh_for_y_and_58_enex5 ) begin
      reg_act_regs_data_3_2_3_enexo_2 <= act_regs_data_and_2571_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_2_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2619_enex5 | Tanh_for_y_and_58_enex5 ) begin
      reg_act_regs_data_2_2_3_enexo_2 <= act_regs_data_and_2619_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_2_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2665_enex5 | Tanh_for_y_and_58_enex5 ) begin
      reg_act_regs_data_1_2_1_enexo_2 <= act_regs_data_and_2665_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_2_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2666_enex5 | Tanh_for_y_and_58_enex5 ) begin
      reg_act_regs_data_1_2_2_enexo_2 <= act_regs_data_and_2666_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_2_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2570_enex5 | Tanh_for_y_and_58_enex5 ) begin
      reg_act_regs_data_3_2_2_enexo_2 <= act_regs_data_and_2570_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_2_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2618_enex5 | Tanh_for_y_and_58_enex5 ) begin
      reg_act_regs_data_2_2_2_enexo_2 <= act_regs_data_and_2618_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_2_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2703_enex5 | Tanh_for_y_and_58_enex5 ) begin
      reg_act_regs_data_0_2_3_enexo_2 <= act_regs_data_and_2703_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_2_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2701_enex5 | Tanh_for_y_and_58_enex5 ) begin
      reg_act_regs_data_0_2_1_enexo_2 <= act_regs_data_and_2701_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_2_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2667_enex5 | Tanh_for_y_and_58_enex5 ) begin
      reg_act_regs_data_1_2_3_enexo_2 <= act_regs_data_and_2667_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_76 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Tanh_for_y_and_59_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_76 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_76 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Tanh_for_y_and_59_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_76 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_1_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2620_enex5 | Tanh_for_y_and_59_enex5 ) begin
      reg_act_regs_data_2_1_1_enexo_1 <= act_regs_data_and_2620_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_76 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Tanh_for_y_and_59_enex5 ) begin
      reg_act_config_inst_counter_enexo_76 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_1_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2669_enex5 | Tanh_for_y_and_59_enex5 ) begin
      reg_act_regs_data_1_1_2_enexo_1 <= act_regs_data_and_2669_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_1_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2763_enex5 | Tanh_for_y_and_59_enex5 ) begin
      reg_act_regs_data_0_1_3_enexo_1 <= act_regs_data_and_2763_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_1_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2572_enex5 | Tanh_for_y_and_59_enex5 ) begin
      reg_act_regs_data_3_1_1_enexo_1 <= act_regs_data_and_2572_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_1_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Tanh_for_y_and_59_enex5 ) begin
      reg_act_regs_data_2_1_enexo <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_1_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2761_enex5 | Tanh_for_y_and_59_enex5 ) begin
      reg_act_regs_data_0_1_1_enexo_1 <= act_regs_data_and_2761_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_1_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2573_enex5 | Tanh_for_y_and_59_enex5 ) begin
      reg_act_regs_data_3_1_2_enexo_1 <= act_regs_data_and_2573_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_1_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2668_enex5 | Tanh_for_y_and_59_enex5 ) begin
      reg_act_regs_data_1_1_1_enexo_1 <= act_regs_data_and_2668_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_1_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2762_enex5 | Tanh_for_y_and_59_enex5 ) begin
      reg_act_regs_data_0_1_2_enexo_1 <= act_regs_data_and_2762_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_1_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2621_enex5 | Tanh_for_y_and_59_enex5 ) begin
      reg_act_regs_data_2_1_2_enexo_1 <= act_regs_data_and_2621_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_1_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2574_enex5 | Tanh_for_y_and_59_enex5 ) begin
      reg_act_regs_data_3_1_3_enexo_1 <= act_regs_data_and_2574_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_1_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2670_enex5 | Tanh_for_y_and_59_enex5 ) begin
      reg_act_regs_data_1_1_3_enexo_1 <= act_regs_data_and_2670_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_1_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2622_enex5 | Tanh_for_y_and_59_enex5 ) begin
      reg_act_regs_data_2_1_3_enexo_1 <= act_regs_data_and_2622_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_77 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Tanh_for_y_and_60_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_77 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_77 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Tanh_for_y_and_60_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_77 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_1_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2620_enex5 | Tanh_for_y_and_60_enex5 ) begin
      reg_act_regs_data_2_1_1_enexo_2 <= act_regs_data_and_2620_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_77 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Tanh_for_y_and_60_enex5 ) begin
      reg_act_config_inst_counter_enexo_77 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_1_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2669_enex5 | Tanh_for_y_and_60_enex5 ) begin
      reg_act_regs_data_1_1_2_enexo_2 <= act_regs_data_and_2669_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_1_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2763_enex5 | Tanh_for_y_and_60_enex5 ) begin
      reg_act_regs_data_0_1_3_enexo_2 <= act_regs_data_and_2763_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_1_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2572_enex5 | Tanh_for_y_and_60_enex5 ) begin
      reg_act_regs_data_3_1_1_enexo_2 <= act_regs_data_and_2572_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Tanh_for_y_and_60_enex5 ) begin
      reg_act_regs_data_2_1_enexo_1 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_1_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2761_enex5 | Tanh_for_y_and_60_enex5 ) begin
      reg_act_regs_data_0_1_1_enexo_2 <= act_regs_data_and_2761_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_1_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2573_enex5 | Tanh_for_y_and_60_enex5 ) begin
      reg_act_regs_data_3_1_2_enexo_2 <= act_regs_data_and_2573_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_1_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2668_enex5 | Tanh_for_y_and_60_enex5 ) begin
      reg_act_regs_data_1_1_1_enexo_2 <= act_regs_data_and_2668_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_1_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2762_enex5 | Tanh_for_y_and_60_enex5 ) begin
      reg_act_regs_data_0_1_2_enexo_2 <= act_regs_data_and_2762_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_1_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2621_enex5 | Tanh_for_y_and_60_enex5 ) begin
      reg_act_regs_data_2_1_2_enexo_2 <= act_regs_data_and_2621_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_1_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2574_enex5 | Tanh_for_y_and_60_enex5 ) begin
      reg_act_regs_data_3_1_3_enexo_2 <= act_regs_data_and_2574_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_1_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2670_enex5 | Tanh_for_y_and_60_enex5 ) begin
      reg_act_regs_data_1_1_3_enexo_2 <= act_regs_data_and_2670_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_1_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2622_enex5 | Tanh_for_y_and_60_enex5 ) begin
      reg_act_regs_data_2_1_3_enexo_2 <= act_regs_data_and_2622_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_78 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Tanh_for_y_and_61_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_78 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_0_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2575_enex5 | Tanh_for_y_and_61_enex5 ) begin
      reg_act_regs_data_3_0_1_enexo_1 <= act_regs_data_and_2575_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_0_enexo <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Tanh_for_y_and_61_enex5 ) begin
      reg_act_regs_data_3_0_enexo <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_78 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Tanh_for_y_and_61_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_78 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_78 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Tanh_for_y_and_61_enex5 ) begin
      reg_act_config_inst_counter_enexo_78 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_0_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2577_enex5 | Tanh_for_y_and_61_enex5 ) begin
      reg_act_regs_data_3_0_3_enexo_1 <= act_regs_data_and_2577_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_0_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2766_enex5 | Tanh_for_y_and_61_enex5 ) begin
      reg_act_regs_data_0_0_3_enexo_1 <= act_regs_data_and_2766_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_0_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2764_enex5 | Tanh_for_y_and_61_enex5 ) begin
      reg_act_regs_data_0_0_1_enexo_1 <= act_regs_data_and_2764_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_0_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2576_enex5 | Tanh_for_y_and_61_enex5 ) begin
      reg_act_regs_data_3_0_2_enexo_1 <= act_regs_data_and_2576_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_0_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2623_enex5 | Tanh_for_y_and_61_enex5 ) begin
      reg_act_regs_data_2_0_1_enexo_1 <= act_regs_data_and_2623_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_0_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2765_enex5 | Tanh_for_y_and_61_enex5 ) begin
      reg_act_regs_data_0_0_2_enexo_1 <= act_regs_data_and_2765_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_0_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2672_enex5 | Tanh_for_y_and_61_enex5 ) begin
      reg_act_regs_data_1_0_2_enexo_1 <= act_regs_data_and_2672_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_0_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2625_enex5 | Tanh_for_y_and_61_enex5 ) begin
      reg_act_regs_data_2_0_3_enexo_1 <= act_regs_data_and_2625_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_0_1_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2671_enex5 | Tanh_for_y_and_61_enex5 ) begin
      reg_act_regs_data_1_0_1_enexo_1 <= act_regs_data_and_2671_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_0_2_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2624_enex5 | Tanh_for_y_and_61_enex5 ) begin
      reg_act_regs_data_2_0_2_enexo_1 <= act_regs_data_and_2624_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_0_3_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_2673_enex5 | Tanh_for_y_and_61_enex5 ) begin
      reg_act_regs_data_1_0_3_enexo_1 <= act_regs_data_and_2673_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_79 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Tanh_for_y_and_62_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_79 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_0_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2575_enex5 | Tanh_for_y_and_62_enex5 ) begin
      reg_act_regs_data_3_0_1_enexo_2 <= act_regs_data_and_2575_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Tanh_for_y_and_62_enex5 ) begin
      reg_act_regs_data_3_0_enexo_1 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_79 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Tanh_for_y_and_62_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_79 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_79 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Tanh_for_y_and_62_enex5 ) begin
      reg_act_config_inst_counter_enexo_79 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_0_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2577_enex5 | Tanh_for_y_and_62_enex5 ) begin
      reg_act_regs_data_3_0_3_enexo_2 <= act_regs_data_and_2577_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_0_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2766_enex5 | Tanh_for_y_and_62_enex5 ) begin
      reg_act_regs_data_0_0_3_enexo_2 <= act_regs_data_and_2766_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_0_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2764_enex5 | Tanh_for_y_and_62_enex5 ) begin
      reg_act_regs_data_0_0_1_enexo_2 <= act_regs_data_and_2764_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_0_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2576_enex5 | Tanh_for_y_and_62_enex5 ) begin
      reg_act_regs_data_3_0_2_enexo_2 <= act_regs_data_and_2576_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_0_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2623_enex5 | Tanh_for_y_and_62_enex5 ) begin
      reg_act_regs_data_2_0_1_enexo_2 <= act_regs_data_and_2623_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_0_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2765_enex5 | Tanh_for_y_and_62_enex5 ) begin
      reg_act_regs_data_0_0_2_enexo_2 <= act_regs_data_and_2765_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_0_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2672_enex5 | Tanh_for_y_and_62_enex5 ) begin
      reg_act_regs_data_1_0_2_enexo_2 <= act_regs_data_and_2672_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_0_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2625_enex5 | Tanh_for_y_and_62_enex5 ) begin
      reg_act_regs_data_2_0_3_enexo_2 <= act_regs_data_and_2625_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_0_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2671_enex5 | Tanh_for_y_and_62_enex5 ) begin
      reg_act_regs_data_1_0_1_enexo_2 <= act_regs_data_and_2671_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_0_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2624_enex5 | Tanh_for_y_and_62_enex5 ) begin
      reg_act_regs_data_2_0_2_enexo_2 <= act_regs_data_and_2624_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_0_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_2673_enex5 | Tanh_for_y_and_62_enex5 ) begin
      reg_act_regs_data_1_0_3_enexo_2 <= act_regs_data_and_2673_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_80 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_31_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_80 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_80 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_31_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_80 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_80 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_31_enex5 ) begin
      reg_act_config_inst_counter_enexo_80 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_15_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_31_enex5 ) begin
      reg_act_regs_data_1_15_enexo_2 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_15_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2674_enex5 | Relu_for_y_qelse_and_31_enex5 ) begin
      reg_act_regs_data_0_15_1_enexo_3 <= act_regs_data_and_2674_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_15_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2626_enex5 | Relu_for_y_qelse_and_31_enex5 ) begin
      reg_act_regs_data_1_15_1_enexo_3 <= act_regs_data_and_2626_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_15_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2578_enex5 | Relu_for_y_qelse_and_31_enex5 ) begin
      reg_act_regs_data_2_15_1_enexo_3 <= act_regs_data_and_2578_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_15_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2530_enex5 | Relu_for_y_qelse_and_31_enex5 ) begin
      reg_act_regs_data_3_15_1_enexo_3 <= act_regs_data_and_2530_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_81 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_32_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_81 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_81 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_32_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_81 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_81 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_32_enex5 ) begin
      reg_act_config_inst_counter_enexo_81 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_15_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_32_enex5 ) begin
      reg_act_regs_data_1_15_enexo_3 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_15_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2531_enex5 | Relu_for_y_qelse_and_32_enex5 ) begin
      reg_act_regs_data_3_15_2_enexo_3 <= act_regs_data_and_2531_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_15_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2579_enex5 | Relu_for_y_qelse_and_32_enex5 ) begin
      reg_act_regs_data_2_15_2_enexo_3 <= act_regs_data_and_2579_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_15_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2675_enex5 | Relu_for_y_qelse_and_32_enex5 ) begin
      reg_act_regs_data_0_15_2_enexo_3 <= act_regs_data_and_2675_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_15_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2627_enex5 | Relu_for_y_qelse_and_32_enex5 ) begin
      reg_act_regs_data_1_15_2_enexo_3 <= act_regs_data_and_2627_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_82 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_33_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_82 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_82 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_33_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_82 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_15_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2580_enex5 | Relu_for_y_qelse_and_33_enex5 ) begin
      reg_act_regs_data_2_15_3_enexo_3 <= act_regs_data_and_2580_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_82 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_33_enex5 ) begin
      reg_act_config_inst_counter_enexo_82 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_15_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_33_enex5 ) begin
      reg_act_regs_data_1_15_enexo_4 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_15_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2676_enex5 | Relu_for_y_qelse_and_33_enex5 ) begin
      reg_act_regs_data_0_15_3_enexo_3 <= act_regs_data_and_2676_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_15_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2628_enex5 | Relu_for_y_qelse_and_33_enex5 ) begin
      reg_act_regs_data_1_15_3_enexo_3 <= act_regs_data_and_2628_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_15_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2532_enex5 | Relu_for_y_qelse_and_33_enex5 ) begin
      reg_act_regs_data_3_15_3_enexo_3 <= act_regs_data_and_2532_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_83 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_34_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_83 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_14_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2629_enex5 | Relu_for_y_qelse_and_34_enex5 ) begin
      reg_act_regs_data_1_14_1_enexo_3 <= act_regs_data_and_2629_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_83 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_34_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_83 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_83 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_34_enex5 ) begin
      reg_act_config_inst_counter_enexo_83 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_14_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_34_enex5 ) begin
      reg_act_regs_data_0_14_enexo_2 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_14_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2581_enex5 | Relu_for_y_qelse_and_34_enex5 ) begin
      reg_act_regs_data_2_14_1_enexo_3 <= act_regs_data_and_2581_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_14_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2533_enex5 | Relu_for_y_qelse_and_34_enex5 ) begin
      reg_act_regs_data_3_14_1_enexo_3 <= act_regs_data_and_2533_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_14_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2677_enex5 | Relu_for_y_qelse_and_34_enex5 ) begin
      reg_act_regs_data_0_14_1_enexo_3 <= act_regs_data_and_2677_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_84 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_35_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_84 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_14_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2678_enex5 | Relu_for_y_qelse_and_35_enex5 ) begin
      reg_act_regs_data_0_14_2_enexo_3 <= act_regs_data_and_2678_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_84 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_35_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_84 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_84 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_35_enex5 ) begin
      reg_act_config_inst_counter_enexo_84 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_14_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_35_enex5 ) begin
      reg_act_regs_data_0_14_enexo_3 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_14_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2582_enex5 | Relu_for_y_qelse_and_35_enex5 ) begin
      reg_act_regs_data_2_14_2_enexo_3 <= act_regs_data_and_2582_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_14_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2534_enex5 | Relu_for_y_qelse_and_35_enex5 ) begin
      reg_act_regs_data_3_14_2_enexo_3 <= act_regs_data_and_2534_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_14_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2630_enex5 | Relu_for_y_qelse_and_35_enex5 ) begin
      reg_act_regs_data_1_14_2_enexo_3 <= act_regs_data_and_2630_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_85 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_36_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_85 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_85 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_36_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_85 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_85 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_36_enex5 ) begin
      reg_act_config_inst_counter_enexo_85 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_14_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_36_enex5 ) begin
      reg_act_regs_data_0_14_enexo_4 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_14_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2679_enex5 | Relu_for_y_qelse_and_36_enex5 ) begin
      reg_act_regs_data_0_14_3_enexo_3 <= act_regs_data_and_2679_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_14_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2583_enex5 | Relu_for_y_qelse_and_36_enex5 ) begin
      reg_act_regs_data_2_14_3_enexo_3 <= act_regs_data_and_2583_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_14_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2535_enex5 | Relu_for_y_qelse_and_36_enex5 ) begin
      reg_act_regs_data_3_14_3_enexo_3 <= act_regs_data_and_2535_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_14_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2631_enex5 | Relu_for_y_qelse_and_36_enex5 ) begin
      reg_act_regs_data_1_14_3_enexo_3 <= act_regs_data_and_2631_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_86 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_37_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_86 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_13_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2632_enex5 | Relu_for_y_qelse_and_37_enex5 ) begin
      reg_act_regs_data_1_13_1_enexo_3 <= act_regs_data_and_2632_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_13_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2584_enex5 | Relu_for_y_qelse_and_37_enex5 ) begin
      reg_act_regs_data_2_13_1_enexo_3 <= act_regs_data_and_2584_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_86 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_37_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_86 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_86 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_37_enex5 ) begin
      reg_act_config_inst_counter_enexo_86 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_13_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2749_enex5 | Relu_for_y_qelse_and_37_enex5 ) begin
      reg_act_regs_data_0_13_1_enexo_3 <= act_regs_data_and_2749_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_13_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_37_enex5 ) begin
      reg_act_regs_data_3_13_enexo_2 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_13_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2536_enex5 | Relu_for_y_qelse_and_37_enex5 ) begin
      reg_act_regs_data_3_13_1_enexo_3 <= act_regs_data_and_2536_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_13_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2537_enex5 | Relu_for_y_qelse_and_38_enex5 ) begin
      reg_act_regs_data_3_13_2_enexo_3 <= act_regs_data_and_2537_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_87 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_38_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_87 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_87 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_38_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_87 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_13_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2750_enex5 | Relu_for_y_qelse_and_38_enex5 ) begin
      reg_act_regs_data_0_13_2_enexo_3 <= act_regs_data_and_2750_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_87 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_38_enex5 ) begin
      reg_act_config_inst_counter_enexo_87 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_13_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2633_enex5 | Relu_for_y_qelse_and_38_enex5 ) begin
      reg_act_regs_data_1_13_2_enexo_3 <= act_regs_data_and_2633_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_13_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_38_enex5 ) begin
      reg_act_regs_data_3_13_enexo_3 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_13_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2585_enex5 | Relu_for_y_qelse_and_38_enex5 ) begin
      reg_act_regs_data_2_13_2_enexo_3 <= act_regs_data_and_2585_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_88 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_39_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_88 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_88 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_39_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_88 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_88 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_39_enex5 ) begin
      reg_act_config_inst_counter_enexo_88 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_13_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_39_enex5 ) begin
      reg_act_regs_data_3_13_enexo_4 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_13_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2586_enex5 | Relu_for_y_qelse_and_39_enex5 ) begin
      reg_act_regs_data_2_13_3_enexo_3 <= act_regs_data_and_2586_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_13_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2538_enex5 | Relu_for_y_qelse_and_39_enex5 ) begin
      reg_act_regs_data_3_13_3_enexo_3 <= act_regs_data_and_2538_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_13_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2634_enex5 | Relu_for_y_qelse_and_39_enex5 ) begin
      reg_act_regs_data_1_13_3_enexo_3 <= act_regs_data_and_2634_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_13_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2751_enex5 | Relu_for_y_qelse_and_39_enex5 ) begin
      reg_act_regs_data_0_13_3_enexo_3 <= act_regs_data_and_2751_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_89 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_40_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_89 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_89 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_40_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_89 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_89 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_40_enex5 ) begin
      reg_act_config_inst_counter_enexo_89 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_12_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2587_enex5 | Relu_for_y_qelse_and_40_enex5 ) begin
      reg_act_regs_data_2_12_1_enexo_3 <= act_regs_data_and_2587_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_12_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_40_enex5 ) begin
      reg_act_regs_data_0_12_enexo_2 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_12_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2752_enex5 | Relu_for_y_qelse_and_40_enex5 ) begin
      reg_act_regs_data_0_12_1_enexo_3 <= act_regs_data_and_2752_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_12_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2635_enex5 | Relu_for_y_qelse_and_40_enex5 ) begin
      reg_act_regs_data_1_12_1_enexo_3 <= act_regs_data_and_2635_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_12_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2539_enex5 | Relu_for_y_qelse_and_40_enex5 ) begin
      reg_act_regs_data_3_12_1_enexo_3 <= act_regs_data_and_2539_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_90 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_41_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_90 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_90 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_41_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_90 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_12_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2588_enex5 | Relu_for_y_qelse_and_41_enex5 ) begin
      reg_act_regs_data_2_12_2_enexo_3 <= act_regs_data_and_2588_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_90 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_41_enex5 ) begin
      reg_act_config_inst_counter_enexo_90 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_12_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_41_enex5 ) begin
      reg_act_regs_data_0_12_enexo_3 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_12_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2753_enex5 | Relu_for_y_qelse_and_41_enex5 ) begin
      reg_act_regs_data_0_12_2_enexo_3 <= act_regs_data_and_2753_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_12_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2540_enex5 | Relu_for_y_qelse_and_41_enex5 ) begin
      reg_act_regs_data_3_12_2_enexo_3 <= act_regs_data_and_2540_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_12_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2636_enex5 | Relu_for_y_qelse_and_41_enex5 ) begin
      reg_act_regs_data_1_12_2_enexo_3 <= act_regs_data_and_2636_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_91 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_42_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_91 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_91 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_42_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_91 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_91 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_42_enex5 ) begin
      reg_act_config_inst_counter_enexo_91 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_12_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_42_enex5 ) begin
      reg_act_regs_data_0_12_enexo_4 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_12_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2754_enex5 | Relu_for_y_qelse_and_42_enex5 ) begin
      reg_act_regs_data_0_12_3_enexo_3 <= act_regs_data_and_2754_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_12_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2589_enex5 | Relu_for_y_qelse_and_42_enex5 ) begin
      reg_act_regs_data_2_12_3_enexo_3 <= act_regs_data_and_2589_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_12_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2541_enex5 | Relu_for_y_qelse_and_42_enex5 ) begin
      reg_act_regs_data_3_12_3_enexo_3 <= act_regs_data_and_2541_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_12_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2637_enex5 | Relu_for_y_qelse_and_42_enex5 ) begin
      reg_act_regs_data_1_12_3_enexo_3 <= act_regs_data_and_2637_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_92 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_43_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_92 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_11_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_43_enex5 ) begin
      reg_act_regs_data_2_11_enexo_2 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_92 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_43_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_92 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_92 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_43_enex5 ) begin
      reg_act_config_inst_counter_enexo_92 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_11_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2590_enex5 | Relu_for_y_qelse_and_43_enex5 ) begin
      reg_act_regs_data_2_11_1_enexo_3 <= act_regs_data_and_2590_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_11_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2542_enex5 | Relu_for_y_qelse_and_43_enex5 ) begin
      reg_act_regs_data_3_11_1_enexo_3 <= act_regs_data_and_2542_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_11_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2755_enex5 | Relu_for_y_qelse_and_43_enex5 ) begin
      reg_act_regs_data_0_11_1_enexo_3 <= act_regs_data_and_2755_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_11_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2638_enex5 | Relu_for_y_qelse_and_43_enex5 ) begin
      reg_act_regs_data_1_11_1_enexo_3 <= act_regs_data_and_2638_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_93 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_44_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_93 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_11_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_44_enex5 ) begin
      reg_act_regs_data_2_11_enexo_3 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_93 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_44_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_93 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_93 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_44_enex5 ) begin
      reg_act_config_inst_counter_enexo_93 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_11_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2591_enex5 | Relu_for_y_qelse_and_44_enex5 ) begin
      reg_act_regs_data_2_11_2_enexo_3 <= act_regs_data_and_2591_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_11_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2756_enex5 | Relu_for_y_qelse_and_44_enex5 ) begin
      reg_act_regs_data_0_11_2_enexo_3 <= act_regs_data_and_2756_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_11_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2543_enex5 | Relu_for_y_qelse_and_44_enex5 ) begin
      reg_act_regs_data_3_11_2_enexo_3 <= act_regs_data_and_2543_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_11_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2639_enex5 | Relu_for_y_qelse_and_44_enex5 ) begin
      reg_act_regs_data_1_11_2_enexo_3 <= act_regs_data_and_2639_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_94 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_45_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_94 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_11_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_45_enex5 ) begin
      reg_act_regs_data_2_11_enexo_4 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_94 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_45_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_94 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_94 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_45_enex5 ) begin
      reg_act_config_inst_counter_enexo_94 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_11_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2757_enex5 | Relu_for_y_qelse_and_45_enex5 ) begin
      reg_act_regs_data_0_11_3_enexo_3 <= act_regs_data_and_2757_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_11_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2640_enex5 | Relu_for_y_qelse_and_45_enex5 ) begin
      reg_act_regs_data_1_11_3_enexo_3 <= act_regs_data_and_2640_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_11_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2592_enex5 | Relu_for_y_qelse_and_45_enex5 ) begin
      reg_act_regs_data_2_11_3_enexo_3 <= act_regs_data_and_2592_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_11_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2544_enex5 | Relu_for_y_qelse_and_45_enex5 ) begin
      reg_act_regs_data_3_11_3_enexo_3 <= act_regs_data_and_2544_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_95 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_46_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_95 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_95 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_46_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_95 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_95 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_46_enex5 ) begin
      reg_act_config_inst_counter_enexo_95 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_10_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2641_enex5 | Relu_for_y_qelse_and_46_enex5 ) begin
      reg_act_regs_data_1_10_1_enexo_3 <= act_regs_data_and_2641_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_10_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2593_enex5 | Relu_for_y_qelse_and_46_enex5 ) begin
      reg_act_regs_data_2_10_1_enexo_3 <= act_regs_data_and_2593_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_10_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_46_enex5 ) begin
      reg_act_regs_data_0_10_enexo_2 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_10_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2545_enex5 | Relu_for_y_qelse_and_46_enex5 ) begin
      reg_act_regs_data_3_10_1_enexo_3 <= act_regs_data_and_2545_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_10_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2758_enex5 | Relu_for_y_qelse_and_46_enex5 ) begin
      reg_act_regs_data_0_10_1_enexo_3 <= act_regs_data_and_2758_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_96 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_47_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_96 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_96 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_47_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_96 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_96 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_47_enex5 ) begin
      reg_act_config_inst_counter_enexo_96 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_10_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2642_enex5 | Relu_for_y_qelse_and_47_enex5 ) begin
      reg_act_regs_data_1_10_2_enexo_3 <= act_regs_data_and_2642_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_10_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_47_enex5 ) begin
      reg_act_regs_data_0_10_enexo_3 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_10_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2759_enex5 | Relu_for_y_qelse_and_47_enex5 ) begin
      reg_act_regs_data_0_10_2_enexo_3 <= act_regs_data_and_2759_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_10_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2546_enex5 | Relu_for_y_qelse_and_47_enex5 ) begin
      reg_act_regs_data_3_10_2_enexo_3 <= act_regs_data_and_2546_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_10_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2594_enex5 | Relu_for_y_qelse_and_47_enex5 ) begin
      reg_act_regs_data_2_10_2_enexo_3 <= act_regs_data_and_2594_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_97 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_48_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_97 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_97 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_48_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_97 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_97 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_48_enex5 ) begin
      reg_act_config_inst_counter_enexo_97 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_10_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2547_enex5 | Relu_for_y_qelse_and_48_enex5 ) begin
      reg_act_regs_data_3_10_3_enexo_3 <= act_regs_data_and_2547_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_10_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_48_enex5 ) begin
      reg_act_regs_data_0_10_enexo_4 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_10_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2760_enex5 | Relu_for_y_qelse_and_48_enex5 ) begin
      reg_act_regs_data_0_10_3_enexo_3 <= act_regs_data_and_2760_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_10_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2595_enex5 | Relu_for_y_qelse_and_48_enex5 ) begin
      reg_act_regs_data_2_10_3_enexo_3 <= act_regs_data_and_2595_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_10_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2643_enex5 | Relu_for_y_qelse_and_48_enex5 ) begin
      reg_act_regs_data_1_10_3_enexo_3 <= act_regs_data_and_2643_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_98 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_49_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_98 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_98 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_49_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_98 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_98 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_49_enex5 ) begin
      reg_act_config_inst_counter_enexo_98 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_9_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2644_enex5 | Relu_for_y_qelse_and_49_enex5 ) begin
      reg_act_regs_data_1_9_1_enexo_3 <= act_regs_data_and_2644_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_9_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_49_enex5 ) begin
      reg_act_regs_data_1_9_enexo_2 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_9_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2548_enex5 | Relu_for_y_qelse_and_49_enex5 ) begin
      reg_act_regs_data_3_9_1_enexo_3 <= act_regs_data_and_2548_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_9_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2680_enex5 | Relu_for_y_qelse_and_49_enex5 ) begin
      reg_act_regs_data_0_9_1_enexo_3 <= act_regs_data_and_2680_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_9_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2596_enex5 | Relu_for_y_qelse_and_49_enex5 ) begin
      reg_act_regs_data_2_9_1_enexo_3 <= act_regs_data_and_2596_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_99 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_50_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_99 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_99 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_50_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_99 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_99 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_50_enex5 ) begin
      reg_act_config_inst_counter_enexo_99 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_9_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2681_enex5 | Relu_for_y_qelse_and_50_enex5 ) begin
      reg_act_regs_data_0_9_2_enexo_3 <= act_regs_data_and_2681_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_9_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_50_enex5 ) begin
      reg_act_regs_data_1_9_enexo_3 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_9_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2597_enex5 | Relu_for_y_qelse_and_50_enex5 ) begin
      reg_act_regs_data_2_9_2_enexo_3 <= act_regs_data_and_2597_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_9_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2645_enex5 | Relu_for_y_qelse_and_50_enex5 ) begin
      reg_act_regs_data_1_9_2_enexo_3 <= act_regs_data_and_2645_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_9_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2549_enex5 | Relu_for_y_qelse_and_50_enex5 ) begin
      reg_act_regs_data_3_9_2_enexo_3 <= act_regs_data_and_2549_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_100 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_51_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_100 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_100 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_51_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_100 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_100 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_51_enex5 ) begin
      reg_act_config_inst_counter_enexo_100 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_9_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2646_enex5 | Relu_for_y_qelse_and_51_enex5 ) begin
      reg_act_regs_data_1_9_3_enexo_3 <= act_regs_data_and_2646_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_9_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_51_enex5 ) begin
      reg_act_regs_data_1_9_enexo_4 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_9_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2682_enex5 | Relu_for_y_qelse_and_51_enex5 ) begin
      reg_act_regs_data_0_9_3_enexo_3 <= act_regs_data_and_2682_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_9_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2598_enex5 | Relu_for_y_qelse_and_51_enex5 ) begin
      reg_act_regs_data_2_9_3_enexo_3 <= act_regs_data_and_2598_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_9_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2550_enex5 | Relu_for_y_qelse_and_51_enex5 ) begin
      reg_act_regs_data_3_9_3_enexo_3 <= act_regs_data_and_2550_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_101 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_52_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_101 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_101 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_52_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_101 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_101 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_52_enex5 ) begin
      reg_act_config_inst_counter_enexo_101 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_8_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_52_enex5 ) begin
      reg_act_regs_data_2_8_enexo_2 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_8_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2599_enex5 | Relu_for_y_qelse_and_52_enex5 ) begin
      reg_act_regs_data_2_8_1_enexo_3 <= act_regs_data_and_2599_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_8_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2683_enex5 | Relu_for_y_qelse_and_52_enex5 ) begin
      reg_act_regs_data_0_8_1_enexo_3 <= act_regs_data_and_2683_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_8_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2551_enex5 | Relu_for_y_qelse_and_52_enex5 ) begin
      reg_act_regs_data_3_8_1_enexo_3 <= act_regs_data_and_2551_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_8_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2647_enex5 | Relu_for_y_qelse_and_52_enex5 ) begin
      reg_act_regs_data_1_8_1_enexo_3 <= act_regs_data_and_2647_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_102 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_53_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_102 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_102 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_53_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_102 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_102 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_53_enex5 ) begin
      reg_act_config_inst_counter_enexo_102 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_8_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_53_enex5 ) begin
      reg_act_regs_data_2_8_enexo_3 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_8_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2684_enex5 | Relu_for_y_qelse_and_53_enex5 ) begin
      reg_act_regs_data_0_8_2_enexo_3 <= act_regs_data_and_2684_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_8_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2648_enex5 | Relu_for_y_qelse_and_53_enex5 ) begin
      reg_act_regs_data_1_8_2_enexo_3 <= act_regs_data_and_2648_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_8_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2600_enex5 | Relu_for_y_qelse_and_53_enex5 ) begin
      reg_act_regs_data_2_8_2_enexo_3 <= act_regs_data_and_2600_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_8_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2552_enex5 | Relu_for_y_qelse_and_53_enex5 ) begin
      reg_act_regs_data_3_8_2_enexo_3 <= act_regs_data_and_2552_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_103 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_54_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_103 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_103 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_54_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_103 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_103 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_54_enex5 ) begin
      reg_act_config_inst_counter_enexo_103 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_8_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_54_enex5 ) begin
      reg_act_regs_data_2_8_enexo_4 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_8_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2685_enex5 | Relu_for_y_qelse_and_54_enex5 ) begin
      reg_act_regs_data_0_8_3_enexo_3 <= act_regs_data_and_2685_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_8_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2601_enex5 | Relu_for_y_qelse_and_54_enex5 ) begin
      reg_act_regs_data_2_8_3_enexo_3 <= act_regs_data_and_2601_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_8_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2649_enex5 | Relu_for_y_qelse_and_54_enex5 ) begin
      reg_act_regs_data_1_8_3_enexo_3 <= act_regs_data_and_2649_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_8_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2553_enex5 | Relu_for_y_qelse_and_54_enex5 ) begin
      reg_act_regs_data_3_8_3_enexo_3 <= act_regs_data_and_2553_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_104 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_55_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_104 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_104 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_55_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_104 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_104 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_55_enex5 ) begin
      reg_act_config_inst_counter_enexo_104 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_7_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_55_enex5 ) begin
      reg_act_regs_data_1_7_enexo_2 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_7_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2554_enex5 | Relu_for_y_qelse_and_55_enex5 ) begin
      reg_act_regs_data_3_7_1_enexo_3 <= act_regs_data_and_2554_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_7_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2650_enex5 | Relu_for_y_qelse_and_55_enex5 ) begin
      reg_act_regs_data_1_7_1_enexo_3 <= act_regs_data_and_2650_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_7_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2686_enex5 | Relu_for_y_qelse_and_55_enex5 ) begin
      reg_act_regs_data_0_7_1_enexo_3 <= act_regs_data_and_2686_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_7_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2602_enex5 | Relu_for_y_qelse_and_55_enex5 ) begin
      reg_act_regs_data_2_7_1_enexo_3 <= act_regs_data_and_2602_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_105 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_56_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_105 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_105 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_56_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_105 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_105 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_56_enex5 ) begin
      reg_act_config_inst_counter_enexo_105 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_7_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_56_enex5 ) begin
      reg_act_regs_data_1_7_enexo_3 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_7_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2687_enex5 | Relu_for_y_qelse_and_56_enex5 ) begin
      reg_act_regs_data_0_7_2_enexo_3 <= act_regs_data_and_2687_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_7_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2603_enex5 | Relu_for_y_qelse_and_56_enex5 ) begin
      reg_act_regs_data_2_7_2_enexo_3 <= act_regs_data_and_2603_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_7_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2555_enex5 | Relu_for_y_qelse_and_56_enex5 ) begin
      reg_act_regs_data_3_7_2_enexo_3 <= act_regs_data_and_2555_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_7_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2651_enex5 | Relu_for_y_qelse_and_56_enex5 ) begin
      reg_act_regs_data_1_7_2_enexo_3 <= act_regs_data_and_2651_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_106 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_57_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_106 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_106 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_57_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_106 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_106 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_57_enex5 ) begin
      reg_act_config_inst_counter_enexo_106 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_7_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2688_enex5 | Relu_for_y_qelse_and_57_enex5 ) begin
      reg_act_regs_data_0_7_3_enexo_3 <= act_regs_data_and_2688_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_7_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2652_enex5 | Relu_for_y_qelse_and_57_enex5 ) begin
      reg_act_regs_data_1_7_3_enexo_3 <= act_regs_data_and_2652_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_7_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2556_enex5 | Relu_for_y_qelse_and_57_enex5 ) begin
      reg_act_regs_data_3_7_3_enexo_3 <= act_regs_data_and_2556_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_7_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_57_enex5 ) begin
      reg_act_regs_data_1_7_enexo_4 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_7_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2604_enex5 | Relu_for_y_qelse_and_57_enex5 ) begin
      reg_act_regs_data_2_7_3_enexo_3 <= act_regs_data_and_2604_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_107 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_58_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_107 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_107 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_58_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_107 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_107 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_58_enex5 ) begin
      reg_act_config_inst_counter_enexo_107 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_6_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2557_enex5 | Relu_for_y_qelse_and_58_enex5 ) begin
      reg_act_regs_data_3_6_1_enexo_3 <= act_regs_data_and_2557_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_6_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2653_enex5 | Relu_for_y_qelse_and_58_enex5 ) begin
      reg_act_regs_data_1_6_1_enexo_3 <= act_regs_data_and_2653_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_6_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_58_enex5 ) begin
      reg_act_regs_data_3_6_enexo_2 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_6_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2605_enex5 | Relu_for_y_qelse_and_58_enex5 ) begin
      reg_act_regs_data_2_6_1_enexo_3 <= act_regs_data_and_2605_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_6_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2689_enex5 | Relu_for_y_qelse_and_58_enex5 ) begin
      reg_act_regs_data_0_6_1_enexo_3 <= act_regs_data_and_2689_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_108 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_59_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_108 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_108 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_59_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_108 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_108 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_59_enex5 ) begin
      reg_act_config_inst_counter_enexo_108 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_6_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_59_enex5 ) begin
      reg_act_regs_data_3_6_enexo_3 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_6_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2606_enex5 | Relu_for_y_qelse_and_59_enex5 ) begin
      reg_act_regs_data_2_6_2_enexo_3 <= act_regs_data_and_2606_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_6_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2654_enex5 | Relu_for_y_qelse_and_59_enex5 ) begin
      reg_act_regs_data_1_6_2_enexo_3 <= act_regs_data_and_2654_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_6_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2558_enex5 | Relu_for_y_qelse_and_59_enex5 ) begin
      reg_act_regs_data_3_6_2_enexo_3 <= act_regs_data_and_2558_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_6_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2690_enex5 | Relu_for_y_qelse_and_59_enex5 ) begin
      reg_act_regs_data_0_6_2_enexo_3 <= act_regs_data_and_2690_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_109 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_60_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_109 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_109 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_60_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_109 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_109 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_60_enex5 ) begin
      reg_act_config_inst_counter_enexo_109 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_6_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2607_enex5 | Relu_for_y_qelse_and_60_enex5 ) begin
      reg_act_regs_data_2_6_3_enexo_3 <= act_regs_data_and_2607_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_6_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2559_enex5 | Relu_for_y_qelse_and_60_enex5 ) begin
      reg_act_regs_data_3_6_3_enexo_3 <= act_regs_data_and_2559_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_6_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_60_enex5 ) begin
      reg_act_regs_data_3_6_enexo_4 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_6_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2691_enex5 | Relu_for_y_qelse_and_60_enex5 ) begin
      reg_act_regs_data_0_6_3_enexo_3 <= act_regs_data_and_2691_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_6_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2655_enex5 | Relu_for_y_qelse_and_60_enex5 ) begin
      reg_act_regs_data_1_6_3_enexo_3 <= act_regs_data_and_2655_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_110 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_61_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_110 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_110 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_61_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_110 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_110 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_61_enex5 ) begin
      reg_act_config_inst_counter_enexo_110 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_5_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2560_enex5 | Relu_for_y_qelse_and_61_enex5 ) begin
      reg_act_regs_data_3_5_1_enexo_3 <= act_regs_data_and_2560_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_5_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2692_enex5 | Relu_for_y_qelse_and_61_enex5 ) begin
      reg_act_regs_data_0_5_1_enexo_3 <= act_regs_data_and_2692_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_5_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_61_enex5 ) begin
      reg_act_regs_data_1_5_enexo_2 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_5_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2656_enex5 | Relu_for_y_qelse_and_61_enex5 ) begin
      reg_act_regs_data_1_5_1_enexo_3 <= act_regs_data_and_2656_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_5_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2608_enex5 | Relu_for_y_qelse_and_61_enex5 ) begin
      reg_act_regs_data_2_5_1_enexo_3 <= act_regs_data_and_2608_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_111 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_62_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_111 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_111 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_62_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_111 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_111 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_62_enex5 ) begin
      reg_act_config_inst_counter_enexo_111 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_5_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2609_enex5 | Relu_for_y_qelse_and_62_enex5 ) begin
      reg_act_regs_data_2_5_2_enexo_3 <= act_regs_data_and_2609_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_5_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_62_enex5 ) begin
      reg_act_regs_data_1_5_enexo_3 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_5_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2657_enex5 | Relu_for_y_qelse_and_62_enex5 ) begin
      reg_act_regs_data_1_5_2_enexo_3 <= act_regs_data_and_2657_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_5_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2561_enex5 | Relu_for_y_qelse_and_62_enex5 ) begin
      reg_act_regs_data_3_5_2_enexo_3 <= act_regs_data_and_2561_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_5_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2693_enex5 | Relu_for_y_qelse_and_62_enex5 ) begin
      reg_act_regs_data_0_5_2_enexo_3 <= act_regs_data_and_2693_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_112 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_63_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_112 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_112 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_63_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_112 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_5_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2694_enex5 | Relu_for_y_qelse_and_63_enex5 ) begin
      reg_act_regs_data_0_5_3_enexo_3 <= act_regs_data_and_2694_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_112 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_63_enex5 ) begin
      reg_act_config_inst_counter_enexo_112 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_5_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_63_enex5 ) begin
      reg_act_regs_data_1_5_enexo_4 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_5_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2658_enex5 | Relu_for_y_qelse_and_63_enex5 ) begin
      reg_act_regs_data_1_5_3_enexo_3 <= act_regs_data_and_2658_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_5_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2562_enex5 | Relu_for_y_qelse_and_63_enex5 ) begin
      reg_act_regs_data_3_5_3_enexo_3 <= act_regs_data_and_2562_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_5_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2610_enex5 | Relu_for_y_qelse_and_63_enex5 ) begin
      reg_act_regs_data_2_5_3_enexo_3 <= act_regs_data_and_2610_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_113 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_64_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_113 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_113 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_64_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_113 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_113 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_64_enex5 ) begin
      reg_act_config_inst_counter_enexo_113 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_4_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2563_enex5 | Relu_for_y_qelse_and_64_enex5 ) begin
      reg_act_regs_data_3_4_1_enexo_3 <= act_regs_data_and_2563_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_4_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2695_enex5 | Relu_for_y_qelse_and_64_enex5 ) begin
      reg_act_regs_data_0_4_1_enexo_3 <= act_regs_data_and_2695_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_4_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2611_enex5 | Relu_for_y_qelse_and_64_enex5 ) begin
      reg_act_regs_data_2_4_1_enexo_3 <= act_regs_data_and_2611_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_4_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_64_enex5 ) begin
      reg_act_regs_data_3_4_enexo_2 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_4_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2659_enex5 | Relu_for_y_qelse_and_64_enex5 ) begin
      reg_act_regs_data_1_4_1_enexo_3 <= act_regs_data_and_2659_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_114 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_65_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_114 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_114 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_65_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_114 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_114 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_65_enex5 ) begin
      reg_act_config_inst_counter_enexo_114 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_4_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2564_enex5 | Relu_for_y_qelse_and_65_enex5 ) begin
      reg_act_regs_data_3_4_2_enexo_3 <= act_regs_data_and_2564_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_4_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2660_enex5 | Relu_for_y_qelse_and_65_enex5 ) begin
      reg_act_regs_data_1_4_2_enexo_3 <= act_regs_data_and_2660_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_4_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_65_enex5 ) begin
      reg_act_regs_data_3_4_enexo_3 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_4_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2696_enex5 | Relu_for_y_qelse_and_65_enex5 ) begin
      reg_act_regs_data_0_4_2_enexo_3 <= act_regs_data_and_2696_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_4_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2612_enex5 | Relu_for_y_qelse_and_65_enex5 ) begin
      reg_act_regs_data_2_4_2_enexo_3 <= act_regs_data_and_2612_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_115 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_66_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_115 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_115 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_66_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_115 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_115 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_66_enex5 ) begin
      reg_act_config_inst_counter_enexo_115 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_4_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2697_enex5 | Relu_for_y_qelse_and_66_enex5 ) begin
      reg_act_regs_data_0_4_3_enexo_3 <= act_regs_data_and_2697_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_4_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2661_enex5 | Relu_for_y_qelse_and_66_enex5 ) begin
      reg_act_regs_data_1_4_3_enexo_3 <= act_regs_data_and_2661_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_4_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2565_enex5 | Relu_for_y_qelse_and_66_enex5 ) begin
      reg_act_regs_data_3_4_3_enexo_3 <= act_regs_data_and_2565_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_4_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_66_enex5 ) begin
      reg_act_regs_data_3_4_enexo_4 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_4_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2613_enex5 | Relu_for_y_qelse_and_66_enex5 ) begin
      reg_act_regs_data_2_4_3_enexo_3 <= act_regs_data_and_2613_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_116 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_67_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_116 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_116 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_67_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_116 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_116 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_67_enex5 ) begin
      reg_act_config_inst_counter_enexo_116 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_3_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2698_enex5 | Relu_for_y_qelse_and_67_enex5 ) begin
      reg_act_regs_data_0_3_1_enexo_3 <= act_regs_data_and_2698_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_3_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_67_enex5 ) begin
      reg_act_regs_data_3_3_enexo_2 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_3_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2566_enex5 | Relu_for_y_qelse_and_67_enex5 ) begin
      reg_act_regs_data_3_3_1_enexo_3 <= act_regs_data_and_2566_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_3_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2662_enex5 | Relu_for_y_qelse_and_67_enex5 ) begin
      reg_act_regs_data_1_3_1_enexo_3 <= act_regs_data_and_2662_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_3_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2614_enex5 | Relu_for_y_qelse_and_67_enex5 ) begin
      reg_act_regs_data_2_3_1_enexo_3 <= act_regs_data_and_2614_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_117 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_68_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_117 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_117 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_68_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_117 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_117 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_68_enex5 ) begin
      reg_act_config_inst_counter_enexo_117 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_68_enex5 ) begin
      reg_act_regs_data_3_3_enexo_3 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_3_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2699_enex5 | Relu_for_y_qelse_and_68_enex5 ) begin
      reg_act_regs_data_0_3_2_enexo_3 <= act_regs_data_and_2699_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_3_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2663_enex5 | Relu_for_y_qelse_and_68_enex5 ) begin
      reg_act_regs_data_1_3_2_enexo_3 <= act_regs_data_and_2663_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_3_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2567_enex5 | Relu_for_y_qelse_and_68_enex5 ) begin
      reg_act_regs_data_3_3_2_enexo_3 <= act_regs_data_and_2567_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_3_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2615_enex5 | Relu_for_y_qelse_and_68_enex5 ) begin
      reg_act_regs_data_2_3_2_enexo_3 <= act_regs_data_and_2615_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_118 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_69_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_118 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_118 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_69_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_118 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_118 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_69_enex5 ) begin
      reg_act_config_inst_counter_enexo_118 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_3_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2700_enex5 | Relu_for_y_qelse_and_69_enex5 ) begin
      reg_act_regs_data_0_3_3_enexo_3 <= act_regs_data_and_2700_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_3_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2568_enex5 | Relu_for_y_qelse_and_69_enex5 ) begin
      reg_act_regs_data_3_3_3_enexo_3 <= act_regs_data_and_2568_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_69_enex5 ) begin
      reg_act_regs_data_3_3_enexo_4 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_3_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2664_enex5 | Relu_for_y_qelse_and_69_enex5 ) begin
      reg_act_regs_data_1_3_3_enexo_3 <= act_regs_data_and_2664_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_3_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2616_enex5 | Relu_for_y_qelse_and_69_enex5 ) begin
      reg_act_regs_data_2_3_3_enexo_3 <= act_regs_data_and_2616_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_2_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2617_enex5 | Relu_for_y_qelse_and_70_enex5 ) begin
      reg_act_regs_data_2_2_1_enexo_3 <= act_regs_data_and_2617_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_119 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_70_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_119 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_119 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_70_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_119 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_119 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_70_enex5 ) begin
      reg_act_config_inst_counter_enexo_119 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_2_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_70_enex5 ) begin
      reg_act_regs_data_3_2_enexo_2 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_2_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2569_enex5 | Relu_for_y_qelse_and_70_enex5 ) begin
      reg_act_regs_data_3_2_1_enexo_3 <= act_regs_data_and_2569_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_2_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2665_enex5 | Relu_for_y_qelse_and_70_enex5 ) begin
      reg_act_regs_data_1_2_1_enexo_3 <= act_regs_data_and_2665_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_2_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2701_enex5 | Relu_for_y_qelse_and_70_enex5 ) begin
      reg_act_regs_data_0_2_1_enexo_3 <= act_regs_data_and_2701_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_120 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_71_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_120 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_120 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_71_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_120 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_120 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_71_enex5 ) begin
      reg_act_config_inst_counter_enexo_120 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_71_enex5 ) begin
      reg_act_regs_data_3_2_enexo_3 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_2_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2702_enex5 | Relu_for_y_qelse_and_71_enex5 ) begin
      reg_act_regs_data_0_2_2_enexo_3 <= act_regs_data_and_2702_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_2_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2666_enex5 | Relu_for_y_qelse_and_71_enex5 ) begin
      reg_act_regs_data_1_2_2_enexo_3 <= act_regs_data_and_2666_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_2_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2570_enex5 | Relu_for_y_qelse_and_71_enex5 ) begin
      reg_act_regs_data_3_2_2_enexo_3 <= act_regs_data_and_2570_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_2_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2618_enex5 | Relu_for_y_qelse_and_71_enex5 ) begin
      reg_act_regs_data_2_2_2_enexo_3 <= act_regs_data_and_2618_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_121 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_72_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_121 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_121 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_72_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_121 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_121 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_72_enex5 ) begin
      reg_act_config_inst_counter_enexo_121 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_72_enex5 ) begin
      reg_act_regs_data_3_2_enexo_4 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_2_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2571_enex5 | Relu_for_y_qelse_and_72_enex5 ) begin
      reg_act_regs_data_3_2_3_enexo_3 <= act_regs_data_and_2571_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_2_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2619_enex5 | Relu_for_y_qelse_and_72_enex5 ) begin
      reg_act_regs_data_2_2_3_enexo_3 <= act_regs_data_and_2619_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_2_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2703_enex5 | Relu_for_y_qelse_and_72_enex5 ) begin
      reg_act_regs_data_0_2_3_enexo_3 <= act_regs_data_and_2703_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_2_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2667_enex5 | Relu_for_y_qelse_and_72_enex5 ) begin
      reg_act_regs_data_1_2_3_enexo_3 <= act_regs_data_and_2667_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_122 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_73_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_122 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_122 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_73_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_122 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_1_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2620_enex5 | Relu_for_y_qelse_and_73_enex5 ) begin
      reg_act_regs_data_2_1_1_enexo_3 <= act_regs_data_and_2620_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_122 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_73_enex5 ) begin
      reg_act_config_inst_counter_enexo_122 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_1_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2572_enex5 | Relu_for_y_qelse_and_73_enex5 ) begin
      reg_act_regs_data_3_1_1_enexo_3 <= act_regs_data_and_2572_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_1_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_73_enex5 ) begin
      reg_act_regs_data_2_1_enexo_2 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_1_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2761_enex5 | Relu_for_y_qelse_and_73_enex5 ) begin
      reg_act_regs_data_0_1_1_enexo_3 <= act_regs_data_and_2761_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_1_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2668_enex5 | Relu_for_y_qelse_and_73_enex5 ) begin
      reg_act_regs_data_1_1_1_enexo_3 <= act_regs_data_and_2668_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_123 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_74_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_123 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_123 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_74_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_123 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_123 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_74_enex5 ) begin
      reg_act_config_inst_counter_enexo_123 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_1_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2669_enex5 | Relu_for_y_qelse_and_74_enex5 ) begin
      reg_act_regs_data_1_1_2_enexo_3 <= act_regs_data_and_2669_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_74_enex5 ) begin
      reg_act_regs_data_2_1_enexo_3 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_1_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2573_enex5 | Relu_for_y_qelse_and_74_enex5 ) begin
      reg_act_regs_data_3_1_2_enexo_3 <= act_regs_data_and_2573_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_1_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2762_enex5 | Relu_for_y_qelse_and_74_enex5 ) begin
      reg_act_regs_data_0_1_2_enexo_3 <= act_regs_data_and_2762_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_1_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2621_enex5 | Relu_for_y_qelse_and_74_enex5 ) begin
      reg_act_regs_data_2_1_2_enexo_3 <= act_regs_data_and_2621_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_124 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_75_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_124 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_124 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_75_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_124 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_124 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_75_enex5 ) begin
      reg_act_config_inst_counter_enexo_124 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_1_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2763_enex5 | Relu_for_y_qelse_and_75_enex5 ) begin
      reg_act_regs_data_0_1_3_enexo_3 <= act_regs_data_and_2763_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_75_enex5 ) begin
      reg_act_regs_data_2_1_enexo_4 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_1_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2574_enex5 | Relu_for_y_qelse_and_75_enex5 ) begin
      reg_act_regs_data_3_1_3_enexo_3 <= act_regs_data_and_2574_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_1_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2670_enex5 | Relu_for_y_qelse_and_75_enex5 ) begin
      reg_act_regs_data_1_1_3_enexo_3 <= act_regs_data_and_2670_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_1_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2622_enex5 | Relu_for_y_qelse_and_75_enex5 ) begin
      reg_act_regs_data_2_1_3_enexo_3 <= act_regs_data_and_2622_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_125 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_76_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_125 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_0_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2575_enex5 | Relu_for_y_qelse_and_76_enex5 ) begin
      reg_act_regs_data_3_0_1_enexo_3 <= act_regs_data_and_2575_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_0_enexo_2 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_76_enex5 ) begin
      reg_act_regs_data_3_0_enexo_2 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_125 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_76_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_125 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_125 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_76_enex5 ) begin
      reg_act_config_inst_counter_enexo_125 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_0_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2764_enex5 | Relu_for_y_qelse_and_76_enex5 ) begin
      reg_act_regs_data_0_0_1_enexo_3 <= act_regs_data_and_2764_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_0_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2623_enex5 | Relu_for_y_qelse_and_76_enex5 ) begin
      reg_act_regs_data_2_0_1_enexo_3 <= act_regs_data_and_2623_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_0_1_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2671_enex5 | Relu_for_y_qelse_and_76_enex5 ) begin
      reg_act_regs_data_1_0_1_enexo_3 <= act_regs_data_and_2671_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_126 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_77_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_126 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_0_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_77_enex5 ) begin
      reg_act_regs_data_3_0_enexo_3 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_126 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_77_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_126 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_126 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_77_enex5 ) begin
      reg_act_config_inst_counter_enexo_126 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_0_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2576_enex5 | Relu_for_y_qelse_and_77_enex5 ) begin
      reg_act_regs_data_3_0_2_enexo_3 <= act_regs_data_and_2576_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_0_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2765_enex5 | Relu_for_y_qelse_and_77_enex5 ) begin
      reg_act_regs_data_0_0_2_enexo_3 <= act_regs_data_and_2765_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_0_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2672_enex5 | Relu_for_y_qelse_and_77_enex5 ) begin
      reg_act_regs_data_1_0_2_enexo_3 <= act_regs_data_and_2672_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_0_2_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2624_enex5 | Relu_for_y_qelse_and_77_enex5 ) begin
      reg_act_regs_data_2_0_2_enexo_3 <= act_regs_data_and_2624_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_127 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | Relu_for_y_qelse_and_78_enex5 ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_127 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_0_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_ssc | Relu_for_y_qelse_and_78_enex5 ) begin
      reg_act_regs_data_3_0_enexo_4 <= act_regs_data_and_ssc;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_127 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | Relu_for_y_qelse_and_78_enex5 ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_127 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_127 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | Relu_for_y_qelse_and_78_enex5 ) begin
      reg_act_config_inst_counter_enexo_127 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_0_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2577_enex5 | Relu_for_y_qelse_and_78_enex5 ) begin
      reg_act_regs_data_3_0_3_enexo_3 <= act_regs_data_and_2577_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_0_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2766_enex5 | Relu_for_y_qelse_and_78_enex5 ) begin
      reg_act_regs_data_0_0_3_enexo_3 <= act_regs_data_and_2766_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_0_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2625_enex5 | Relu_for_y_qelse_and_78_enex5 ) begin
      reg_act_regs_data_2_0_3_enexo_3 <= act_regs_data_and_2625_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_0_3_enexo_3 <= 1'b1;
    end
    else if ( act_regs_data_and_2673_enex5 | Relu_for_y_qelse_and_78_enex5 ) begin
      reg_act_regs_data_1_0_3_enexo_3 <= act_regs_data_and_2673_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_128 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | ActUnit_RunInst_curr_inst_and_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_128 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_128 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | ActUnit_RunInst_curr_inst_and_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_128 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_128 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | ActUnit_RunInst_curr_inst_and_enex5
        ) begin
      reg_act_config_inst_counter_enexo_128 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_129 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | ActUnit_RunInst_switch_lp_and_813_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_129 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_129 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | ActUnit_RunInst_switch_lp_and_813_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_129 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_129 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | ActUnit_RunInst_switch_lp_and_813_enex5
        ) begin
      reg_act_config_inst_counter_enexo_129 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_0_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2576_enex5 | ActUnit_RunInst_switch_lp_and_813_enex5
        ) begin
      reg_act_regs_data_3_0_2_enexo_4 <= act_regs_data_and_2576_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_0_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2765_enex5 | ActUnit_RunInst_switch_lp_and_813_enex5
        ) begin
      reg_act_regs_data_0_0_2_enexo_4 <= act_regs_data_and_2765_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_0_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2672_enex5 | ActUnit_RunInst_switch_lp_and_813_enex5
        ) begin
      reg_act_regs_data_1_0_2_enexo_4 <= act_regs_data_and_2672_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_0_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2624_enex5 | ActUnit_RunInst_switch_lp_and_813_enex5
        ) begin
      reg_act_regs_data_2_0_2_enexo_4 <= act_regs_data_and_2624_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_130 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | ActUnit_RunInst_switch_lp_and_814_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_130 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_130 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | ActUnit_RunInst_switch_lp_and_814_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_130 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_130 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | ActUnit_RunInst_switch_lp_and_814_enex5
        ) begin
      reg_act_config_inst_counter_enexo_130 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_0_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2577_enex5 | ActUnit_RunInst_switch_lp_and_814_enex5
        ) begin
      reg_act_regs_data_3_0_3_enexo_4 <= act_regs_data_and_2577_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_0_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2766_enex5 | ActUnit_RunInst_switch_lp_and_814_enex5
        ) begin
      reg_act_regs_data_0_0_3_enexo_4 <= act_regs_data_and_2766_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_0_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2625_enex5 | ActUnit_RunInst_switch_lp_and_814_enex5
        ) begin
      reg_act_regs_data_2_0_3_enexo_4 <= act_regs_data_and_2625_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_0_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2673_enex5 | ActUnit_RunInst_switch_lp_and_814_enex5
        ) begin
      reg_act_regs_data_1_0_3_enexo_4 <= act_regs_data_and_2673_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_131 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | ActUnit_RunInst_switch_lp_and_815_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_131 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_0_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2575_enex5 | ActUnit_RunInst_switch_lp_and_815_enex5
        ) begin
      reg_act_regs_data_3_0_1_enexo_4 <= act_regs_data_and_2575_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_131 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | ActUnit_RunInst_switch_lp_and_815_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_131 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_131 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | ActUnit_RunInst_switch_lp_and_815_enex5
        ) begin
      reg_act_config_inst_counter_enexo_131 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_0_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2764_enex5 | ActUnit_RunInst_switch_lp_and_815_enex5
        ) begin
      reg_act_regs_data_0_0_1_enexo_4 <= act_regs_data_and_2764_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_0_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2623_enex5 | ActUnit_RunInst_switch_lp_and_815_enex5
        ) begin
      reg_act_regs_data_2_0_1_enexo_4 <= act_regs_data_and_2623_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_0_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2671_enex5 | ActUnit_RunInst_switch_lp_and_815_enex5
        ) begin
      reg_act_regs_data_1_0_1_enexo_4 <= act_regs_data_and_2671_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_132 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_132 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_132 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_132 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_132 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_enex5
        ) begin
      reg_act_config_inst_counter_enexo_132 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_1_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2669_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_enex5
        ) begin
      reg_act_regs_data_1_1_2_enexo_4 <= act_regs_data_and_2669_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_1_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2573_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_enex5
        ) begin
      reg_act_regs_data_3_1_2_enexo_4 <= act_regs_data_and_2573_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_1_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2762_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_enex5
        ) begin
      reg_act_regs_data_0_1_2_enexo_4 <= act_regs_data_and_2762_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_1_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2621_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_enex5
        ) begin
      reg_act_regs_data_2_1_2_enexo_4 <= act_regs_data_and_2621_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_133 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_15_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_133 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_133 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_15_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_133 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_133 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_15_enex5
        ) begin
      reg_act_config_inst_counter_enexo_133 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_1_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2763_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_15_enex5
        ) begin
      reg_act_regs_data_0_1_3_enexo_4 <= act_regs_data_and_2763_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_1_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2574_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_15_enex5
        ) begin
      reg_act_regs_data_3_1_3_enexo_4 <= act_regs_data_and_2574_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_1_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2670_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_15_enex5
        ) begin
      reg_act_regs_data_1_1_3_enexo_4 <= act_regs_data_and_2670_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_1_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2622_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_15_enex5
        ) begin
      reg_act_regs_data_2_1_3_enexo_4 <= act_regs_data_and_2622_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_134 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_16_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_134 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_134 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_16_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_134 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_1_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2620_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_16_enex5
        ) begin
      reg_act_regs_data_2_1_1_enexo_4 <= act_regs_data_and_2620_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_134 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_16_enex5
        ) begin
      reg_act_config_inst_counter_enexo_134 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_1_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2572_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_16_enex5
        ) begin
      reg_act_regs_data_3_1_1_enexo_4 <= act_regs_data_and_2572_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_1_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2761_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_16_enex5
        ) begin
      reg_act_regs_data_0_1_1_enexo_4 <= act_regs_data_and_2761_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_1_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2668_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_16_enex5
        ) begin
      reg_act_regs_data_1_1_1_enexo_4 <= act_regs_data_and_2668_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_135 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_17_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_135 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_135 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_17_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_135 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_135 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_17_enex5
        ) begin
      reg_act_config_inst_counter_enexo_135 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_2_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2702_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_17_enex5
        ) begin
      reg_act_regs_data_0_2_2_enexo_4 <= act_regs_data_and_2702_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_2_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2666_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_17_enex5
        ) begin
      reg_act_regs_data_1_2_2_enexo_4 <= act_regs_data_and_2666_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_2_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2570_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_17_enex5
        ) begin
      reg_act_regs_data_3_2_2_enexo_4 <= act_regs_data_and_2570_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_2_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2618_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_17_enex5
        ) begin
      reg_act_regs_data_2_2_2_enexo_4 <= act_regs_data_and_2618_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_136 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_18_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_136 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_136 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_18_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_136 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_136 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_18_enex5
        ) begin
      reg_act_config_inst_counter_enexo_136 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_2_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2571_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_18_enex5
        ) begin
      reg_act_regs_data_3_2_3_enexo_4 <= act_regs_data_and_2571_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_2_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2619_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_18_enex5
        ) begin
      reg_act_regs_data_2_2_3_enexo_4 <= act_regs_data_and_2619_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_2_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2703_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_18_enex5
        ) begin
      reg_act_regs_data_0_2_3_enexo_4 <= act_regs_data_and_2703_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_2_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2667_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_18_enex5
        ) begin
      reg_act_regs_data_1_2_3_enexo_4 <= act_regs_data_and_2667_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_2_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2617_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_19_enex5
        ) begin
      reg_act_regs_data_2_2_1_enexo_4 <= act_regs_data_and_2617_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_137 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_19_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_137 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_137 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_19_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_137 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_137 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_19_enex5
        ) begin
      reg_act_config_inst_counter_enexo_137 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_2_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2569_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_19_enex5
        ) begin
      reg_act_regs_data_3_2_1_enexo_4 <= act_regs_data_and_2569_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_2_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2665_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_19_enex5
        ) begin
      reg_act_regs_data_1_2_1_enexo_4 <= act_regs_data_and_2665_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_2_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2701_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_19_enex5
        ) begin
      reg_act_regs_data_0_2_1_enexo_4 <= act_regs_data_and_2701_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_138 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_20_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_138 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_138 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_20_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_138 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_138 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_20_enex5
        ) begin
      reg_act_config_inst_counter_enexo_138 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_3_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2699_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_20_enex5
        ) begin
      reg_act_regs_data_0_3_2_enexo_4 <= act_regs_data_and_2699_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_3_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2663_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_20_enex5
        ) begin
      reg_act_regs_data_1_3_2_enexo_4 <= act_regs_data_and_2663_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_3_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2567_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_20_enex5
        ) begin
      reg_act_regs_data_3_3_2_enexo_4 <= act_regs_data_and_2567_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_3_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2615_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_20_enex5
        ) begin
      reg_act_regs_data_2_3_2_enexo_4 <= act_regs_data_and_2615_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_139 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_21_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_139 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_139 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_21_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_139 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_139 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_21_enex5
        ) begin
      reg_act_config_inst_counter_enexo_139 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_3_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2700_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_21_enex5
        ) begin
      reg_act_regs_data_0_3_3_enexo_4 <= act_regs_data_and_2700_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_3_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2568_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_21_enex5
        ) begin
      reg_act_regs_data_3_3_3_enexo_4 <= act_regs_data_and_2568_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_3_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2664_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_21_enex5
        ) begin
      reg_act_regs_data_1_3_3_enexo_4 <= act_regs_data_and_2664_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_3_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2616_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_21_enex5
        ) begin
      reg_act_regs_data_2_3_3_enexo_4 <= act_regs_data_and_2616_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_140 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_22_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_140 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_140 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_22_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_140 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_140 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_22_enex5
        ) begin
      reg_act_config_inst_counter_enexo_140 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_3_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2698_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_22_enex5
        ) begin
      reg_act_regs_data_0_3_1_enexo_4 <= act_regs_data_and_2698_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_3_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2566_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_22_enex5
        ) begin
      reg_act_regs_data_3_3_1_enexo_4 <= act_regs_data_and_2566_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_3_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2662_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_22_enex5
        ) begin
      reg_act_regs_data_1_3_1_enexo_4 <= act_regs_data_and_2662_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_3_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2614_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_22_enex5
        ) begin
      reg_act_regs_data_2_3_1_enexo_4 <= act_regs_data_and_2614_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_141 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_23_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_141 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_141 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_23_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_141 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_141 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_23_enex5
        ) begin
      reg_act_config_inst_counter_enexo_141 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_4_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2564_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_23_enex5
        ) begin
      reg_act_regs_data_3_4_2_enexo_4 <= act_regs_data_and_2564_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_4_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2660_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_23_enex5
        ) begin
      reg_act_regs_data_1_4_2_enexo_4 <= act_regs_data_and_2660_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_4_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2696_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_23_enex5
        ) begin
      reg_act_regs_data_0_4_2_enexo_4 <= act_regs_data_and_2696_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_4_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2612_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_23_enex5
        ) begin
      reg_act_regs_data_2_4_2_enexo_4 <= act_regs_data_and_2612_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_142 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_24_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_142 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_142 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_24_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_142 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_142 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_24_enex5
        ) begin
      reg_act_config_inst_counter_enexo_142 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_4_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2697_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_24_enex5
        ) begin
      reg_act_regs_data_0_4_3_enexo_4 <= act_regs_data_and_2697_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_4_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2661_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_24_enex5
        ) begin
      reg_act_regs_data_1_4_3_enexo_4 <= act_regs_data_and_2661_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_4_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2565_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_24_enex5
        ) begin
      reg_act_regs_data_3_4_3_enexo_4 <= act_regs_data_and_2565_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_4_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2613_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_24_enex5
        ) begin
      reg_act_regs_data_2_4_3_enexo_4 <= act_regs_data_and_2613_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_143 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_25_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_143 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_143 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_25_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_143 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_143 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_25_enex5
        ) begin
      reg_act_config_inst_counter_enexo_143 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_4_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2563_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_25_enex5
        ) begin
      reg_act_regs_data_3_4_1_enexo_4 <= act_regs_data_and_2563_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_4_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2695_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_25_enex5
        ) begin
      reg_act_regs_data_0_4_1_enexo_4 <= act_regs_data_and_2695_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_4_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2611_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_25_enex5
        ) begin
      reg_act_regs_data_2_4_1_enexo_4 <= act_regs_data_and_2611_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_4_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2659_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_25_enex5
        ) begin
      reg_act_regs_data_1_4_1_enexo_4 <= act_regs_data_and_2659_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_144 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_26_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_144 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_144 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_26_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_144 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_144 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_26_enex5
        ) begin
      reg_act_config_inst_counter_enexo_144 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_5_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2609_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_26_enex5
        ) begin
      reg_act_regs_data_2_5_2_enexo_4 <= act_regs_data_and_2609_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_5_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2657_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_26_enex5
        ) begin
      reg_act_regs_data_1_5_2_enexo_4 <= act_regs_data_and_2657_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_5_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2561_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_26_enex5
        ) begin
      reg_act_regs_data_3_5_2_enexo_4 <= act_regs_data_and_2561_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_5_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2693_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_26_enex5
        ) begin
      reg_act_regs_data_0_5_2_enexo_4 <= act_regs_data_and_2693_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_145 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_27_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_145 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_145 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_27_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_145 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_5_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2694_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_27_enex5
        ) begin
      reg_act_regs_data_0_5_3_enexo_4 <= act_regs_data_and_2694_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_145 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_27_enex5
        ) begin
      reg_act_config_inst_counter_enexo_145 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_5_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2658_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_27_enex5
        ) begin
      reg_act_regs_data_1_5_3_enexo_4 <= act_regs_data_and_2658_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_5_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2562_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_27_enex5
        ) begin
      reg_act_regs_data_3_5_3_enexo_4 <= act_regs_data_and_2562_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_5_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2610_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_27_enex5
        ) begin
      reg_act_regs_data_2_5_3_enexo_4 <= act_regs_data_and_2610_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_146 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_28_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_146 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_146 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_28_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_146 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_146 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_28_enex5
        ) begin
      reg_act_config_inst_counter_enexo_146 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_5_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2560_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_28_enex5
        ) begin
      reg_act_regs_data_3_5_1_enexo_4 <= act_regs_data_and_2560_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_5_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2692_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_28_enex5
        ) begin
      reg_act_regs_data_0_5_1_enexo_4 <= act_regs_data_and_2692_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_5_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2656_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_28_enex5
        ) begin
      reg_act_regs_data_1_5_1_enexo_4 <= act_regs_data_and_2656_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_5_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2608_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_28_enex5
        ) begin
      reg_act_regs_data_2_5_1_enexo_4 <= act_regs_data_and_2608_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_147 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_29_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_147 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_147 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_29_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_147 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_147 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_29_enex5
        ) begin
      reg_act_config_inst_counter_enexo_147 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_6_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2606_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_29_enex5
        ) begin
      reg_act_regs_data_2_6_2_enexo_4 <= act_regs_data_and_2606_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_6_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2654_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_29_enex5
        ) begin
      reg_act_regs_data_1_6_2_enexo_4 <= act_regs_data_and_2654_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_6_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2558_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_29_enex5
        ) begin
      reg_act_regs_data_3_6_2_enexo_4 <= act_regs_data_and_2558_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_6_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2690_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_29_enex5
        ) begin
      reg_act_regs_data_0_6_2_enexo_4 <= act_regs_data_and_2690_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_148 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_30_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_148 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_148 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_30_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_148 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_148 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_30_enex5
        ) begin
      reg_act_config_inst_counter_enexo_148 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_6_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2607_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_30_enex5
        ) begin
      reg_act_regs_data_2_6_3_enexo_4 <= act_regs_data_and_2607_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_6_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2559_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_30_enex5
        ) begin
      reg_act_regs_data_3_6_3_enexo_4 <= act_regs_data_and_2559_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_6_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2691_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_30_enex5
        ) begin
      reg_act_regs_data_0_6_3_enexo_4 <= act_regs_data_and_2691_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_6_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2655_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_30_enex5
        ) begin
      reg_act_regs_data_1_6_3_enexo_4 <= act_regs_data_and_2655_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_149 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_31_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_149 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_149 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_31_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_149 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_149 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_31_enex5
        ) begin
      reg_act_config_inst_counter_enexo_149 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_6_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2557_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_31_enex5
        ) begin
      reg_act_regs_data_3_6_1_enexo_4 <= act_regs_data_and_2557_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_6_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2653_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_31_enex5
        ) begin
      reg_act_regs_data_1_6_1_enexo_4 <= act_regs_data_and_2653_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_6_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2605_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_31_enex5
        ) begin
      reg_act_regs_data_2_6_1_enexo_4 <= act_regs_data_and_2605_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_6_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2689_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_31_enex5
        ) begin
      reg_act_regs_data_0_6_1_enexo_4 <= act_regs_data_and_2689_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_150 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_32_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_150 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_150 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_32_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_150 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_150 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_32_enex5
        ) begin
      reg_act_config_inst_counter_enexo_150 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_7_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2687_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_32_enex5
        ) begin
      reg_act_regs_data_0_7_2_enexo_4 <= act_regs_data_and_2687_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_7_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2603_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_32_enex5
        ) begin
      reg_act_regs_data_2_7_2_enexo_4 <= act_regs_data_and_2603_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_7_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2555_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_32_enex5
        ) begin
      reg_act_regs_data_3_7_2_enexo_4 <= act_regs_data_and_2555_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_7_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2651_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_32_enex5
        ) begin
      reg_act_regs_data_1_7_2_enexo_4 <= act_regs_data_and_2651_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_151 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_33_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_151 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_151 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_33_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_151 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_151 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_33_enex5
        ) begin
      reg_act_config_inst_counter_enexo_151 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_7_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2688_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_33_enex5
        ) begin
      reg_act_regs_data_0_7_3_enexo_4 <= act_regs_data_and_2688_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_7_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2652_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_33_enex5
        ) begin
      reg_act_regs_data_1_7_3_enexo_4 <= act_regs_data_and_2652_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_7_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2556_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_33_enex5
        ) begin
      reg_act_regs_data_3_7_3_enexo_4 <= act_regs_data_and_2556_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_7_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2604_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_33_enex5
        ) begin
      reg_act_regs_data_2_7_3_enexo_4 <= act_regs_data_and_2604_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_152 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_34_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_152 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_152 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_34_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_152 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_152 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_34_enex5
        ) begin
      reg_act_config_inst_counter_enexo_152 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_7_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2554_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_34_enex5
        ) begin
      reg_act_regs_data_3_7_1_enexo_4 <= act_regs_data_and_2554_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_7_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2650_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_34_enex5
        ) begin
      reg_act_regs_data_1_7_1_enexo_4 <= act_regs_data_and_2650_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_7_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2686_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_34_enex5
        ) begin
      reg_act_regs_data_0_7_1_enexo_4 <= act_regs_data_and_2686_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_7_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2602_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_34_enex5
        ) begin
      reg_act_regs_data_2_7_1_enexo_4 <= act_regs_data_and_2602_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_153 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_35_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_153 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_153 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_35_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_153 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_153 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_35_enex5
        ) begin
      reg_act_config_inst_counter_enexo_153 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_8_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2684_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_35_enex5
        ) begin
      reg_act_regs_data_0_8_2_enexo_4 <= act_regs_data_and_2684_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_8_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2648_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_35_enex5
        ) begin
      reg_act_regs_data_1_8_2_enexo_4 <= act_regs_data_and_2648_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_8_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2600_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_35_enex5
        ) begin
      reg_act_regs_data_2_8_2_enexo_4 <= act_regs_data_and_2600_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_8_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2552_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_35_enex5
        ) begin
      reg_act_regs_data_3_8_2_enexo_4 <= act_regs_data_and_2552_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_154 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_36_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_154 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_154 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_36_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_154 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_154 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_36_enex5
        ) begin
      reg_act_config_inst_counter_enexo_154 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_8_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2685_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_36_enex5
        ) begin
      reg_act_regs_data_0_8_3_enexo_4 <= act_regs_data_and_2685_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_8_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2601_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_36_enex5
        ) begin
      reg_act_regs_data_2_8_3_enexo_4 <= act_regs_data_and_2601_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_8_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2649_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_36_enex5
        ) begin
      reg_act_regs_data_1_8_3_enexo_4 <= act_regs_data_and_2649_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_8_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2553_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_36_enex5
        ) begin
      reg_act_regs_data_3_8_3_enexo_4 <= act_regs_data_and_2553_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_155 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_37_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_155 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_155 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_37_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_155 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_155 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_37_enex5
        ) begin
      reg_act_config_inst_counter_enexo_155 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_8_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2599_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_37_enex5
        ) begin
      reg_act_regs_data_2_8_1_enexo_4 <= act_regs_data_and_2599_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_8_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2683_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_37_enex5
        ) begin
      reg_act_regs_data_0_8_1_enexo_4 <= act_regs_data_and_2683_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_8_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2551_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_37_enex5
        ) begin
      reg_act_regs_data_3_8_1_enexo_4 <= act_regs_data_and_2551_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_8_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2647_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_37_enex5
        ) begin
      reg_act_regs_data_1_8_1_enexo_4 <= act_regs_data_and_2647_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_156 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_38_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_156 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_156 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_38_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_156 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_156 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_38_enex5
        ) begin
      reg_act_config_inst_counter_enexo_156 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_9_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2681_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_38_enex5
        ) begin
      reg_act_regs_data_0_9_2_enexo_4 <= act_regs_data_and_2681_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_9_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2597_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_38_enex5
        ) begin
      reg_act_regs_data_2_9_2_enexo_4 <= act_regs_data_and_2597_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_9_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2645_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_38_enex5
        ) begin
      reg_act_regs_data_1_9_2_enexo_4 <= act_regs_data_and_2645_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_9_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2549_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_38_enex5
        ) begin
      reg_act_regs_data_3_9_2_enexo_4 <= act_regs_data_and_2549_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_157 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_39_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_157 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_157 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_39_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_157 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_157 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_39_enex5
        ) begin
      reg_act_config_inst_counter_enexo_157 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_9_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2646_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_39_enex5
        ) begin
      reg_act_regs_data_1_9_3_enexo_4 <= act_regs_data_and_2646_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_9_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2682_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_39_enex5
        ) begin
      reg_act_regs_data_0_9_3_enexo_4 <= act_regs_data_and_2682_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_9_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2598_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_39_enex5
        ) begin
      reg_act_regs_data_2_9_3_enexo_4 <= act_regs_data_and_2598_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_9_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2550_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_39_enex5
        ) begin
      reg_act_regs_data_3_9_3_enexo_4 <= act_regs_data_and_2550_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_158 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_40_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_158 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_158 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_40_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_158 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_158 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_40_enex5
        ) begin
      reg_act_config_inst_counter_enexo_158 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_9_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2644_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_40_enex5
        ) begin
      reg_act_regs_data_1_9_1_enexo_4 <= act_regs_data_and_2644_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_9_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2548_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_40_enex5
        ) begin
      reg_act_regs_data_3_9_1_enexo_4 <= act_regs_data_and_2548_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_9_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2680_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_40_enex5
        ) begin
      reg_act_regs_data_0_9_1_enexo_4 <= act_regs_data_and_2680_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_9_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2596_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_40_enex5
        ) begin
      reg_act_regs_data_2_9_1_enexo_4 <= act_regs_data_and_2596_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_159 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_41_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_159 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_159 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_41_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_159 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_159 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_41_enex5
        ) begin
      reg_act_config_inst_counter_enexo_159 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_10_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2642_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_41_enex5
        ) begin
      reg_act_regs_data_1_10_2_enexo_4 <= act_regs_data_and_2642_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_10_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2759_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_41_enex5
        ) begin
      reg_act_regs_data_0_10_2_enexo_4 <= act_regs_data_and_2759_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_10_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2546_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_41_enex5
        ) begin
      reg_act_regs_data_3_10_2_enexo_4 <= act_regs_data_and_2546_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_10_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2594_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_41_enex5
        ) begin
      reg_act_regs_data_2_10_2_enexo_4 <= act_regs_data_and_2594_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_160 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_42_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_160 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_160 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_42_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_160 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_160 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_42_enex5
        ) begin
      reg_act_config_inst_counter_enexo_160 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_10_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2547_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_42_enex5
        ) begin
      reg_act_regs_data_3_10_3_enexo_4 <= act_regs_data_and_2547_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_10_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2760_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_42_enex5
        ) begin
      reg_act_regs_data_0_10_3_enexo_4 <= act_regs_data_and_2760_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_10_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2595_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_42_enex5
        ) begin
      reg_act_regs_data_2_10_3_enexo_4 <= act_regs_data_and_2595_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_10_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2643_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_42_enex5
        ) begin
      reg_act_regs_data_1_10_3_enexo_4 <= act_regs_data_and_2643_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_161 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_43_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_161 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_161 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_43_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_161 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_161 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_43_enex5
        ) begin
      reg_act_config_inst_counter_enexo_161 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_10_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2641_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_43_enex5
        ) begin
      reg_act_regs_data_1_10_1_enexo_4 <= act_regs_data_and_2641_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_10_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2593_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_43_enex5
        ) begin
      reg_act_regs_data_2_10_1_enexo_4 <= act_regs_data_and_2593_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_10_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2545_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_43_enex5
        ) begin
      reg_act_regs_data_3_10_1_enexo_4 <= act_regs_data_and_2545_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_10_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2758_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_43_enex5
        ) begin
      reg_act_regs_data_0_10_1_enexo_4 <= act_regs_data_and_2758_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_162 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_44_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_162 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_162 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_44_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_162 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_162 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_44_enex5
        ) begin
      reg_act_config_inst_counter_enexo_162 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_11_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2591_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_44_enex5
        ) begin
      reg_act_regs_data_2_11_2_enexo_4 <= act_regs_data_and_2591_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_11_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2756_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_44_enex5
        ) begin
      reg_act_regs_data_0_11_2_enexo_4 <= act_regs_data_and_2756_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_11_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2543_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_44_enex5
        ) begin
      reg_act_regs_data_3_11_2_enexo_4 <= act_regs_data_and_2543_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_11_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2639_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_44_enex5
        ) begin
      reg_act_regs_data_1_11_2_enexo_4 <= act_regs_data_and_2639_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_163 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_45_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_163 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_163 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_45_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_163 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_163 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_45_enex5
        ) begin
      reg_act_config_inst_counter_enexo_163 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_11_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2757_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_45_enex5
        ) begin
      reg_act_regs_data_0_11_3_enexo_4 <= act_regs_data_and_2757_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_11_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2640_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_45_enex5
        ) begin
      reg_act_regs_data_1_11_3_enexo_4 <= act_regs_data_and_2640_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_11_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2592_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_45_enex5
        ) begin
      reg_act_regs_data_2_11_3_enexo_4 <= act_regs_data_and_2592_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_11_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2544_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_45_enex5
        ) begin
      reg_act_regs_data_3_11_3_enexo_4 <= act_regs_data_and_2544_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_164 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_46_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_164 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_164 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_46_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_164 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_164 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_46_enex5
        ) begin
      reg_act_config_inst_counter_enexo_164 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_11_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2590_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_46_enex5
        ) begin
      reg_act_regs_data_2_11_1_enexo_4 <= act_regs_data_and_2590_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_11_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2542_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_46_enex5
        ) begin
      reg_act_regs_data_3_11_1_enexo_4 <= act_regs_data_and_2542_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_11_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2755_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_46_enex5
        ) begin
      reg_act_regs_data_0_11_1_enexo_4 <= act_regs_data_and_2755_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_11_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2638_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_46_enex5
        ) begin
      reg_act_regs_data_1_11_1_enexo_4 <= act_regs_data_and_2638_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_165 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_47_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_165 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_165 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_47_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_165 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_12_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2588_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_47_enex5
        ) begin
      reg_act_regs_data_2_12_2_enexo_4 <= act_regs_data_and_2588_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_165 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_47_enex5
        ) begin
      reg_act_config_inst_counter_enexo_165 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_12_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2753_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_47_enex5
        ) begin
      reg_act_regs_data_0_12_2_enexo_4 <= act_regs_data_and_2753_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_12_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2540_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_47_enex5
        ) begin
      reg_act_regs_data_3_12_2_enexo_4 <= act_regs_data_and_2540_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_12_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2636_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_47_enex5
        ) begin
      reg_act_regs_data_1_12_2_enexo_4 <= act_regs_data_and_2636_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_166 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_48_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_166 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_166 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_48_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_166 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_166 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_48_enex5
        ) begin
      reg_act_config_inst_counter_enexo_166 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_12_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2754_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_48_enex5
        ) begin
      reg_act_regs_data_0_12_3_enexo_4 <= act_regs_data_and_2754_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_12_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2589_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_48_enex5
        ) begin
      reg_act_regs_data_2_12_3_enexo_4 <= act_regs_data_and_2589_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_12_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2541_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_48_enex5
        ) begin
      reg_act_regs_data_3_12_3_enexo_4 <= act_regs_data_and_2541_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_12_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2637_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_48_enex5
        ) begin
      reg_act_regs_data_1_12_3_enexo_4 <= act_regs_data_and_2637_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_167 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_49_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_167 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_167 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_49_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_167 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_167 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_49_enex5
        ) begin
      reg_act_config_inst_counter_enexo_167 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_12_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2587_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_49_enex5
        ) begin
      reg_act_regs_data_2_12_1_enexo_4 <= act_regs_data_and_2587_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_12_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2752_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_49_enex5
        ) begin
      reg_act_regs_data_0_12_1_enexo_4 <= act_regs_data_and_2752_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_12_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2635_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_49_enex5
        ) begin
      reg_act_regs_data_1_12_1_enexo_4 <= act_regs_data_and_2635_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_12_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2539_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_49_enex5
        ) begin
      reg_act_regs_data_3_12_1_enexo_4 <= act_regs_data_and_2539_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_13_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2537_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_50_enex5
        ) begin
      reg_act_regs_data_3_13_2_enexo_4 <= act_regs_data_and_2537_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_168 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_50_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_168 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_168 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_50_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_168 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_13_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2750_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_50_enex5
        ) begin
      reg_act_regs_data_0_13_2_enexo_4 <= act_regs_data_and_2750_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_168 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_50_enex5
        ) begin
      reg_act_config_inst_counter_enexo_168 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_13_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2633_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_50_enex5
        ) begin
      reg_act_regs_data_1_13_2_enexo_4 <= act_regs_data_and_2633_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_13_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2585_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_50_enex5
        ) begin
      reg_act_regs_data_2_13_2_enexo_4 <= act_regs_data_and_2585_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_169 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_51_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_169 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_169 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_51_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_169 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_169 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_51_enex5
        ) begin
      reg_act_config_inst_counter_enexo_169 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_13_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2586_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_51_enex5
        ) begin
      reg_act_regs_data_2_13_3_enexo_4 <= act_regs_data_and_2586_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_13_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2538_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_51_enex5
        ) begin
      reg_act_regs_data_3_13_3_enexo_4 <= act_regs_data_and_2538_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_13_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2634_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_51_enex5
        ) begin
      reg_act_regs_data_1_13_3_enexo_4 <= act_regs_data_and_2634_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_13_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2751_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_51_enex5
        ) begin
      reg_act_regs_data_0_13_3_enexo_4 <= act_regs_data_and_2751_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_170 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_52_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_170 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_13_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2632_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_52_enex5
        ) begin
      reg_act_regs_data_1_13_1_enexo_4 <= act_regs_data_and_2632_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_13_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2584_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_52_enex5
        ) begin
      reg_act_regs_data_2_13_1_enexo_4 <= act_regs_data_and_2584_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_170 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_52_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_170 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_170 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_52_enex5
        ) begin
      reg_act_config_inst_counter_enexo_170 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_13_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2749_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_52_enex5
        ) begin
      reg_act_regs_data_0_13_1_enexo_4 <= act_regs_data_and_2749_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_13_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2536_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_52_enex5
        ) begin
      reg_act_regs_data_3_13_1_enexo_4 <= act_regs_data_and_2536_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_171 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_53_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_171 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_14_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2678_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_53_enex5
        ) begin
      reg_act_regs_data_0_14_2_enexo_4 <= act_regs_data_and_2678_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_171 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_53_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_171 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_171 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_53_enex5
        ) begin
      reg_act_config_inst_counter_enexo_171 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_14_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2582_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_53_enex5
        ) begin
      reg_act_regs_data_2_14_2_enexo_4 <= act_regs_data_and_2582_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_14_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2534_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_53_enex5
        ) begin
      reg_act_regs_data_3_14_2_enexo_4 <= act_regs_data_and_2534_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_14_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2630_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_53_enex5
        ) begin
      reg_act_regs_data_1_14_2_enexo_4 <= act_regs_data_and_2630_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_172 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_54_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_172 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_172 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_54_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_172 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_172 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_54_enex5
        ) begin
      reg_act_config_inst_counter_enexo_172 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_14_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2679_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_54_enex5
        ) begin
      reg_act_regs_data_0_14_3_enexo_4 <= act_regs_data_and_2679_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_14_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2583_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_54_enex5
        ) begin
      reg_act_regs_data_2_14_3_enexo_4 <= act_regs_data_and_2583_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_14_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2535_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_54_enex5
        ) begin
      reg_act_regs_data_3_14_3_enexo_4 <= act_regs_data_and_2535_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_14_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2631_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_54_enex5
        ) begin
      reg_act_regs_data_1_14_3_enexo_4 <= act_regs_data_and_2631_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_173 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_55_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_173 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_14_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2629_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_55_enex5
        ) begin
      reg_act_regs_data_1_14_1_enexo_4 <= act_regs_data_and_2629_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_173 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_55_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_173 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_173 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_55_enex5
        ) begin
      reg_act_config_inst_counter_enexo_173 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_14_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2581_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_55_enex5
        ) begin
      reg_act_regs_data_2_14_1_enexo_4 <= act_regs_data_and_2581_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_14_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2533_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_55_enex5
        ) begin
      reg_act_regs_data_3_14_1_enexo_4 <= act_regs_data_and_2533_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_14_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2677_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_55_enex5
        ) begin
      reg_act_regs_data_0_14_1_enexo_4 <= act_regs_data_and_2677_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_174 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_56_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_174 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_174 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_56_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_174 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_174 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_56_enex5
        ) begin
      reg_act_config_inst_counter_enexo_174 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_15_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2531_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_56_enex5
        ) begin
      reg_act_regs_data_3_15_2_enexo_4 <= act_regs_data_and_2531_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_15_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2579_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_56_enex5
        ) begin
      reg_act_regs_data_2_15_2_enexo_4 <= act_regs_data_and_2579_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_15_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2675_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_56_enex5
        ) begin
      reg_act_regs_data_0_15_2_enexo_4 <= act_regs_data_and_2675_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_15_2_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2627_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_56_enex5
        ) begin
      reg_act_regs_data_1_15_2_enexo_4 <= act_regs_data_and_2627_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_175 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_57_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_175 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_175 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_57_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_175 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_15_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2580_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_57_enex5
        ) begin
      reg_act_regs_data_2_15_3_enexo_4 <= act_regs_data_and_2580_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_175 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_57_enex5
        ) begin
      reg_act_config_inst_counter_enexo_175 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_15_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2676_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_57_enex5
        ) begin
      reg_act_regs_data_0_15_3_enexo_4 <= act_regs_data_and_2676_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_15_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2628_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_57_enex5
        ) begin
      reg_act_regs_data_1_15_3_enexo_4 <= act_regs_data_and_2628_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_15_3_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2532_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_57_enex5
        ) begin
      reg_act_regs_data_3_15_3_enexo_4 <= act_regs_data_and_2532_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_176 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_6_for_and_58_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_176 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_176 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_6_for_and_58_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_176 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_176 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_6_for_and_58_enex5
        ) begin
      reg_act_config_inst_counter_enexo_176 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_15_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2674_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_58_enex5
        ) begin
      reg_act_regs_data_0_15_1_enexo_4 <= act_regs_data_and_2674_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_15_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2626_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_58_enex5
        ) begin
      reg_act_regs_data_1_15_1_enexo_4 <= act_regs_data_and_2626_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_15_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2578_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_58_enex5
        ) begin
      reg_act_regs_data_2_15_1_enexo_4 <= act_regs_data_and_2578_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_15_1_enexo_4 <= 1'b1;
    end
    else if ( act_regs_data_and_2530_enex5 | nv_scvector_cctor_nv_scvector_6_for_and_58_enex5
        ) begin
      reg_act_regs_data_3_15_1_enexo_4 <= act_regs_data_and_2530_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2704_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2704_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2704_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2704_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2704_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2704_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2704_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2704_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2704_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2704_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2704_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2704_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2704_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2704_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2704_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2704_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_15_sva_dfm_2_30_26_enexo_1 <= 1'b1;
    end
    else if ( and_2189_tmp | act_regs_data_and_2704_enex5 ) begin
      reg_act_regs_data_3_15_sva_dfm_2_30_26_enexo_1 <= and_2189_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2704_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2704_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_1 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2705_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_1 <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_1 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2705_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_1 <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_1 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2705_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_1 <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_15_sva_dfm_2_25_22_enexo_1 <= 1'b1;
    end
    else if ( and_2061_cse | act_regs_data_and_2705_enex5 ) begin
      reg_act_regs_data_3_15_sva_dfm_2_25_22_enexo_1 <= and_2061_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_1 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2705_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_1 <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_1 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2705_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_1 <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_1 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2705_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_1 <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_1 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2705_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_1 <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_1 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2705_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_1 <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_1 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2705_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_1 <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_1 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2705_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_1 <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_1 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2705_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_1 <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_1 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2705_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_1 <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_1 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2705_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_1 <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_1 <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2705_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_1 <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_1 <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2705_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_1 <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_1 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2705_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_1 <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_1 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2705_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_1 <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_1 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2705_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_1 <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_2 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2706_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_2 <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_2 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2706_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_2 <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_2 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2706_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_2 <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_2 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2706_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_2 <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_2 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2706_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_2 <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_2 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2706_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_2 <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_2 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2706_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_2 <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_2 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2706_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_2 <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_2 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2706_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_2 <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_2 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2706_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_2 <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_2 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2706_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_2 <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_2 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2706_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_2 <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_2 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2706_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_2 <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_2 <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2706_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_2 <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_2 <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2706_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_2 <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_2 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2706_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_2 <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_2 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2706_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_2 <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_15_sva_dfm_2_21_0_enexo_1 <= 1'b1;
    end
    else if ( and_2061_cse | act_regs_data_and_2706_enex5 ) begin
      reg_act_regs_data_3_15_sva_dfm_2_21_0_enexo_1 <= and_2061_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_2 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2706_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_2 <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_3 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2707_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_3 <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_3 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2707_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_3 <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_3 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2707_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_3 <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_3 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2707_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_3 <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_3 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2707_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_3 <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_3 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2707_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_3 <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_3 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2707_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_3 <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_3 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2707_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_3 <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_3 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2707_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_3 <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_3 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2707_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_3 <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_3 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2707_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_3 <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_3 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2707_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_3 <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_3 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2707_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_3 <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_3 <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2707_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_3 <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_3 <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2707_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_3 <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_3 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2707_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_3 <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_14_sva_dfm_2_30_26_enexo_1 <= 1'b1;
    end
    else if ( and_2187_tmp | act_regs_data_and_2707_enex5 ) begin
      reg_act_regs_data_3_14_sva_dfm_2_30_26_enexo_1 <= and_2187_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_3 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2707_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_3 <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_3 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2707_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_3 <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_4 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2708_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_4 <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_4 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2708_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_4 <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_4 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2708_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_4 <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_14_sva_dfm_2_25_22_enexo_1 <= 1'b1;
    end
    else if ( and_2059_cse | act_regs_data_and_2708_enex5 ) begin
      reg_act_regs_data_3_14_sva_dfm_2_25_22_enexo_1 <= and_2059_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_4 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2708_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_4 <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_4 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2708_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_4 <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_4 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2708_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_4 <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_4 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2708_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_4 <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_4 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2708_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_4 <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_4 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2708_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_4 <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_4 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2708_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_4 <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_4 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2708_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_4 <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_4 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2708_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_4 <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_4 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2708_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_4 <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_4 <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2708_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_4 <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_4 <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2708_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_4 <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_4 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2708_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_4 <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_4 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2708_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_4 <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_4 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2708_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_4 <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_5 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2709_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_5 <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_5 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2709_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_5 <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_5 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2709_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_5 <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_5 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2709_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_5 <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_5 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2709_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_5 <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_5 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2709_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_5 <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_5 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2709_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_5 <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_5 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2709_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_5 <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_5 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2709_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_5 <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_5 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2709_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_5 <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_5 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2709_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_5 <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_5 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2709_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_5 <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_5 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2709_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_5 <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_5 <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2709_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_5 <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_5 <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2709_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_5 <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_5 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2709_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_5 <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_5 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2709_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_5 <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_14_sva_dfm_2_21_0_enexo_1 <= 1'b1;
    end
    else if ( and_2059_cse | act_regs_data_and_2709_enex5 ) begin
      reg_act_regs_data_3_14_sva_dfm_2_21_0_enexo_1 <= and_2059_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_5 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2709_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_5 <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_6 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2710_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_6 <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_6 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2710_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_6 <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_6 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2710_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_6 <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_6 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2710_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_6 <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_6 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2710_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_6 <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_6 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2710_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_6 <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_6 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2710_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_6 <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_6 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2710_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_6 <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_6 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2710_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_6 <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_6 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2710_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_6 <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_6 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2710_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_6 <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_6 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2710_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_6 <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_6 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2710_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_6 <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_6 <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2710_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_6 <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_6 <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2710_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_6 <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_6 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2710_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_6 <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_13_sva_dfm_2_30_26_enexo_1 <= 1'b1;
    end
    else if ( and_2185_tmp | act_regs_data_and_2710_enex5 ) begin
      reg_act_regs_data_3_13_sva_dfm_2_30_26_enexo_1 <= and_2185_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_6 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2710_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_6 <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_6 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2710_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_6 <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_7 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2711_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_7 <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_7 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2711_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_7 <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_7 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2711_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_7 <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_13_sva_dfm_2_25_22_enexo_1 <= 1'b1;
    end
    else if ( and_2057_cse | act_regs_data_and_2711_enex5 ) begin
      reg_act_regs_data_3_13_sva_dfm_2_25_22_enexo_1 <= and_2057_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_7 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2711_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_7 <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_7 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2711_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_7 <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_7 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2711_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_7 <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_7 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2711_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_7 <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_7 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2711_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_7 <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_7 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2711_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_7 <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_7 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2711_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_7 <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_7 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2711_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_7 <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_7 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2711_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_7 <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_7 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2711_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_7 <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_7 <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2711_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_7 <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_7 <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2711_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_7 <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_7 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2711_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_7 <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_7 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2711_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_7 <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_7 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2711_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_7 <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_8 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2712_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_8 <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_8 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2712_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_8 <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_8 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2712_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_8 <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_8 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2712_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_8 <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_8 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2712_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_8 <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_8 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2712_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_8 <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_8 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2712_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_8 <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_8 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2712_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_8 <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_8 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2712_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_8 <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_8 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2712_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_8 <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_8 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2712_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_8 <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_8 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2712_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_8 <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_8 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2712_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_8 <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_8 <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2712_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_8 <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_8 <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2712_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_8 <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_8 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2712_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_8 <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_8 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2712_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_8 <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_13_sva_dfm_2_21_0_enexo_1 <= 1'b1;
    end
    else if ( and_2057_cse | act_regs_data_and_2712_enex5 ) begin
      reg_act_regs_data_3_13_sva_dfm_2_21_0_enexo_1 <= and_2057_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_8 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2712_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_8 <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_9 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2713_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_9 <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_9 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2713_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_9 <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_9 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2713_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_9 <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_9 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2713_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_9 <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_9 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2713_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_9 <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_9 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2713_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_9 <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_9 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2713_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_9 <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_9 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2713_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_9 <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_9 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2713_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_9 <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_9 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2713_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_9 <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_9 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2713_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_9 <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_9 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2713_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_9 <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_9 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2713_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_9 <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_9 <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2713_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_9 <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_9 <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2713_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_9 <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_9 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2713_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_9 <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_12_sva_dfm_2_30_26_enexo_1 <= 1'b1;
    end
    else if ( and_2183_tmp | act_regs_data_and_2713_enex5 ) begin
      reg_act_regs_data_3_12_sva_dfm_2_30_26_enexo_1 <= and_2183_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_9 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2713_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_9 <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_9 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2713_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_9 <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_10 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2714_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_10 <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_10 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2714_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_10 <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_10 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2714_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_10 <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_12_sva_dfm_2_25_22_enexo_1 <= 1'b1;
    end
    else if ( and_2055_cse | act_regs_data_and_2714_enex5 ) begin
      reg_act_regs_data_3_12_sva_dfm_2_25_22_enexo_1 <= and_2055_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_10 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2714_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_10 <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_10 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2714_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_10 <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_10 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2714_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_10 <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_10 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2714_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_10 <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_10 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2714_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_10 <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_10 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2714_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_10 <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_10 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2714_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_10 <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_10 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2714_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_10 <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_10 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2714_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_10 <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_10 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2714_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_10 <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_10 <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2714_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_10 <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_10 <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2714_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_10 <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_10 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2714_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_10 <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_10 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2714_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_10 <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_10 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2714_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_10 <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_11 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2715_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_11 <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_11 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2715_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_11 <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_11 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2715_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_11 <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_11 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2715_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_11 <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_11 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2715_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_11 <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_11 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2715_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_11 <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_11 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2715_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_11 <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_11 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2715_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_11 <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_11 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2715_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_11 <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_11 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2715_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_11 <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_11 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2715_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_11 <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_11 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2715_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_11 <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_11 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2715_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_11 <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_11 <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2715_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_11 <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_11 <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2715_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_11 <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_11 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2715_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_11 <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_11 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2715_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_11 <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_12_sva_dfm_2_21_0_enexo_1 <= 1'b1;
    end
    else if ( and_2055_cse | act_regs_data_and_2715_enex5 ) begin
      reg_act_regs_data_3_12_sva_dfm_2_21_0_enexo_1 <= and_2055_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_11 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2715_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_11 <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_12 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2716_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_12 <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_12 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2716_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_12 <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_12 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2716_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_12 <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_12 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2716_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_12 <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_12 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2716_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_12 <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_12 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2716_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_12 <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_12 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2716_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_12 <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_12 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2716_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_12 <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_12 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2716_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_12 <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_12 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2716_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_12 <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_12 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2716_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_12 <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_12 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2716_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_12 <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_12 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2716_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_12 <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_12 <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2716_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_12 <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_12 <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2716_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_12 <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_12 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2716_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_12 <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_11_sva_dfm_2_30_26_enexo_1 <= 1'b1;
    end
    else if ( and_2181_tmp | act_regs_data_and_2716_enex5 ) begin
      reg_act_regs_data_3_11_sva_dfm_2_30_26_enexo_1 <= and_2181_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_12 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2716_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_12 <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_12 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2716_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_12 <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_13 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2717_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_13 <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_13 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2717_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_13 <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_13 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2717_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_13 <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_11_sva_dfm_2_25_22_enexo_1 <= 1'b1;
    end
    else if ( and_2053_cse | act_regs_data_and_2717_enex5 ) begin
      reg_act_regs_data_3_11_sva_dfm_2_25_22_enexo_1 <= and_2053_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_13 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2717_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_13 <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_13 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2717_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_13 <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_13 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2717_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_13 <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_13 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2717_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_13 <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_13 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2717_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_13 <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_13 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2717_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_13 <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_13 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2717_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_13 <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_13 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2717_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_13 <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_13 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2717_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_13 <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_13 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2717_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_13 <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_13 <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2717_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_13 <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_13 <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2717_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_13 <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_13 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2717_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_13 <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_13 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2717_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_13 <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_13 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2717_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_13 <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_14 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2718_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_14 <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_14 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2718_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_14 <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_14 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2718_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_14 <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_14 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2718_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_14 <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_14 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2718_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_14 <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_14 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2718_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_14 <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_14 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2718_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_14 <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_14 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2718_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_14 <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_14 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2718_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_14 <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_14 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2718_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_14 <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_14 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2718_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_14 <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_14 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2718_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_14 <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_14 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2718_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_14 <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_14 <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2718_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_14 <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_14 <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2718_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_14 <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_14 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2718_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_14 <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_14 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2718_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_14 <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_11_sva_dfm_2_21_0_enexo_1 <= 1'b1;
    end
    else if ( and_2053_cse | act_regs_data_and_2718_enex5 ) begin
      reg_act_regs_data_3_11_sva_dfm_2_21_0_enexo_1 <= and_2053_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_14 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2718_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_14 <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_15 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2719_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_15 <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_15 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2719_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_15 <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_15 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2719_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_15 <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_15 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2719_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_15 <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_15 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2719_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_15 <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_15 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2719_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_15 <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_15 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2719_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_15 <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_15 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2719_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_15 <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_15 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2719_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_15 <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_15 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2719_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_15 <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_15 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2719_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_15 <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_15 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2719_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_15 <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_15 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2719_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_15 <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_15 <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2719_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_15 <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_15 <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2719_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_15 <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_15 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2719_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_15 <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_10_sva_dfm_2_30_26_enexo_1 <= 1'b1;
    end
    else if ( and_2179_tmp | act_regs_data_and_2719_enex5 ) begin
      reg_act_regs_data_3_10_sva_dfm_2_30_26_enexo_1 <= and_2179_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_15 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2719_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_15 <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_15 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2719_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_15 <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_16 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2720_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_16 <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_16 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2720_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_16 <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_16 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2720_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_16 <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_10_sva_dfm_2_25_22_enexo_1 <= 1'b1;
    end
    else if ( and_2051_cse | act_regs_data_and_2720_enex5 ) begin
      reg_act_regs_data_3_10_sva_dfm_2_25_22_enexo_1 <= and_2051_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_16 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2720_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_16 <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_16 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2720_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_16 <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_16 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2720_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_16 <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_16 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2720_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_16 <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_16 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2720_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_16 <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_16 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2720_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_16 <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_16 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2720_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_16 <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_16 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2720_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_16 <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_16 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2720_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_16 <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_16 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2720_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_16 <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_16 <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2720_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_16 <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_16 <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2720_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_16 <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_16 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2720_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_16 <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_16 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2720_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_16 <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_16 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2720_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_16 <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_17 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2721_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_17 <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_17 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2721_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_17 <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_17 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2721_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_17 <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_17 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2721_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_17 <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_17 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2721_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_17 <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_17 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2721_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_17 <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_17 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2721_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_17 <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_17 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2721_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_17 <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_17 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2721_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_17 <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_17 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2721_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_17 <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_17 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2721_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_17 <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_17 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2721_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_17 <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_17 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2721_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_17 <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_17 <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2721_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_17 <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_17 <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2721_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_17 <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_17 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2721_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_17 <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_17 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2721_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_17 <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_10_sva_dfm_2_21_0_enexo_1 <= 1'b1;
    end
    else if ( and_2051_cse | act_regs_data_and_2721_enex5 ) begin
      reg_act_regs_data_3_10_sva_dfm_2_21_0_enexo_1 <= and_2051_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_17 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2721_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_17 <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_18 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2722_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_18 <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_18 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2722_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_18 <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_18 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2722_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_18 <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_18 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2722_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_18 <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_18 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2722_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_18 <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_18 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2722_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_18 <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_18 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2722_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_18 <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_18 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2722_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_18 <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_18 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2722_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_18 <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_18 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2722_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_18 <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_18 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2722_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_18 <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_18 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2722_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_18 <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_18 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2722_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_18 <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_18 <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2722_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_18 <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_18 <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2722_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_18 <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_18 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2722_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_18 <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_9_sva_dfm_2_30_26_enexo_1 <= 1'b1;
    end
    else if ( and_2177_tmp | act_regs_data_and_2722_enex5 ) begin
      reg_act_regs_data_3_9_sva_dfm_2_30_26_enexo_1 <= and_2177_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_18 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2722_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_18 <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_18 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2722_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_18 <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_19 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2723_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_19 <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_19 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2723_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_19 <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_19 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2723_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_19 <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_9_sva_dfm_2_25_22_enexo_1 <= 1'b1;
    end
    else if ( and_2049_cse | act_regs_data_and_2723_enex5 ) begin
      reg_act_regs_data_3_9_sva_dfm_2_25_22_enexo_1 <= and_2049_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_19 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2723_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_19 <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_19 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2723_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_19 <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_19 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2723_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_19 <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_19 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2723_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_19 <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_19 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2723_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_19 <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_19 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2723_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_19 <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_19 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2723_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_19 <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_19 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2723_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_19 <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_19 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2723_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_19 <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_19 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2723_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_19 <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_19 <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2723_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_19 <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_19 <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2723_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_19 <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_19 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2723_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_19 <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_19 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2723_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_19 <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_19 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2723_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_19 <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_20 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2724_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_20 <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_20 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2724_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_20 <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_20 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2724_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_20 <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_20 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2724_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_20 <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_20 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2724_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_20 <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_20 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2724_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_20 <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_20 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2724_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_20 <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_20 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2724_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_20 <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_20 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2724_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_20 <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_20 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2724_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_20 <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_20 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2724_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_20 <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_20 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2724_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_20 <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_20 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2724_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_20 <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_20 <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2724_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_20 <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_20 <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2724_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_20 <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_20 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2724_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_20 <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_20 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2724_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_20 <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_9_sva_dfm_2_21_0_enexo_1 <= 1'b1;
    end
    else if ( and_2049_cse | act_regs_data_and_2724_enex5 ) begin
      reg_act_regs_data_3_9_sva_dfm_2_21_0_enexo_1 <= and_2049_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_20 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2724_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_20 <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_21 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2725_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_21 <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_21 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2725_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_21 <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_21 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2725_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_21 <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_21 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2725_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_21 <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_21 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2725_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_21 <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_21 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2725_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_21 <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_21 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2725_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_21 <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_21 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2725_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_21 <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_21 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2725_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_21 <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_21 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2725_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_21 <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_21 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2725_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_21 <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_21 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2725_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_21 <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_21 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2725_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_21 <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_21 <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2725_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_21 <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_21 <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2725_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_21 <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_21 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2725_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_21 <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_8_sva_dfm_2_30_26_enexo_1 <= 1'b1;
    end
    else if ( and_2175_tmp | act_regs_data_and_2725_enex5 ) begin
      reg_act_regs_data_3_8_sva_dfm_2_30_26_enexo_1 <= and_2175_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_21 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2725_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_21 <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_21 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2725_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_21 <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_22 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2726_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_22 <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_22 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2726_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_22 <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_22 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2726_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_22 <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_8_sva_dfm_2_25_22_enexo_1 <= 1'b1;
    end
    else if ( and_2047_cse | act_regs_data_and_2726_enex5 ) begin
      reg_act_regs_data_3_8_sva_dfm_2_25_22_enexo_1 <= and_2047_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_22 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2726_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_22 <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_22 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2726_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_22 <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_22 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2726_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_22 <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_22 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2726_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_22 <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_22 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2726_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_22 <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_22 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2726_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_22 <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_22 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2726_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_22 <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_22 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2726_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_22 <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_22 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2726_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_22 <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_22 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2726_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_22 <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_22 <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2726_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_22 <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_22 <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2726_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_22 <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_22 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2726_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_22 <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_22 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2726_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_22 <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_22 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2726_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_22 <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_23 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2727_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_23 <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_23 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2727_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_23 <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_23 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2727_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_23 <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_23 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2727_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_23 <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_23 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2727_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_23 <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_23 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2727_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_23 <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_23 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2727_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_23 <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_23 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2727_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_23 <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_23 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2727_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_23 <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_23 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2727_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_23 <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_23 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2727_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_23 <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_23 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2727_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_23 <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_23 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2727_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_23 <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_23 <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2727_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_23 <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_23 <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2727_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_23 <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_23 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2727_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_23 <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_23 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2727_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_23 <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_8_sva_dfm_2_21_0_enexo_1 <= 1'b1;
    end
    else if ( and_2047_cse | act_regs_data_and_2727_enex5 ) begin
      reg_act_regs_data_3_8_sva_dfm_2_21_0_enexo_1 <= and_2047_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_23 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2727_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_23 <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_24 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2728_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_24 <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_24 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2728_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_24 <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_24 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2728_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_24 <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_24 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2728_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_24 <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_24 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2728_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_24 <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_24 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2728_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_24 <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_24 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2728_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_24 <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_24 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2728_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_24 <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_24 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2728_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_24 <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_24 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2728_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_24 <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_24 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2728_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_24 <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_24 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2728_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_24 <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_24 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2728_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_24 <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_24 <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2728_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_24 <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_24 <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2728_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_24 <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_24 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2728_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_24 <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_7_sva_dfm_2_30_26_enexo_1 <= 1'b1;
    end
    else if ( and_2173_tmp | act_regs_data_and_2728_enex5 ) begin
      reg_act_regs_data_3_7_sva_dfm_2_30_26_enexo_1 <= and_2173_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_24 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2728_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_24 <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_24 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2728_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_24 <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_25 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2729_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_25 <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_25 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2729_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_25 <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_25 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2729_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_25 <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_7_sva_dfm_2_25_22_enexo_1 <= 1'b1;
    end
    else if ( and_2045_cse | act_regs_data_and_2729_enex5 ) begin
      reg_act_regs_data_3_7_sva_dfm_2_25_22_enexo_1 <= and_2045_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_25 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2729_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_25 <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_25 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2729_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_25 <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_25 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2729_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_25 <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_25 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2729_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_25 <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_25 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2729_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_25 <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_25 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2729_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_25 <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_25 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2729_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_25 <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_25 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2729_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_25 <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_25 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2729_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_25 <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_25 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2729_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_25 <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_25 <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2729_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_25 <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_25 <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2729_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_25 <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_25 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2729_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_25 <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_25 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2729_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_25 <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_25 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2729_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_25 <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_26 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2730_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_26 <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_26 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2730_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_26 <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_26 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2730_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_26 <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_26 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2730_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_26 <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_26 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2730_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_26 <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_26 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2730_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_26 <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_26 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2730_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_26 <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_26 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2730_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_26 <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_26 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2730_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_26 <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_26 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2730_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_26 <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_26 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2730_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_26 <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_26 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2730_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_26 <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_26 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2730_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_26 <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_26 <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2730_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_26 <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_26 <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2730_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_26 <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_26 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2730_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_26 <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_26 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2730_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_26 <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_7_sva_dfm_2_21_0_enexo_1 <= 1'b1;
    end
    else if ( and_2045_cse | act_regs_data_and_2730_enex5 ) begin
      reg_act_regs_data_3_7_sva_dfm_2_21_0_enexo_1 <= and_2045_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_26 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2730_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_26 <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_27 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2731_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_27 <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_27 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2731_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_27 <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_27 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2731_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_27 <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_27 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2731_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_27 <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_27 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2731_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_27 <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_27 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2731_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_27 <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_27 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2731_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_27 <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_27 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2731_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_27 <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_27 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2731_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_27 <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_27 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2731_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_27 <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_27 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2731_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_27 <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_27 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2731_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_27 <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_27 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2731_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_27 <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_27 <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2731_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_27 <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_27 <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2731_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_27 <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_27 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2731_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_27 <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_6_sva_dfm_2_30_26_enexo_1 <= 1'b1;
    end
    else if ( and_2171_tmp | act_regs_data_and_2731_enex5 ) begin
      reg_act_regs_data_3_6_sva_dfm_2_30_26_enexo_1 <= and_2171_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_27 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2731_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_27 <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_27 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2731_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_27 <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_28 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2732_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_28 <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_28 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2732_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_28 <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_28 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2732_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_28 <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_6_sva_dfm_2_25_22_enexo_1 <= 1'b1;
    end
    else if ( and_2043_cse | act_regs_data_and_2732_enex5 ) begin
      reg_act_regs_data_3_6_sva_dfm_2_25_22_enexo_1 <= and_2043_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_28 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2732_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_28 <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_28 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2732_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_28 <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_28 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2732_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_28 <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_28 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2732_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_28 <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_28 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2732_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_28 <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_28 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2732_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_28 <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_28 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2732_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_28 <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_28 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2732_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_28 <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_28 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2732_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_28 <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_28 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2732_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_28 <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_28 <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2732_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_28 <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_28 <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2732_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_28 <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_28 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2732_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_28 <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_28 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2732_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_28 <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_28 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2732_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_28 <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_29 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2733_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_29 <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_29 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2733_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_29 <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_29 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2733_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_29 <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_29 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2733_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_29 <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_29 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2733_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_29 <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_29 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2733_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_29 <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_29 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2733_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_29 <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_29 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2733_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_29 <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_29 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2733_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_29 <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_29 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2733_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_29 <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_29 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2733_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_29 <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_29 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2733_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_29 <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_29 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2733_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_29 <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_29 <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2733_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_29 <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_29 <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2733_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_29 <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_29 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2733_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_29 <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_29 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2733_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_29 <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_6_sva_dfm_2_21_0_enexo_1 <= 1'b1;
    end
    else if ( and_2043_cse | act_regs_data_and_2733_enex5 ) begin
      reg_act_regs_data_3_6_sva_dfm_2_21_0_enexo_1 <= and_2043_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_29 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2733_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_29 <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_30 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2734_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_30 <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_30 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2734_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_30 <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_30 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2734_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_30 <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_30 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2734_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_30 <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_30 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2734_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_30 <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_30 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2734_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_30 <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_30 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2734_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_30 <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_30 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2734_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_30 <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_30 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2734_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_30 <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_30 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2734_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_30 <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_30 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2734_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_30 <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_30 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2734_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_30 <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_30 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2734_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_30 <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_30 <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2734_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_30 <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_30 <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2734_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_30 <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_30 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2734_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_30 <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_5_sva_dfm_2_30_26_enexo_1 <= 1'b1;
    end
    else if ( and_2169_tmp | act_regs_data_and_2734_enex5 ) begin
      reg_act_regs_data_3_5_sva_dfm_2_30_26_enexo_1 <= and_2169_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_30 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2734_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_30 <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_30 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2734_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_30 <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_31 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2735_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_31 <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_31 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2735_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_31 <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_31 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2735_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_31 <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_5_sva_dfm_2_25_22_enexo_1 <= 1'b1;
    end
    else if ( and_2041_cse | act_regs_data_and_2735_enex5 ) begin
      reg_act_regs_data_3_5_sva_dfm_2_25_22_enexo_1 <= and_2041_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_31 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2735_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_31 <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_31 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2735_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_31 <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_31 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2735_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_31 <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_31 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2735_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_31 <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_31 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2735_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_31 <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_31 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2735_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_31 <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_31 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2735_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_31 <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_31 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2735_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_31 <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_31 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2735_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_31 <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_31 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2735_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_31 <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_31 <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2735_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_31 <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_31 <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2735_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_31 <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_31 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2735_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_31 <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_31 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2735_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_31 <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_31 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2735_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_31 <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_32 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2736_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_32 <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_32 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2736_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_32 <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_32 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2736_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_32 <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_32 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2736_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_32 <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_32 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2736_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_32 <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_32 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2736_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_32 <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_32 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2736_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_32 <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_32 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2736_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_32 <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_32 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2736_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_32 <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_32 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2736_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_32 <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_32 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2736_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_32 <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_32 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2736_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_32 <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_32 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2736_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_32 <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_32 <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2736_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_32 <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_32 <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2736_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_32 <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_32 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2736_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_32 <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_32 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2736_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_32 <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_5_sva_dfm_2_21_0_enexo_1 <= 1'b1;
    end
    else if ( and_2041_cse | act_regs_data_and_2736_enex5 ) begin
      reg_act_regs_data_3_5_sva_dfm_2_21_0_enexo_1 <= and_2041_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_32 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2736_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_32 <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_33 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2737_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_33 <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_33 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2737_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_33 <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_33 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2737_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_33 <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_33 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2737_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_33 <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_33 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2737_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_33 <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_33 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2737_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_33 <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_33 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2737_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_33 <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_33 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2737_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_33 <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_33 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2737_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_33 <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_33 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2737_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_33 <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_33 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2737_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_33 <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_33 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2737_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_33 <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_33 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2737_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_33 <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_33 <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2737_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_33 <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_33 <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2737_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_33 <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_33 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2737_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_33 <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_4_sva_dfm_2_30_26_enexo_1 <= 1'b1;
    end
    else if ( and_2167_tmp | act_regs_data_and_2737_enex5 ) begin
      reg_act_regs_data_3_4_sva_dfm_2_30_26_enexo_1 <= and_2167_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_33 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2737_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_33 <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_33 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2737_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_33 <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_34 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2738_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_34 <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_34 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2738_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_34 <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_34 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2738_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_34 <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_4_sva_dfm_2_25_22_enexo_1 <= 1'b1;
    end
    else if ( and_2039_cse | act_regs_data_and_2738_enex5 ) begin
      reg_act_regs_data_3_4_sva_dfm_2_25_22_enexo_1 <= and_2039_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_34 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2738_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_34 <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_34 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2738_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_34 <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_34 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2738_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_34 <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_34 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2738_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_34 <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_34 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2738_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_34 <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_34 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2738_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_34 <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_34 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2738_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_34 <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_34 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2738_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_34 <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_34 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2738_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_34 <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_34 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2738_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_34 <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_34 <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2738_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_34 <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_34 <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2738_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_34 <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_34 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2738_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_34 <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_34 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2738_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_34 <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_34 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2738_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_34 <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_35 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2739_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_35 <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_35 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2739_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_35 <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_35 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2739_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_35 <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_35 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2739_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_35 <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_35 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2739_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_35 <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_35 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2739_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_35 <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_35 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2739_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_35 <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_35 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2739_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_35 <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_35 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2739_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_35 <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_35 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2739_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_35 <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_35 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2739_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_35 <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_35 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2739_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_35 <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_35 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2739_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_35 <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_35 <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2739_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_35 <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_35 <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2739_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_35 <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_35 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2739_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_35 <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_35 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2739_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_35 <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_4_sva_dfm_2_21_0_enexo_1 <= 1'b1;
    end
    else if ( and_2039_cse | act_regs_data_and_2739_enex5 ) begin
      reg_act_regs_data_3_4_sva_dfm_2_21_0_enexo_1 <= and_2039_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_35 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2739_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_35 <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_36 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2740_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_36 <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_36 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2740_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_36 <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_36 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2740_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_36 <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_36 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2740_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_36 <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_36 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2740_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_36 <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_36 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2740_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_36 <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_36 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2740_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_36 <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_36 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2740_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_36 <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_36 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2740_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_36 <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_36 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2740_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_36 <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_36 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2740_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_36 <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_36 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2740_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_36 <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_36 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2740_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_36 <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_36 <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2740_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_36 <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_36 <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2740_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_36 <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_36 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2740_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_36 <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_3_sva_dfm_2_30_26_enexo_1 <= 1'b1;
    end
    else if ( and_2165_tmp | act_regs_data_and_2740_enex5 ) begin
      reg_act_regs_data_3_3_sva_dfm_2_30_26_enexo_1 <= and_2165_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_36 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2740_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_36 <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_36 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2740_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_36 <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_37 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2741_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_37 <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_37 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2741_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_37 <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_37 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2741_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_37 <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_3_sva_dfm_2_25_22_enexo_1 <= 1'b1;
    end
    else if ( and_2037_cse | act_regs_data_and_2741_enex5 ) begin
      reg_act_regs_data_3_3_sva_dfm_2_25_22_enexo_1 <= and_2037_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_37 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2741_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_37 <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_37 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2741_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_37 <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_37 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2741_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_37 <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_37 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2741_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_37 <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_37 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2741_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_37 <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_37 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2741_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_37 <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_37 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2741_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_37 <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_37 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2741_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_37 <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_37 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2741_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_37 <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_37 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2741_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_37 <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_37 <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2741_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_37 <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_37 <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2741_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_37 <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_37 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2741_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_37 <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_37 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2741_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_37 <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_37 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2741_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_37 <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_38 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2742_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_38 <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_38 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2742_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_38 <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_38 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2742_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_38 <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_38 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2742_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_38 <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_38 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2742_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_38 <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_38 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2742_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_38 <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_38 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2742_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_38 <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_38 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2742_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_38 <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_38 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2742_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_38 <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_38 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2742_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_38 <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_38 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2742_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_38 <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_38 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2742_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_38 <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_38 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2742_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_38 <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_38 <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2742_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_38 <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_38 <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2742_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_38 <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_38 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2742_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_38 <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_38 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2742_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_38 <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_3_sva_dfm_2_21_0_enexo_1 <= 1'b1;
    end
    else if ( and_2037_cse | act_regs_data_and_2742_enex5 ) begin
      reg_act_regs_data_3_3_sva_dfm_2_21_0_enexo_1 <= and_2037_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_38 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2742_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_38 <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_39 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2743_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_39 <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_39 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2743_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_39 <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_39 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2743_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_39 <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_39 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2743_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_39 <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_39 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2743_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_39 <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_39 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2743_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_39 <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_39 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2743_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_39 <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_39 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2743_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_39 <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_39 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2743_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_39 <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_39 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2743_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_39 <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_39 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2743_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_39 <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_39 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2743_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_39 <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_39 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2743_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_39 <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_39 <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2743_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_39 <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_39 <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2743_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_39 <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_39 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2743_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_39 <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_2_sva_dfm_2_30_26_enexo_1 <= 1'b1;
    end
    else if ( and_2163_tmp | act_regs_data_and_2743_enex5 ) begin
      reg_act_regs_data_3_2_sva_dfm_2_30_26_enexo_1 <= and_2163_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_39 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2743_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_39 <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_39 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2743_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_39 <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_40 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2744_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_40 <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_40 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2744_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_40 <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_40 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2744_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_40 <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_2_sva_dfm_2_25_22_enexo_1 <= 1'b1;
    end
    else if ( and_2035_cse | act_regs_data_and_2744_enex5 ) begin
      reg_act_regs_data_3_2_sva_dfm_2_25_22_enexo_1 <= and_2035_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_40 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2744_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_40 <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_40 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2744_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_40 <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_40 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2744_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_40 <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_40 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2744_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_40 <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_40 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2744_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_40 <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_40 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2744_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_40 <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_40 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2744_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_40 <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_40 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2744_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_40 <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_40 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2744_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_40 <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_40 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2744_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_40 <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_40 <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2744_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_40 <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_40 <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2744_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_40 <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_40 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2744_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_40 <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_40 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2744_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_40 <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_40 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2744_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_40 <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_41 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2745_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_41 <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_41 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2745_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_41 <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_41 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2745_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_41 <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_41 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2745_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_41 <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_41 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2745_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_41 <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_41 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2745_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_41 <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_41 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2745_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_41 <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_41 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2745_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_41 <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_41 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2745_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_41 <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_41 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2745_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_41 <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_41 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2745_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_41 <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_41 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2745_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_41 <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_41 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2745_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_41 <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_41 <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2745_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_41 <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_41 <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2745_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_41 <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_41 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2745_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_41 <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_41 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2745_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_41 <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_2_sva_dfm_2_21_0_enexo_1 <= 1'b1;
    end
    else if ( and_2035_cse | act_regs_data_and_2745_enex5 ) begin
      reg_act_regs_data_3_2_sva_dfm_2_21_0_enexo_1 <= and_2035_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_41 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2745_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_41 <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_42 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2746_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_42 <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_42 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2746_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_42 <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_42 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2746_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_42 <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_42 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2746_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_42 <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_42 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2746_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_42 <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_42 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2746_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_42 <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_42 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2746_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_42 <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_42 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2746_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_42 <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_42 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2746_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_42 <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_42 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2746_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_42 <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_42 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2746_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_42 <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_42 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2746_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_42 <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_42 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2746_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_42 <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_42 <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2746_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_42 <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_42 <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2746_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_42 <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_42 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2746_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_42 <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_1_sva_dfm_2_30_26_enexo_1 <= 1'b1;
    end
    else if ( and_2161_tmp | act_regs_data_and_2746_enex5 ) begin
      reg_act_regs_data_3_1_sva_dfm_2_30_26_enexo_1 <= and_2161_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_42 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2746_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_42 <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_42 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2746_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_42 <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_43 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2747_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_43 <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_43 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2747_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_43 <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_43 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2747_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_43 <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_1_sva_dfm_2_25_22_enexo_1 <= 1'b1;
    end
    else if ( and_2033_cse | act_regs_data_and_2747_enex5 ) begin
      reg_act_regs_data_3_1_sva_dfm_2_25_22_enexo_1 <= and_2033_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_43 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2747_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_43 <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_43 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2747_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_43 <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_43 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2747_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_43 <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_43 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2747_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_43 <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_43 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2747_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_43 <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_43 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2747_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_43 <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_43 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2747_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_43 <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_43 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2747_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_43 <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_43 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2747_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_43 <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_43 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2747_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_43 <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_43 <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2747_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_43 <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_43 <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2747_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_43 <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_43 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2747_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_43 <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_43 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2747_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_43 <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_43 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2747_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_43 <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_44 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_21_enex5 | act_regs_data_and_2748_enex5
        ) begin
      reg_act_port_read_out_data_0_5_sva_dfm_enexo_44 <= act_port_read_out_data_and_21_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_44 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_22_enex5 | act_regs_data_and_2748_enex5
        ) begin
      reg_act_port_read_out_data_0_6_sva_dfm_enexo_44 <= act_port_read_out_data_and_22_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_44 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_29_enex5 | act_regs_data_and_2748_enex5
        ) begin
      reg_act_port_read_out_data_0_13_sva_dfm_enexo_44 <= act_port_read_out_data_and_29_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_44 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_26_enex5 | act_regs_data_and_2748_enex5
        ) begin
      reg_act_port_read_out_data_0_10_sva_dfm_enexo_44 <= act_port_read_out_data_and_26_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_44 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_27_enex5 | act_regs_data_and_2748_enex5
        ) begin
      reg_act_port_read_out_data_0_11_sva_dfm_enexo_44 <= act_port_read_out_data_and_27_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_44 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_31_enex5 | act_regs_data_and_2748_enex5
        ) begin
      reg_act_port_read_out_data_0_15_sva_dfm_enexo_44 <= act_port_read_out_data_and_31_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_44 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_23_enex5 | act_regs_data_and_2748_enex5
        ) begin
      reg_act_port_read_out_data_0_7_sva_dfm_enexo_44 <= act_port_read_out_data_and_23_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_44 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_24_enex5 | act_regs_data_and_2748_enex5
        ) begin
      reg_act_port_read_out_data_0_8_sva_dfm_enexo_44 <= act_port_read_out_data_and_24_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_44 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_16_enex5 | act_regs_data_and_2748_enex5
        ) begin
      reg_act_port_read_out_data_0_0_sva_dfm_enexo_44 <= act_port_read_out_data_and_16_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_44 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_28_enex5 | act_regs_data_and_2748_enex5
        ) begin
      reg_act_port_read_out_data_0_12_sva_dfm_enexo_44 <= act_port_read_out_data_and_28_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_44 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_19_enex5 | act_regs_data_and_2748_enex5
        ) begin
      reg_act_port_read_out_data_0_3_sva_dfm_enexo_44 <= act_port_read_out_data_and_19_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_44 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_25_enex5 | act_regs_data_and_2748_enex5
        ) begin
      reg_act_port_read_out_data_0_9_sva_dfm_enexo_44 <= act_port_read_out_data_and_25_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_44 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_17_enex5 | act_regs_data_and_2748_enex5
        ) begin
      reg_act_port_read_out_data_0_1_sva_dfm_enexo_44 <= act_port_read_out_data_and_17_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_44 <= 1'b1;
    end
    else if ( ActUnit_PushOutput_if_for_i_and_tmp | act_regs_data_and_2748_enex5
        ) begin
      reg_ActUnit_PushOutput_if_for_i_4_0_sva_3_0_enexo_44 <= ActUnit_PushOutput_if_for_i_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_44 <= 1'b1;
    end
    else if ( ActUnit_RunLoad_if_a2_and_tmp | act_regs_data_and_2748_enex5 ) begin
      reg_nvhls_get_slc_2U_NVUINT8_return_3_enexo_44 <= ActUnit_RunLoad_if_a2_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_44 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_30_enex5 | act_regs_data_and_2748_enex5
        ) begin
      reg_act_port_read_out_data_0_14_sva_dfm_enexo_44 <= act_port_read_out_data_and_30_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_44 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_20_enex5 | act_regs_data_and_2748_enex5
        ) begin
      reg_act_port_read_out_data_0_4_sva_dfm_enexo_44 <= act_port_read_out_data_and_20_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_1_sva_dfm_2_21_0_enexo_1 <= 1'b1;
    end
    else if ( and_2033_cse | act_regs_data_and_2748_enex5 ) begin
      reg_act_regs_data_3_1_sva_dfm_2_21_0_enexo_1 <= and_2033_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_44 <= 1'b1;
    end
    else if ( act_port_read_out_data_and_18_enex5 | act_regs_data_and_2748_enex5
        ) begin
      reg_act_port_read_out_data_0_2_sva_dfm_enexo_44 <= act_port_read_out_data_and_18_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_174 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2749_enex5 ) begin
      reg_is_start_enexo_174 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_174 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2749_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_174 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_13_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_264_cse | act_regs_data_and_2749_enex5 ) begin
      reg_act_regs_data_0_13_sva_8_30_26_enexo_1 <= act_regs_data_and_264_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_1_30_26_enexo <=
          1'b1;
    end
    else if ( and_1927_tmp | act_regs_data_and_2749_enex5 ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_1_30_26_enexo <=
          and_1927_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_13_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2089_tmp | act_regs_data_and_2749_enex5 ) begin
      reg_act_regs_data_0_13_sva_dfm_2_30_26_enexo <= and_2089_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_174 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2749_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_174 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_175 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2750_enex5 ) begin
      reg_is_start_enexo_175 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_175 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2750_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_175 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_1_25_22_enexo <=
          1'b1;
    end
    else if ( and_1887_tmp | act_regs_data_and_2750_enex5 ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_1_25_22_enexo <=
          and_1887_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_13_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_264_cse | act_regs_data_and_2750_enex5 ) begin
      reg_act_regs_data_0_13_sva_8_25_22_enexo_1 <= act_regs_data_and_264_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_13_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_1961_cse | act_regs_data_and_2750_enex5 ) begin
      reg_act_regs_data_0_13_sva_dfm_2_25_22_enexo <= and_1961_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_175 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2750_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_175 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_176 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2751_enex5 ) begin
      reg_is_start_enexo_176 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_176 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2751_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_176 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_13_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_264_cse | act_regs_data_and_2751_enex5 ) begin
      reg_act_regs_data_0_13_sva_8_21_0_enexo_1 <= act_regs_data_and_264_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Silu_for_16_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo
          <= 1'b1;
    end
    else if ( and_2328_tmp | act_regs_data_and_2751_enex5 ) begin
      reg_Silu_for_16_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo
          <= and_2328_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_13_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_1961_cse | act_regs_data_and_2751_enex5 ) begin
      reg_act_regs_data_0_13_sva_dfm_2_21_0_enexo <= and_1961_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_176 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2751_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_176 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_177 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2752_enex5 ) begin
      reg_is_start_enexo_177 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_177 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2752_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_177 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_12_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_268_cse | act_regs_data_and_2752_enex5 ) begin
      reg_act_regs_data_0_12_sva_8_30_26_enexo_1 <= act_regs_data_and_268_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_1_30_26_enexo <=
          1'b1;
    end
    else if ( and_1921_tmp | act_regs_data_and_2752_enex5 ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_1_30_26_enexo <=
          and_1921_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_12_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2087_tmp | act_regs_data_and_2752_enex5 ) begin
      reg_act_regs_data_0_12_sva_dfm_2_30_26_enexo <= and_2087_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_177 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2752_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_177 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_178 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2753_enex5 ) begin
      reg_is_start_enexo_178 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_178 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2753_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_178 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_1_25_22_enexo <=
          1'b1;
    end
    else if ( and_1885_tmp | act_regs_data_and_2753_enex5 ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_1_25_22_enexo <=
          and_1885_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_12_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_268_cse | act_regs_data_and_2753_enex5 ) begin
      reg_act_regs_data_0_12_sva_8_25_22_enexo_1 <= act_regs_data_and_268_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_12_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_1959_cse | act_regs_data_and_2753_enex5 ) begin
      reg_act_regs_data_0_12_sva_dfm_2_25_22_enexo <= and_1959_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_178 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2753_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_178 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_179 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2754_enex5 ) begin
      reg_is_start_enexo_179 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_179 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2754_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_179 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_12_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_268_cse | act_regs_data_and_2754_enex5 ) begin
      reg_act_regs_data_0_12_sva_8_21_0_enexo_1 <= act_regs_data_and_268_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Silu_for_15_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo
          <= 1'b1;
    end
    else if ( and_2327_tmp | act_regs_data_and_2754_enex5 ) begin
      reg_Silu_for_15_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo
          <= and_2327_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_12_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_1959_cse | act_regs_data_and_2754_enex5 ) begin
      reg_act_regs_data_0_12_sva_dfm_2_21_0_enexo <= and_1959_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_179 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2754_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_179 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_180 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2755_enex5 ) begin
      reg_is_start_enexo_180 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_180 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2755_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_180 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_11_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_272_cse | act_regs_data_and_2755_enex5 ) begin
      reg_act_regs_data_0_11_sva_8_30_26_enexo_1 <= act_regs_data_and_272_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_1_30_26_enexo <=
          1'b1;
    end
    else if ( and_1915_tmp | act_regs_data_and_2755_enex5 ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_1_30_26_enexo <=
          and_1915_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_11_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2085_tmp | act_regs_data_and_2755_enex5 ) begin
      reg_act_regs_data_0_11_sva_dfm_2_30_26_enexo <= and_2085_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_180 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2755_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_180 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_181 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2756_enex5 ) begin
      reg_is_start_enexo_181 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_181 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2756_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_181 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_1_25_22_enexo <=
          1'b1;
    end
    else if ( and_1883_tmp | act_regs_data_and_2756_enex5 ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_1_25_22_enexo <=
          and_1883_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_11_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_272_cse | act_regs_data_and_2756_enex5 ) begin
      reg_act_regs_data_0_11_sva_8_25_22_enexo_1 <= act_regs_data_and_272_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_11_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_1957_cse | act_regs_data_and_2756_enex5 ) begin
      reg_act_regs_data_0_11_sva_dfm_2_25_22_enexo <= and_1957_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_181 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2756_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_181 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_182 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2757_enex5 ) begin
      reg_is_start_enexo_182 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_182 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2757_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_182 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_11_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_272_cse | act_regs_data_and_2757_enex5 ) begin
      reg_act_regs_data_0_11_sva_8_21_0_enexo_1 <= act_regs_data_and_272_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_11_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_1957_cse | act_regs_data_and_2757_enex5 ) begin
      reg_act_regs_data_0_11_sva_dfm_2_21_0_enexo <= and_1957_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_182 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2757_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_182 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Silu_for_14_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo
          <= 1'b1;
    end
    else if ( and_2326_tmp | act_regs_data_and_2757_enex5 ) begin
      reg_Silu_for_14_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo
          <= and_2326_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_183 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2758_enex5 ) begin
      reg_is_start_enexo_183 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_183 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2758_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_183 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_10_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_276_cse | act_regs_data_and_2758_enex5 ) begin
      reg_act_regs_data_0_10_sva_8_30_26_enexo_1 <= act_regs_data_and_276_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_1_30_26_enexo <=
          1'b1;
    end
    else if ( and_1909_tmp | act_regs_data_and_2758_enex5 ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_1_30_26_enexo <=
          and_1909_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_10_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2083_tmp | act_regs_data_and_2758_enex5 ) begin
      reg_act_regs_data_0_10_sva_dfm_2_30_26_enexo <= and_2083_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_183 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2758_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_183 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_184 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2759_enex5 ) begin
      reg_is_start_enexo_184 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_184 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2759_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_184 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_1_25_22_enexo <=
          1'b1;
    end
    else if ( and_1881_tmp | act_regs_data_and_2759_enex5 ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_1_25_22_enexo <=
          and_1881_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_10_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_276_cse | act_regs_data_and_2759_enex5 ) begin
      reg_act_regs_data_0_10_sva_8_25_22_enexo_1 <= act_regs_data_and_276_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_10_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_1955_cse | act_regs_data_and_2759_enex5 ) begin
      reg_act_regs_data_0_10_sva_dfm_2_25_22_enexo <= and_1955_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_184 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2759_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_184 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_185 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2760_enex5 ) begin
      reg_is_start_enexo_185 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_185 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2760_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_185 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_10_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_276_cse | act_regs_data_and_2760_enex5 ) begin
      reg_act_regs_data_0_10_sva_8_21_0_enexo_1 <= act_regs_data_and_276_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_10_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_1955_cse | act_regs_data_and_2760_enex5 ) begin
      reg_act_regs_data_0_10_sva_dfm_2_21_0_enexo <= and_1955_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_185 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2760_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_185 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Silu_for_13_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo
          <= 1'b1;
    end
    else if ( and_2325_tmp | act_regs_data_and_2760_enex5 ) begin
      reg_Silu_for_13_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo
          <= and_2325_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_186 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2761_enex5 ) begin
      reg_is_start_enexo_186 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_1_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_312_cse | act_regs_data_and_2761_enex5 ) begin
      reg_act_regs_data_0_1_sva_8_30_26_enexo_1 <= act_regs_data_and_312_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_186 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2761_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_186 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_71_64_sva_dfm_6_1_enexo <= 1'b1;
    end
    else if ( and_1803_tmp | act_regs_data_and_2761_enex5 ) begin
      reg_rva_out_reg_data_71_64_sva_dfm_6_1_enexo <= and_1803_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_1_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2065_tmp | act_regs_data_and_2761_enex5 ) begin
      reg_act_regs_data_0_1_sva_dfm_2_30_26_enexo <= and_2065_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_186 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2761_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_186 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_187 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2762_enex5 ) begin
      reg_is_start_enexo_187 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_1_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_312_cse | act_regs_data_and_2762_enex5 ) begin
      reg_act_regs_data_0_1_sva_8_25_22_enexo_1 <= act_regs_data_and_312_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_187 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2762_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_187 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_39_32_sva_dfm_6_1_enexo <= 1'b1;
    end
    else if ( and_1801_tmp | act_regs_data_and_2762_enex5 ) begin
      reg_rva_out_reg_data_39_32_sva_dfm_6_1_enexo <= and_1801_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_1_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_1937_cse | act_regs_data_and_2762_enex5 ) begin
      reg_act_regs_data_0_1_sva_dfm_2_25_22_enexo <= and_1937_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_187 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2762_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_187 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_188 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2763_enex5 ) begin
      reg_is_start_enexo_188 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_1_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_312_cse | act_regs_data_and_2763_enex5 ) begin
      reg_act_regs_data_0_1_sva_8_21_0_enexo_1 <= act_regs_data_and_312_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_188 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2763_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_188 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_1_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_1937_cse | act_regs_data_and_2763_enex5 ) begin
      reg_act_regs_data_0_1_sva_dfm_2_21_0_enexo <= and_1937_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_188 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2763_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_188 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Silu_for_12_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo
          <= 1'b1;
    end
    else if ( and_2324_tmp | act_regs_data_and_2763_enex5 ) begin
      reg_Silu_for_12_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo
          <= and_2324_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_1_30_26_enexo <=
          1'b1;
    end
    else if ( and_1808_tmp | act_regs_data_and_2764_enex5 ) begin
      reg_ActUnit_PushOutput_if_output_port_reg_data_data_0_sva_1_30_26_enexo <=
          and_1808_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_189 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2764_enex5 ) begin
      reg_is_start_enexo_189 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_189 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2764_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_189 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_0_sva_8_30_26_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_316_cse | act_regs_data_and_2764_enex5 ) begin
      reg_act_regs_data_0_0_sva_8_30_26_enexo_1 <= act_regs_data_and_316_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_0_sva_dfm_2_30_26_enexo <= 1'b1;
    end
    else if ( and_2063_tmp | act_regs_data_and_2764_enex5 ) begin
      reg_act_regs_data_0_0_sva_dfm_2_30_26_enexo <= and_2063_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_189 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2764_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_189 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_190 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2765_enex5 ) begin
      reg_is_start_enexo_190 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_190 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2765_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_190 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_rva_out_reg_data_29_24_sva_dfm_6_1_enexo <= 1'b1;
    end
    else if ( rva_out_reg_data_and_61_tmp | act_regs_data_and_2765_enex5 ) begin
      reg_rva_out_reg_data_29_24_sva_dfm_6_1_enexo <= rva_out_reg_data_and_61_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_0_sva_8_25_22_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_316_cse | act_regs_data_and_2765_enex5 ) begin
      reg_act_regs_data_0_0_sva_8_25_22_enexo_1 <= act_regs_data_and_316_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_0_sva_dfm_2_25_22_enexo <= 1'b1;
    end
    else if ( and_1935_cse | act_regs_data_and_2765_enex5 ) begin
      reg_act_regs_data_0_0_sva_dfm_2_25_22_enexo <= and_1935_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_190 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2765_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_190 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_is_start_enexo_191 <= 1'b1;
    end
    else if ( is_start_and_tmp | act_regs_data_and_2766_enex5 ) begin
      reg_is_start_enexo_191 <= is_start_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_191 <= 1'b1;
    end
    else if ( act_config_output_counter_and_1_cse | act_regs_data_and_2766_enex5
        ) begin
      reg_act_config_is_zero_first_sva_dfm_4_enexo_191 <= act_config_output_counter_and_1_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_0_sva_8_21_0_enexo_1 <= 1'b1;
    end
    else if ( act_regs_data_and_316_cse | act_regs_data_and_2766_enex5 ) begin
      reg_act_regs_data_0_0_sva_8_21_0_enexo_1 <= act_regs_data_and_316_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_0_sva_dfm_2_21_0_enexo <= 1'b1;
    end
    else if ( and_1935_cse | act_regs_data_and_2766_enex5 ) begin
      reg_act_regs_data_0_0_sva_dfm_2_21_0_enexo <= and_1935_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_Silu_for_11_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo
          <= 1'b1;
    end
    else if ( Silu_for_else_else_else_if_and_tmp | act_regs_data_and_2766_enex5 )
        begin
      reg_Silu_for_11_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_1_enexo
          <= Silu_for_else_else_else_if_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_w_load_lpi_1_dfm_1_enexo_191 <= 1'b1;
    end
    else if ( w_load_and_tmp | act_regs_data_and_2766_enex5 ) begin
      reg_w_load_lpi_1_dfm_1_enexo_191 <= w_load_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_177 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | ActUnit_RunInst_switch_lp_and_816_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_177 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_177 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | ActUnit_RunInst_switch_lp_and_816_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_177 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_177 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | ActUnit_RunInst_switch_lp_and_816_enex5
        ) begin
      reg_act_config_inst_counter_enexo_177 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_0_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2576_enex5 | ActUnit_RunInst_switch_lp_and_816_enex5
        ) begin
      reg_act_regs_data_3_0_2_enexo_5 <= act_regs_data_and_2576_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_0_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2765_enex5 | ActUnit_RunInst_switch_lp_and_816_enex5
        ) begin
      reg_act_regs_data_0_0_2_enexo_5 <= act_regs_data_and_2765_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_0_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2672_enex5 | ActUnit_RunInst_switch_lp_and_816_enex5
        ) begin
      reg_act_regs_data_1_0_2_enexo_5 <= act_regs_data_and_2672_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_0_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2624_enex5 | ActUnit_RunInst_switch_lp_and_816_enex5
        ) begin
      reg_act_regs_data_2_0_2_enexo_5 <= act_regs_data_and_2624_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_178 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | ActUnit_RunInst_switch_lp_and_817_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_178 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_178 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | ActUnit_RunInst_switch_lp_and_817_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_178 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_178 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | ActUnit_RunInst_switch_lp_and_817_enex5
        ) begin
      reg_act_config_inst_counter_enexo_178 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_0_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2577_enex5 | ActUnit_RunInst_switch_lp_and_817_enex5
        ) begin
      reg_act_regs_data_3_0_3_enexo_5 <= act_regs_data_and_2577_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_0_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2766_enex5 | ActUnit_RunInst_switch_lp_and_817_enex5
        ) begin
      reg_act_regs_data_0_0_3_enexo_5 <= act_regs_data_and_2766_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_0_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2625_enex5 | ActUnit_RunInst_switch_lp_and_817_enex5
        ) begin
      reg_act_regs_data_2_0_3_enexo_5 <= act_regs_data_and_2625_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_0_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2673_enex5 | ActUnit_RunInst_switch_lp_and_817_enex5
        ) begin
      reg_act_regs_data_1_0_3_enexo_5 <= act_regs_data_and_2673_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_179 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | ActUnit_RunInst_switch_lp_and_818_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_179 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_0_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2575_enex5 | ActUnit_RunInst_switch_lp_and_818_enex5
        ) begin
      reg_act_regs_data_3_0_1_enexo_5 <= act_regs_data_and_2575_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_179 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | ActUnit_RunInst_switch_lp_and_818_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_179 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_179 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | ActUnit_RunInst_switch_lp_and_818_enex5
        ) begin
      reg_act_config_inst_counter_enexo_179 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_0_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2764_enex5 | ActUnit_RunInst_switch_lp_and_818_enex5
        ) begin
      reg_act_regs_data_0_0_1_enexo_5 <= act_regs_data_and_2764_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_0_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2623_enex5 | ActUnit_RunInst_switch_lp_and_818_enex5
        ) begin
      reg_act_regs_data_2_0_1_enexo_5 <= act_regs_data_and_2623_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_0_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2671_enex5 | ActUnit_RunInst_switch_lp_and_818_enex5
        ) begin
      reg_act_regs_data_1_0_1_enexo_5 <= act_regs_data_and_2671_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_180 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_180 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_180 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_180 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_180 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_enex5
        ) begin
      reg_act_config_inst_counter_enexo_180 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_1_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2669_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_enex5
        ) begin
      reg_act_regs_data_1_1_2_enexo_5 <= act_regs_data_and_2669_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_1_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2573_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_enex5
        ) begin
      reg_act_regs_data_3_1_2_enexo_5 <= act_regs_data_and_2573_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_1_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2762_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_enex5
        ) begin
      reg_act_regs_data_0_1_2_enexo_5 <= act_regs_data_and_2762_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_1_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2621_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_enex5
        ) begin
      reg_act_regs_data_2_1_2_enexo_5 <= act_regs_data_and_2621_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_181 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_15_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_181 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_181 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_15_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_181 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_181 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_15_enex5
        ) begin
      reg_act_config_inst_counter_enexo_181 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_1_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2763_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_15_enex5
        ) begin
      reg_act_regs_data_0_1_3_enexo_5 <= act_regs_data_and_2763_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_1_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2574_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_15_enex5
        ) begin
      reg_act_regs_data_3_1_3_enexo_5 <= act_regs_data_and_2574_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_1_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2670_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_15_enex5
        ) begin
      reg_act_regs_data_1_1_3_enexo_5 <= act_regs_data_and_2670_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_1_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2622_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_15_enex5
        ) begin
      reg_act_regs_data_2_1_3_enexo_5 <= act_regs_data_and_2622_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_182 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_16_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_182 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_182 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_16_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_182 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_1_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2620_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_16_enex5
        ) begin
      reg_act_regs_data_2_1_1_enexo_5 <= act_regs_data_and_2620_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_182 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_16_enex5
        ) begin
      reg_act_config_inst_counter_enexo_182 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_1_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2572_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_16_enex5
        ) begin
      reg_act_regs_data_3_1_1_enexo_5 <= act_regs_data_and_2572_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_1_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2761_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_16_enex5
        ) begin
      reg_act_regs_data_0_1_1_enexo_5 <= act_regs_data_and_2761_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_1_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2668_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_16_enex5
        ) begin
      reg_act_regs_data_1_1_1_enexo_5 <= act_regs_data_and_2668_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_183 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_17_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_183 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_183 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_17_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_183 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_183 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_17_enex5
        ) begin
      reg_act_config_inst_counter_enexo_183 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_2_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2702_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_17_enex5
        ) begin
      reg_act_regs_data_0_2_2_enexo_5 <= act_regs_data_and_2702_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_2_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2666_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_17_enex5
        ) begin
      reg_act_regs_data_1_2_2_enexo_5 <= act_regs_data_and_2666_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_2_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2570_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_17_enex5
        ) begin
      reg_act_regs_data_3_2_2_enexo_5 <= act_regs_data_and_2570_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_2_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2618_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_17_enex5
        ) begin
      reg_act_regs_data_2_2_2_enexo_5 <= act_regs_data_and_2618_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_184 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_18_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_184 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_184 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_18_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_184 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_184 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_18_enex5
        ) begin
      reg_act_config_inst_counter_enexo_184 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_2_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2571_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_18_enex5
        ) begin
      reg_act_regs_data_3_2_3_enexo_5 <= act_regs_data_and_2571_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_2_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2619_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_18_enex5
        ) begin
      reg_act_regs_data_2_2_3_enexo_5 <= act_regs_data_and_2619_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_2_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2703_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_18_enex5
        ) begin
      reg_act_regs_data_0_2_3_enexo_5 <= act_regs_data_and_2703_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_2_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2667_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_18_enex5
        ) begin
      reg_act_regs_data_1_2_3_enexo_5 <= act_regs_data_and_2667_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_2_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2617_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_19_enex5
        ) begin
      reg_act_regs_data_2_2_1_enexo_5 <= act_regs_data_and_2617_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_185 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_19_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_185 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_185 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_19_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_185 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_185 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_19_enex5
        ) begin
      reg_act_config_inst_counter_enexo_185 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_2_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2569_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_19_enex5
        ) begin
      reg_act_regs_data_3_2_1_enexo_5 <= act_regs_data_and_2569_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_2_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2665_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_19_enex5
        ) begin
      reg_act_regs_data_1_2_1_enexo_5 <= act_regs_data_and_2665_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_2_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2701_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_19_enex5
        ) begin
      reg_act_regs_data_0_2_1_enexo_5 <= act_regs_data_and_2701_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_186 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_20_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_186 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_186 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_20_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_186 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_186 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_20_enex5
        ) begin
      reg_act_config_inst_counter_enexo_186 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_3_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2699_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_20_enex5
        ) begin
      reg_act_regs_data_0_3_2_enexo_5 <= act_regs_data_and_2699_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_3_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2663_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_20_enex5
        ) begin
      reg_act_regs_data_1_3_2_enexo_5 <= act_regs_data_and_2663_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_3_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2567_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_20_enex5
        ) begin
      reg_act_regs_data_3_3_2_enexo_5 <= act_regs_data_and_2567_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_3_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2615_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_20_enex5
        ) begin
      reg_act_regs_data_2_3_2_enexo_5 <= act_regs_data_and_2615_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_187 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_21_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_187 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_187 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_21_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_187 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_187 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_21_enex5
        ) begin
      reg_act_config_inst_counter_enexo_187 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_3_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2700_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_21_enex5
        ) begin
      reg_act_regs_data_0_3_3_enexo_5 <= act_regs_data_and_2700_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_3_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2568_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_21_enex5
        ) begin
      reg_act_regs_data_3_3_3_enexo_5 <= act_regs_data_and_2568_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_3_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2664_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_21_enex5
        ) begin
      reg_act_regs_data_1_3_3_enexo_5 <= act_regs_data_and_2664_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_3_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2616_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_21_enex5
        ) begin
      reg_act_regs_data_2_3_3_enexo_5 <= act_regs_data_and_2616_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_188 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_22_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_188 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_188 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_22_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_188 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_188 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_22_enex5
        ) begin
      reg_act_config_inst_counter_enexo_188 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_3_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2698_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_22_enex5
        ) begin
      reg_act_regs_data_0_3_1_enexo_5 <= act_regs_data_and_2698_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_3_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2566_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_22_enex5
        ) begin
      reg_act_regs_data_3_3_1_enexo_5 <= act_regs_data_and_2566_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_3_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2662_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_22_enex5
        ) begin
      reg_act_regs_data_1_3_1_enexo_5 <= act_regs_data_and_2662_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_3_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2614_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_22_enex5
        ) begin
      reg_act_regs_data_2_3_1_enexo_5 <= act_regs_data_and_2614_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_189 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_23_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_189 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_189 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_23_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_189 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_189 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_23_enex5
        ) begin
      reg_act_config_inst_counter_enexo_189 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_4_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2564_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_23_enex5
        ) begin
      reg_act_regs_data_3_4_2_enexo_5 <= act_regs_data_and_2564_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_4_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2660_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_23_enex5
        ) begin
      reg_act_regs_data_1_4_2_enexo_5 <= act_regs_data_and_2660_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_4_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2696_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_23_enex5
        ) begin
      reg_act_regs_data_0_4_2_enexo_5 <= act_regs_data_and_2696_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_4_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2612_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_23_enex5
        ) begin
      reg_act_regs_data_2_4_2_enexo_5 <= act_regs_data_and_2612_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_190 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_24_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_190 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_190 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_24_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_190 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_190 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_24_enex5
        ) begin
      reg_act_config_inst_counter_enexo_190 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_4_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2697_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_24_enex5
        ) begin
      reg_act_regs_data_0_4_3_enexo_5 <= act_regs_data_and_2697_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_4_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2661_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_24_enex5
        ) begin
      reg_act_regs_data_1_4_3_enexo_5 <= act_regs_data_and_2661_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_4_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2565_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_24_enex5
        ) begin
      reg_act_regs_data_3_4_3_enexo_5 <= act_regs_data_and_2565_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_4_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2613_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_24_enex5
        ) begin
      reg_act_regs_data_2_4_3_enexo_5 <= act_regs_data_and_2613_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_191 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_25_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_191 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_191 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_25_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_191 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_191 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_25_enex5
        ) begin
      reg_act_config_inst_counter_enexo_191 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_4_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2563_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_25_enex5
        ) begin
      reg_act_regs_data_3_4_1_enexo_5 <= act_regs_data_and_2563_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_4_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2695_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_25_enex5
        ) begin
      reg_act_regs_data_0_4_1_enexo_5 <= act_regs_data_and_2695_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_4_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2611_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_25_enex5
        ) begin
      reg_act_regs_data_2_4_1_enexo_5 <= act_regs_data_and_2611_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_4_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2659_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_25_enex5
        ) begin
      reg_act_regs_data_1_4_1_enexo_5 <= act_regs_data_and_2659_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_192 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_26_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_192 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_192 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_26_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_192 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_192 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_26_enex5
        ) begin
      reg_act_config_inst_counter_enexo_192 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_5_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2609_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_26_enex5
        ) begin
      reg_act_regs_data_2_5_2_enexo_5 <= act_regs_data_and_2609_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_5_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2657_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_26_enex5
        ) begin
      reg_act_regs_data_1_5_2_enexo_5 <= act_regs_data_and_2657_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_5_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2561_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_26_enex5
        ) begin
      reg_act_regs_data_3_5_2_enexo_5 <= act_regs_data_and_2561_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_5_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2693_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_26_enex5
        ) begin
      reg_act_regs_data_0_5_2_enexo_5 <= act_regs_data_and_2693_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_193 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_27_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_193 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_193 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_27_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_193 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_5_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2694_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_27_enex5
        ) begin
      reg_act_regs_data_0_5_3_enexo_5 <= act_regs_data_and_2694_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_193 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_27_enex5
        ) begin
      reg_act_config_inst_counter_enexo_193 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_5_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2658_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_27_enex5
        ) begin
      reg_act_regs_data_1_5_3_enexo_5 <= act_regs_data_and_2658_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_5_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2562_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_27_enex5
        ) begin
      reg_act_regs_data_3_5_3_enexo_5 <= act_regs_data_and_2562_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_5_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2610_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_27_enex5
        ) begin
      reg_act_regs_data_2_5_3_enexo_5 <= act_regs_data_and_2610_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_194 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_28_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_194 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_194 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_28_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_194 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_194 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_28_enex5
        ) begin
      reg_act_config_inst_counter_enexo_194 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_5_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2560_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_28_enex5
        ) begin
      reg_act_regs_data_3_5_1_enexo_5 <= act_regs_data_and_2560_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_5_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2692_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_28_enex5
        ) begin
      reg_act_regs_data_0_5_1_enexo_5 <= act_regs_data_and_2692_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_5_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2656_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_28_enex5
        ) begin
      reg_act_regs_data_1_5_1_enexo_5 <= act_regs_data_and_2656_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_5_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2608_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_28_enex5
        ) begin
      reg_act_regs_data_2_5_1_enexo_5 <= act_regs_data_and_2608_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_195 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_29_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_195 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_195 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_29_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_195 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_195 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_29_enex5
        ) begin
      reg_act_config_inst_counter_enexo_195 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_6_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2606_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_29_enex5
        ) begin
      reg_act_regs_data_2_6_2_enexo_5 <= act_regs_data_and_2606_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_6_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2654_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_29_enex5
        ) begin
      reg_act_regs_data_1_6_2_enexo_5 <= act_regs_data_and_2654_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_6_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2558_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_29_enex5
        ) begin
      reg_act_regs_data_3_6_2_enexo_5 <= act_regs_data_and_2558_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_6_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2690_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_29_enex5
        ) begin
      reg_act_regs_data_0_6_2_enexo_5 <= act_regs_data_and_2690_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_196 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_30_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_196 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_196 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_30_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_196 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_196 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_30_enex5
        ) begin
      reg_act_config_inst_counter_enexo_196 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_6_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2607_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_30_enex5
        ) begin
      reg_act_regs_data_2_6_3_enexo_5 <= act_regs_data_and_2607_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_6_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2559_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_30_enex5
        ) begin
      reg_act_regs_data_3_6_3_enexo_5 <= act_regs_data_and_2559_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_6_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2691_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_30_enex5
        ) begin
      reg_act_regs_data_0_6_3_enexo_5 <= act_regs_data_and_2691_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_6_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2655_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_30_enex5
        ) begin
      reg_act_regs_data_1_6_3_enexo_5 <= act_regs_data_and_2655_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_197 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_31_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_197 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_197 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_31_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_197 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_197 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_31_enex5
        ) begin
      reg_act_config_inst_counter_enexo_197 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_6_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2557_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_31_enex5
        ) begin
      reg_act_regs_data_3_6_1_enexo_5 <= act_regs_data_and_2557_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_6_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2653_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_31_enex5
        ) begin
      reg_act_regs_data_1_6_1_enexo_5 <= act_regs_data_and_2653_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_6_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2605_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_31_enex5
        ) begin
      reg_act_regs_data_2_6_1_enexo_5 <= act_regs_data_and_2605_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_6_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2689_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_31_enex5
        ) begin
      reg_act_regs_data_0_6_1_enexo_5 <= act_regs_data_and_2689_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_198 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_32_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_198 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_198 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_32_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_198 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_198 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_32_enex5
        ) begin
      reg_act_config_inst_counter_enexo_198 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_7_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2687_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_32_enex5
        ) begin
      reg_act_regs_data_0_7_2_enexo_5 <= act_regs_data_and_2687_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_7_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2603_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_32_enex5
        ) begin
      reg_act_regs_data_2_7_2_enexo_5 <= act_regs_data_and_2603_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_7_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2555_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_32_enex5
        ) begin
      reg_act_regs_data_3_7_2_enexo_5 <= act_regs_data_and_2555_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_7_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2651_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_32_enex5
        ) begin
      reg_act_regs_data_1_7_2_enexo_5 <= act_regs_data_and_2651_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_199 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_33_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_199 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_199 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_33_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_199 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_199 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_33_enex5
        ) begin
      reg_act_config_inst_counter_enexo_199 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_7_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2688_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_33_enex5
        ) begin
      reg_act_regs_data_0_7_3_enexo_5 <= act_regs_data_and_2688_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_7_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2652_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_33_enex5
        ) begin
      reg_act_regs_data_1_7_3_enexo_5 <= act_regs_data_and_2652_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_7_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2556_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_33_enex5
        ) begin
      reg_act_regs_data_3_7_3_enexo_5 <= act_regs_data_and_2556_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_7_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2604_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_33_enex5
        ) begin
      reg_act_regs_data_2_7_3_enexo_5 <= act_regs_data_and_2604_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_200 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_34_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_200 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_200 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_34_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_200 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_200 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_34_enex5
        ) begin
      reg_act_config_inst_counter_enexo_200 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_7_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2554_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_34_enex5
        ) begin
      reg_act_regs_data_3_7_1_enexo_5 <= act_regs_data_and_2554_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_7_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2650_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_34_enex5
        ) begin
      reg_act_regs_data_1_7_1_enexo_5 <= act_regs_data_and_2650_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_7_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2686_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_34_enex5
        ) begin
      reg_act_regs_data_0_7_1_enexo_5 <= act_regs_data_and_2686_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_7_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2602_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_34_enex5
        ) begin
      reg_act_regs_data_2_7_1_enexo_5 <= act_regs_data_and_2602_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_201 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_35_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_201 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_201 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_35_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_201 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_201 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_35_enex5
        ) begin
      reg_act_config_inst_counter_enexo_201 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_8_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2684_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_35_enex5
        ) begin
      reg_act_regs_data_0_8_2_enexo_5 <= act_regs_data_and_2684_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_8_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2648_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_35_enex5
        ) begin
      reg_act_regs_data_1_8_2_enexo_5 <= act_regs_data_and_2648_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_8_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2600_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_35_enex5
        ) begin
      reg_act_regs_data_2_8_2_enexo_5 <= act_regs_data_and_2600_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_8_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2552_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_35_enex5
        ) begin
      reg_act_regs_data_3_8_2_enexo_5 <= act_regs_data_and_2552_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_202 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_36_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_202 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_202 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_36_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_202 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_202 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_36_enex5
        ) begin
      reg_act_config_inst_counter_enexo_202 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_8_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2685_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_36_enex5
        ) begin
      reg_act_regs_data_0_8_3_enexo_5 <= act_regs_data_and_2685_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_8_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2601_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_36_enex5
        ) begin
      reg_act_regs_data_2_8_3_enexo_5 <= act_regs_data_and_2601_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_8_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2649_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_36_enex5
        ) begin
      reg_act_regs_data_1_8_3_enexo_5 <= act_regs_data_and_2649_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_8_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2553_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_36_enex5
        ) begin
      reg_act_regs_data_3_8_3_enexo_5 <= act_regs_data_and_2553_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_203 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_37_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_203 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_203 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_37_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_203 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_203 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_37_enex5
        ) begin
      reg_act_config_inst_counter_enexo_203 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_8_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2599_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_37_enex5
        ) begin
      reg_act_regs_data_2_8_1_enexo_5 <= act_regs_data_and_2599_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_8_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2683_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_37_enex5
        ) begin
      reg_act_regs_data_0_8_1_enexo_5 <= act_regs_data_and_2683_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_8_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2551_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_37_enex5
        ) begin
      reg_act_regs_data_3_8_1_enexo_5 <= act_regs_data_and_2551_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_8_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2647_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_37_enex5
        ) begin
      reg_act_regs_data_1_8_1_enexo_5 <= act_regs_data_and_2647_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_204 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_38_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_204 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_204 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_38_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_204 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_204 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_38_enex5
        ) begin
      reg_act_config_inst_counter_enexo_204 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_9_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2681_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_38_enex5
        ) begin
      reg_act_regs_data_0_9_2_enexo_5 <= act_regs_data_and_2681_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_9_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2597_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_38_enex5
        ) begin
      reg_act_regs_data_2_9_2_enexo_5 <= act_regs_data_and_2597_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_9_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2645_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_38_enex5
        ) begin
      reg_act_regs_data_1_9_2_enexo_5 <= act_regs_data_and_2645_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_9_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2549_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_38_enex5
        ) begin
      reg_act_regs_data_3_9_2_enexo_5 <= act_regs_data_and_2549_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_205 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_39_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_205 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_205 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_39_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_205 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_205 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_39_enex5
        ) begin
      reg_act_config_inst_counter_enexo_205 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_9_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2646_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_39_enex5
        ) begin
      reg_act_regs_data_1_9_3_enexo_5 <= act_regs_data_and_2646_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_9_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2682_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_39_enex5
        ) begin
      reg_act_regs_data_0_9_3_enexo_5 <= act_regs_data_and_2682_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_9_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2598_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_39_enex5
        ) begin
      reg_act_regs_data_2_9_3_enexo_5 <= act_regs_data_and_2598_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_9_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2550_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_39_enex5
        ) begin
      reg_act_regs_data_3_9_3_enexo_5 <= act_regs_data_and_2550_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_206 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_40_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_206 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_206 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_40_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_206 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_206 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_40_enex5
        ) begin
      reg_act_config_inst_counter_enexo_206 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_9_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2644_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_40_enex5
        ) begin
      reg_act_regs_data_1_9_1_enexo_5 <= act_regs_data_and_2644_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_9_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2548_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_40_enex5
        ) begin
      reg_act_regs_data_3_9_1_enexo_5 <= act_regs_data_and_2548_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_9_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2680_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_40_enex5
        ) begin
      reg_act_regs_data_0_9_1_enexo_5 <= act_regs_data_and_2680_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_9_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2596_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_40_enex5
        ) begin
      reg_act_regs_data_2_9_1_enexo_5 <= act_regs_data_and_2596_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_207 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_41_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_207 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_207 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_41_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_207 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_207 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_41_enex5
        ) begin
      reg_act_config_inst_counter_enexo_207 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_10_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2642_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_41_enex5
        ) begin
      reg_act_regs_data_1_10_2_enexo_5 <= act_regs_data_and_2642_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_10_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2759_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_41_enex5
        ) begin
      reg_act_regs_data_0_10_2_enexo_5 <= act_regs_data_and_2759_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_10_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2546_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_41_enex5
        ) begin
      reg_act_regs_data_3_10_2_enexo_5 <= act_regs_data_and_2546_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_10_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2594_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_41_enex5
        ) begin
      reg_act_regs_data_2_10_2_enexo_5 <= act_regs_data_and_2594_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_208 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_42_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_208 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_208 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_42_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_208 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_208 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_42_enex5
        ) begin
      reg_act_config_inst_counter_enexo_208 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_10_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2547_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_42_enex5
        ) begin
      reg_act_regs_data_3_10_3_enexo_5 <= act_regs_data_and_2547_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_10_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2760_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_42_enex5
        ) begin
      reg_act_regs_data_0_10_3_enexo_5 <= act_regs_data_and_2760_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_10_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2595_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_42_enex5
        ) begin
      reg_act_regs_data_2_10_3_enexo_5 <= act_regs_data_and_2595_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_10_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2643_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_42_enex5
        ) begin
      reg_act_regs_data_1_10_3_enexo_5 <= act_regs_data_and_2643_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_209 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_43_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_209 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_209 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_43_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_209 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_209 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_43_enex5
        ) begin
      reg_act_config_inst_counter_enexo_209 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_10_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2641_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_43_enex5
        ) begin
      reg_act_regs_data_1_10_1_enexo_5 <= act_regs_data_and_2641_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_10_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2593_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_43_enex5
        ) begin
      reg_act_regs_data_2_10_1_enexo_5 <= act_regs_data_and_2593_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_10_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2545_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_43_enex5
        ) begin
      reg_act_regs_data_3_10_1_enexo_5 <= act_regs_data_and_2545_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_10_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2758_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_43_enex5
        ) begin
      reg_act_regs_data_0_10_1_enexo_5 <= act_regs_data_and_2758_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_210 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_44_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_210 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_210 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_44_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_210 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_210 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_44_enex5
        ) begin
      reg_act_config_inst_counter_enexo_210 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_11_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2591_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_44_enex5
        ) begin
      reg_act_regs_data_2_11_2_enexo_5 <= act_regs_data_and_2591_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_11_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2756_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_44_enex5
        ) begin
      reg_act_regs_data_0_11_2_enexo_5 <= act_regs_data_and_2756_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_11_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2543_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_44_enex5
        ) begin
      reg_act_regs_data_3_11_2_enexo_5 <= act_regs_data_and_2543_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_11_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2639_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_44_enex5
        ) begin
      reg_act_regs_data_1_11_2_enexo_5 <= act_regs_data_and_2639_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_211 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_45_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_211 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_211 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_45_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_211 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_211 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_45_enex5
        ) begin
      reg_act_config_inst_counter_enexo_211 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_11_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2757_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_45_enex5
        ) begin
      reg_act_regs_data_0_11_3_enexo_5 <= act_regs_data_and_2757_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_11_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2640_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_45_enex5
        ) begin
      reg_act_regs_data_1_11_3_enexo_5 <= act_regs_data_and_2640_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_11_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2592_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_45_enex5
        ) begin
      reg_act_regs_data_2_11_3_enexo_5 <= act_regs_data_and_2592_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_11_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2544_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_45_enex5
        ) begin
      reg_act_regs_data_3_11_3_enexo_5 <= act_regs_data_and_2544_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_212 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_46_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_212 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_212 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_46_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_212 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_212 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_46_enex5
        ) begin
      reg_act_config_inst_counter_enexo_212 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_11_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2590_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_46_enex5
        ) begin
      reg_act_regs_data_2_11_1_enexo_5 <= act_regs_data_and_2590_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_11_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2542_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_46_enex5
        ) begin
      reg_act_regs_data_3_11_1_enexo_5 <= act_regs_data_and_2542_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_11_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2755_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_46_enex5
        ) begin
      reg_act_regs_data_0_11_1_enexo_5 <= act_regs_data_and_2755_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_11_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2638_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_46_enex5
        ) begin
      reg_act_regs_data_1_11_1_enexo_5 <= act_regs_data_and_2638_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_213 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_47_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_213 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_213 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_47_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_213 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_12_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2588_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_47_enex5
        ) begin
      reg_act_regs_data_2_12_2_enexo_5 <= act_regs_data_and_2588_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_213 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_47_enex5
        ) begin
      reg_act_config_inst_counter_enexo_213 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_12_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2753_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_47_enex5
        ) begin
      reg_act_regs_data_0_12_2_enexo_5 <= act_regs_data_and_2753_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_12_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2540_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_47_enex5
        ) begin
      reg_act_regs_data_3_12_2_enexo_5 <= act_regs_data_and_2540_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_12_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2636_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_47_enex5
        ) begin
      reg_act_regs_data_1_12_2_enexo_5 <= act_regs_data_and_2636_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_214 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_48_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_214 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_214 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_48_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_214 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_214 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_48_enex5
        ) begin
      reg_act_config_inst_counter_enexo_214 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_12_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2754_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_48_enex5
        ) begin
      reg_act_regs_data_0_12_3_enexo_5 <= act_regs_data_and_2754_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_12_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2589_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_48_enex5
        ) begin
      reg_act_regs_data_2_12_3_enexo_5 <= act_regs_data_and_2589_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_12_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2541_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_48_enex5
        ) begin
      reg_act_regs_data_3_12_3_enexo_5 <= act_regs_data_and_2541_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_12_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2637_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_48_enex5
        ) begin
      reg_act_regs_data_1_12_3_enexo_5 <= act_regs_data_and_2637_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_215 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_49_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_215 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_215 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_49_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_215 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_215 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_49_enex5
        ) begin
      reg_act_config_inst_counter_enexo_215 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_12_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2587_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_49_enex5
        ) begin
      reg_act_regs_data_2_12_1_enexo_5 <= act_regs_data_and_2587_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_12_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2752_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_49_enex5
        ) begin
      reg_act_regs_data_0_12_1_enexo_5 <= act_regs_data_and_2752_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_12_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2635_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_49_enex5
        ) begin
      reg_act_regs_data_1_12_1_enexo_5 <= act_regs_data_and_2635_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_12_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2539_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_49_enex5
        ) begin
      reg_act_regs_data_3_12_1_enexo_5 <= act_regs_data_and_2539_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_13_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2537_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_50_enex5
        ) begin
      reg_act_regs_data_3_13_2_enexo_5 <= act_regs_data_and_2537_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_216 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_50_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_216 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_216 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_50_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_216 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_13_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2750_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_50_enex5
        ) begin
      reg_act_regs_data_0_13_2_enexo_5 <= act_regs_data_and_2750_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_216 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_50_enex5
        ) begin
      reg_act_config_inst_counter_enexo_216 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_13_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2633_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_50_enex5
        ) begin
      reg_act_regs_data_1_13_2_enexo_5 <= act_regs_data_and_2633_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_13_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2585_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_50_enex5
        ) begin
      reg_act_regs_data_2_13_2_enexo_5 <= act_regs_data_and_2585_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_217 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_51_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_217 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_217 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_51_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_217 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_217 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_51_enex5
        ) begin
      reg_act_config_inst_counter_enexo_217 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_13_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2586_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_51_enex5
        ) begin
      reg_act_regs_data_2_13_3_enexo_5 <= act_regs_data_and_2586_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_13_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2538_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_51_enex5
        ) begin
      reg_act_regs_data_3_13_3_enexo_5 <= act_regs_data_and_2538_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_13_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2634_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_51_enex5
        ) begin
      reg_act_regs_data_1_13_3_enexo_5 <= act_regs_data_and_2634_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_13_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2751_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_51_enex5
        ) begin
      reg_act_regs_data_0_13_3_enexo_5 <= act_regs_data_and_2751_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_218 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_52_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_218 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_13_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2632_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_52_enex5
        ) begin
      reg_act_regs_data_1_13_1_enexo_5 <= act_regs_data_and_2632_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_13_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2584_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_52_enex5
        ) begin
      reg_act_regs_data_2_13_1_enexo_5 <= act_regs_data_and_2584_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_218 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_52_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_218 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_218 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_52_enex5
        ) begin
      reg_act_config_inst_counter_enexo_218 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_13_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2749_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_52_enex5
        ) begin
      reg_act_regs_data_0_13_1_enexo_5 <= act_regs_data_and_2749_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_13_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2536_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_52_enex5
        ) begin
      reg_act_regs_data_3_13_1_enexo_5 <= act_regs_data_and_2536_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_219 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_53_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_219 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_14_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2678_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_53_enex5
        ) begin
      reg_act_regs_data_0_14_2_enexo_5 <= act_regs_data_and_2678_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_219 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_53_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_219 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_219 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_53_enex5
        ) begin
      reg_act_config_inst_counter_enexo_219 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_14_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2582_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_53_enex5
        ) begin
      reg_act_regs_data_2_14_2_enexo_5 <= act_regs_data_and_2582_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_14_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2534_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_53_enex5
        ) begin
      reg_act_regs_data_3_14_2_enexo_5 <= act_regs_data_and_2534_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_14_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2630_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_53_enex5
        ) begin
      reg_act_regs_data_1_14_2_enexo_5 <= act_regs_data_and_2630_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_220 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_54_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_220 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_220 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_54_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_220 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_220 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_54_enex5
        ) begin
      reg_act_config_inst_counter_enexo_220 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_14_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2679_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_54_enex5
        ) begin
      reg_act_regs_data_0_14_3_enexo_5 <= act_regs_data_and_2679_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_14_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2583_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_54_enex5
        ) begin
      reg_act_regs_data_2_14_3_enexo_5 <= act_regs_data_and_2583_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_14_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2535_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_54_enex5
        ) begin
      reg_act_regs_data_3_14_3_enexo_5 <= act_regs_data_and_2535_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_14_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2631_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_54_enex5
        ) begin
      reg_act_regs_data_1_14_3_enexo_5 <= act_regs_data_and_2631_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_221 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_55_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_221 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_14_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2629_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_55_enex5
        ) begin
      reg_act_regs_data_1_14_1_enexo_5 <= act_regs_data_and_2629_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_221 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_55_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_221 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_221 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_55_enex5
        ) begin
      reg_act_config_inst_counter_enexo_221 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_14_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2581_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_55_enex5
        ) begin
      reg_act_regs_data_2_14_1_enexo_5 <= act_regs_data_and_2581_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_14_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2533_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_55_enex5
        ) begin
      reg_act_regs_data_3_14_1_enexo_5 <= act_regs_data_and_2533_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_14_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2677_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_55_enex5
        ) begin
      reg_act_regs_data_0_14_1_enexo_5 <= act_regs_data_and_2677_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_222 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_56_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_222 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_222 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_56_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_222 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_222 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_56_enex5
        ) begin
      reg_act_config_inst_counter_enexo_222 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_15_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2531_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_56_enex5
        ) begin
      reg_act_regs_data_3_15_2_enexo_5 <= act_regs_data_and_2531_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_15_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2579_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_56_enex5
        ) begin
      reg_act_regs_data_2_15_2_enexo_5 <= act_regs_data_and_2579_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_15_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2675_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_56_enex5
        ) begin
      reg_act_regs_data_0_15_2_enexo_5 <= act_regs_data_and_2675_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_15_2_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2627_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_56_enex5
        ) begin
      reg_act_regs_data_1_15_2_enexo_5 <= act_regs_data_and_2627_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_223 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_57_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_223 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_223 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_57_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_223 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_15_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2580_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_57_enex5
        ) begin
      reg_act_regs_data_2_15_3_enexo_5 <= act_regs_data_and_2580_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_223 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_57_enex5
        ) begin
      reg_act_config_inst_counter_enexo_223 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_15_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2676_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_57_enex5
        ) begin
      reg_act_regs_data_0_15_3_enexo_5 <= act_regs_data_and_2676_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_15_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2628_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_57_enex5
        ) begin
      reg_act_regs_data_1_15_3_enexo_5 <= act_regs_data_and_2628_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_15_3_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2532_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_57_enex5
        ) begin
      reg_act_regs_data_3_15_3_enexo_5 <= act_regs_data_and_2532_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_224 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_20_cse | nv_scvector_cctor_nv_scvector_5_for_and_58_enex5
        ) begin
      reg_act_config_inst_regs_4_sva_dfm_5_enexo_224 <= act_config_inst_regs_and_20_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_224 <= 1'b1;
    end
    else if ( act_config_inst_regs_and_4_cse | nv_scvector_cctor_nv_scvector_5_for_and_58_enex5
        ) begin
      reg_act_config_inst_regs_20_sva_dfm_6_enexo_224 <= act_config_inst_regs_and_4_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_config_inst_counter_enexo_224 <= 1'b1;
    end
    else if ( act_config_inst_counter_and_tmp | nv_scvector_cctor_nv_scvector_5_for_and_58_enex5
        ) begin
      reg_act_config_inst_counter_enexo_224 <= act_config_inst_counter_and_tmp;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_15_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2674_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_58_enex5
        ) begin
      reg_act_regs_data_0_15_1_enexo_5 <= act_regs_data_and_2674_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_1_15_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2626_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_58_enex5
        ) begin
      reg_act_regs_data_1_15_1_enexo_5 <= act_regs_data_and_2626_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_2_15_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2578_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_58_enex5
        ) begin
      reg_act_regs_data_2_15_1_enexo_5 <= act_regs_data_and_2578_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_3_15_1_enexo_5 <= 1'b1;
    end
    else if ( act_regs_data_and_2530_enex5 | nv_scvector_cctor_nv_scvector_5_for_and_58_enex5
        ) begin
      reg_act_regs_data_3_15_1_enexo_5 <= act_regs_data_and_2530_enex5;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_29_24_sva_dfm_6_3 <= 1'b0;
      rva_out_reg_data_29_24_sva_dfm_6_2_0 <= 3'b000;
    end
    else if ( rva_out_reg_data_and_61_tmp ) begin
      rva_out_reg_data_29_24_sva_dfm_6_3 <= MUX1HOT_s_1_5_2((Silu_for_12_else_else_else_else_if_acc_sdt[3]),
          ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_25_22_mx0w2_3,
          nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_6_nl, (act_mem_banks_read_read_data_lpi_1_dfm_1_31_0[27]),
          rva_out_reg_data_29_24_sva_dfm_3_3, {and_dcpl_331 , and_dcpl_1390 , and_dcpl_1236
          , and_dcpl_1094 , and_dcpl_1096});
      rva_out_reg_data_29_24_sva_dfm_6_2_0 <= MUX1HOT_v_3_5_2((Silu_for_12_else_else_else_else_if_acc_sdt[2:0]),
          ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_25_22_mx0w2_2_0,
          nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_304_nl, (act_mem_banks_read_read_data_lpi_1_dfm_1_31_0[26:24]),
          rva_out_reg_data_29_24_sva_dfm_3_2_0, {and_dcpl_331 , and_dcpl_1390 , and_dcpl_1236
          , and_dcpl_1094 , and_dcpl_1096});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rva_out_reg_data_39_32_sva_dfm_6_3 <= 1'b0;
      rva_out_reg_data_39_32_sva_dfm_6_2_0 <= 3'b000;
    end
    else if ( and_1801_tmp ) begin
      rva_out_reg_data_39_32_sva_dfm_6_3 <= MUX1HOT_s_1_3_2(and_1711_nl, (act_mem_banks_read_read_data_lpi_1_dfm_1_63_32[3]),
          rva_out_reg_data_39_32_sva_dfm_3_3, {rva_out_reg_data_39_32_sva_dfm_6_mx0c0
          , and_dcpl_1094 , and_dcpl_1096});
      rva_out_reg_data_39_32_sva_dfm_6_2_0 <= MUX1HOT_v_3_3_2(and_3505_nl, (act_mem_banks_read_read_data_lpi_1_dfm_1_63_32[2:0]),
          rva_out_reg_data_39_32_sva_dfm_3_2_0, {rva_out_reg_data_39_32_sva_dfm_6_mx0c0
          , and_dcpl_1094 , and_dcpl_1096});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_15_sva_25 <= 1'b0;
      act_regs_data_3_15_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2531_enex5 ) begin
      act_regs_data_3_15_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_3_15_sva_dfm_2_25_22_rsp_0,
          act_regs_data_2_2_sva_8_25, act_regs_data_3_15_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_3_15_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_3_15_sva_dfm_2_25_22_rsp_1,
          act_regs_data_2_2_sva_8_24_22, act_regs_data_3_15_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_14_sva_25 <= 1'b0;
      act_regs_data_3_14_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2534_enex5 ) begin
      act_regs_data_3_14_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_3_14_sva_dfm_2_25_22_rsp_0,
          act_regs_data_2_15_sva_8_25, act_regs_data_3_14_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_3_14_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_3_14_sva_dfm_2_25_22_rsp_1,
          act_regs_data_2_15_sva_8_24_22, act_regs_data_3_14_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_13_sva_25 <= 1'b0;
      act_regs_data_3_13_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2537_enex5 ) begin
      act_regs_data_3_13_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_3_13_sva_dfm_2_25_22_rsp_0,
          act_regs_data_2_14_sva_8_25, act_regs_data_3_13_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_3_13_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_3_13_sva_dfm_2_25_22_rsp_1,
          act_regs_data_2_14_sva_8_24_22, act_regs_data_3_13_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_12_sva_25 <= 1'b0;
      act_regs_data_3_12_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2540_enex5 ) begin
      act_regs_data_3_12_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_3_12_sva_dfm_2_25_22_rsp_0,
          act_regs_data_2_13_sva_8_25, act_regs_data_3_12_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_3_12_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_3_12_sva_dfm_2_25_22_rsp_1,
          act_regs_data_2_13_sva_8_24_22, act_regs_data_3_12_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_11_sva_25 <= 1'b0;
      act_regs_data_3_11_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2543_enex5 ) begin
      act_regs_data_3_11_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_3_11_sva_dfm_2_25_22_rsp_0,
          act_regs_data_2_12_sva_8_25, act_regs_data_3_11_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_3_11_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_3_11_sva_dfm_2_25_22_rsp_1,
          act_regs_data_2_12_sva_8_24_22, act_regs_data_3_11_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_10_sva_25 <= 1'b0;
      act_regs_data_3_10_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2546_enex5 ) begin
      act_regs_data_3_10_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_3_10_sva_dfm_2_25_22_rsp_0,
          act_regs_data_2_11_sva_8_25, act_regs_data_3_10_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_3_10_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_3_10_sva_dfm_2_25_22_rsp_1,
          act_regs_data_2_11_sva_8_24_22, act_regs_data_3_10_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_9_sva_25 <= 1'b0;
      act_regs_data_3_9_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2549_enex5 ) begin
      act_regs_data_3_9_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_3_9_sva_dfm_2_25_22_rsp_0,
          act_regs_data_3_0_sva_8_25, act_regs_data_3_9_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_3_9_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_3_9_sva_dfm_2_25_22_rsp_1,
          act_regs_data_3_0_sva_8_24_22, act_regs_data_3_9_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_8_sva_25 <= 1'b0;
      act_regs_data_3_8_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2552_enex5 ) begin
      act_regs_data_3_8_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_3_8_sva_dfm_2_25_22_rsp_0,
          act_regs_data_2_9_sva_8_25, act_regs_data_3_8_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_3_8_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_3_8_sva_dfm_2_25_22_rsp_1,
          act_regs_data_2_9_sva_8_24_22, act_regs_data_3_8_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_7_sva_25 <= 1'b0;
      act_regs_data_3_7_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2555_enex5 ) begin
      act_regs_data_3_7_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_3_7_sva_dfm_2_25_22_rsp_0,
          act_regs_data_2_8_sva_8_25, act_regs_data_3_7_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_3_7_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_3_7_sva_dfm_2_25_22_rsp_1,
          act_regs_data_2_8_sva_8_24_22, act_regs_data_3_7_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_6_sva_25 <= 1'b0;
      act_regs_data_3_6_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2558_enex5 ) begin
      act_regs_data_3_6_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_3_6_sva_dfm_2_25_22_rsp_0,
          act_regs_data_2_7_sva_8_25, act_regs_data_3_6_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_3_6_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_3_6_sva_dfm_2_25_22_rsp_1,
          act_regs_data_2_7_sva_8_24_22, act_regs_data_3_6_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_5_sva_25 <= 1'b0;
      act_regs_data_3_5_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2561_enex5 ) begin
      act_regs_data_3_5_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_3_5_sva_dfm_2_25_22_rsp_0,
          act_regs_data_2_6_sva_8_25, act_regs_data_3_5_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_3_5_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_3_5_sva_dfm_2_25_22_rsp_1,
          act_regs_data_2_6_sva_8_24_22, act_regs_data_3_5_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_4_sva_25 <= 1'b0;
      act_regs_data_3_4_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2564_enex5 ) begin
      act_regs_data_3_4_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_3_4_sva_dfm_2_25_22_rsp_0,
          act_regs_data_2_5_sva_8_25, act_regs_data_3_4_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_3_4_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_3_4_sva_dfm_2_25_22_rsp_1,
          act_regs_data_2_5_sva_8_24_22, act_regs_data_3_4_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_3_sva_25 <= 1'b0;
      act_regs_data_3_3_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2567_enex5 ) begin
      act_regs_data_3_3_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_3_3_sva_dfm_2_25_22_rsp_0,
          act_regs_data_2_4_sva_8_25, act_regs_data_3_3_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_3_3_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_3_3_sva_dfm_2_25_22_rsp_1,
          act_regs_data_2_4_sva_8_24_22, act_regs_data_3_3_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_2_sva_25 <= 1'b0;
      act_regs_data_3_2_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2570_enex5 ) begin
      act_regs_data_3_2_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_3_2_sva_dfm_2_25_22_rsp_0,
          act_regs_data_2_3_sva_8_25, act_regs_data_3_2_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_3_2_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_3_2_sva_dfm_2_25_22_rsp_1,
          act_regs_data_2_3_sva_8_24_22, act_regs_data_3_2_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_1_sva_25 <= 1'b0;
      act_regs_data_3_1_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2573_enex5 ) begin
      act_regs_data_3_1_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_3_1_sva_dfm_2_25_22_rsp_0,
          act_regs_data_2_10_sva_8_25, act_regs_data_3_1_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_3_1_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_3_1_sva_dfm_2_25_22_rsp_1,
          act_regs_data_2_10_sva_8_24_22, act_regs_data_3_1_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_0_sva_25 <= 1'b0;
      act_regs_data_3_0_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2576_enex5 ) begin
      act_regs_data_3_0_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_3_0_sva_dfm_2_25_22_rsp_0,
          act_regs_data_2_1_sva_8_25, act_regs_data_3_0_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_3_0_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_3_0_sva_dfm_2_25_22_rsp_1,
          act_regs_data_2_1_sva_8_24_22, act_regs_data_3_0_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_15_sva_25 <= 1'b0;
      act_regs_data_2_15_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2579_enex5 ) begin
      act_regs_data_2_15_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_2_15_sva_dfm_2_25_22_rsp_0,
          act_regs_data_1_2_sva_8_25, act_regs_data_2_15_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_2_15_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_2_15_sva_dfm_2_25_22_rsp_1,
          act_regs_data_1_2_sva_8_24_22, act_regs_data_2_15_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_14_sva_25 <= 1'b0;
      act_regs_data_2_14_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2582_enex5 ) begin
      act_regs_data_2_14_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_2_14_sva_dfm_2_25_22_rsp_0,
          act_regs_data_1_15_sva_8_25, act_regs_data_2_14_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_2_14_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_2_14_sva_dfm_2_25_22_rsp_1,
          act_regs_data_1_15_sva_8_24_22, act_regs_data_2_14_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_13_sva_25 <= 1'b0;
      act_regs_data_2_13_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2585_enex5 ) begin
      act_regs_data_2_13_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_2_13_sva_dfm_2_25_22_rsp_0,
          act_regs_data_1_14_sva_8_25, act_regs_data_2_13_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_2_13_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_2_13_sva_dfm_2_25_22_rsp_1,
          act_regs_data_1_14_sva_8_24_22, act_regs_data_2_13_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_12_sva_25 <= 1'b0;
      act_regs_data_2_12_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2588_enex5 ) begin
      act_regs_data_2_12_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_2_12_sva_dfm_2_25_22_rsp_0,
          act_regs_data_1_13_sva_8_25, act_regs_data_2_12_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_2_12_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_2_12_sva_dfm_2_25_22_rsp_1,
          act_regs_data_1_13_sva_8_24_22, act_regs_data_2_12_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_11_sva_25 <= 1'b0;
      act_regs_data_2_11_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2591_enex5 ) begin
      act_regs_data_2_11_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_2_11_sva_dfm_2_25_22_rsp_0,
          act_regs_data_1_12_sva_8_25, act_regs_data_2_11_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_2_11_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_2_11_sva_dfm_2_25_22_rsp_1,
          act_regs_data_1_12_sva_8_24_22, act_regs_data_2_11_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_10_sva_25 <= 1'b0;
      act_regs_data_2_10_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2594_enex5 ) begin
      act_regs_data_2_10_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_2_10_sva_dfm_2_25_22_rsp_0,
          act_regs_data_1_11_sva_8_25, act_regs_data_2_10_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_2_10_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_2_10_sva_dfm_2_25_22_rsp_1,
          act_regs_data_1_11_sva_8_24_22, act_regs_data_2_10_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_9_sva_25 <= 1'b0;
      act_regs_data_2_9_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2597_enex5 ) begin
      act_regs_data_2_9_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_2_9_sva_dfm_2_25_22_rsp_0,
          act_regs_data_2_0_sva_8_25, act_regs_data_2_9_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_2_9_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_2_9_sva_dfm_2_25_22_rsp_1,
          act_regs_data_2_0_sva_8_24_22, act_regs_data_2_9_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_8_sva_25 <= 1'b0;
      act_regs_data_2_8_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2600_enex5 ) begin
      act_regs_data_2_8_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_2_8_sva_dfm_2_25_22_rsp_0,
          act_regs_data_1_9_sva_8_25, act_regs_data_2_8_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_2_8_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_2_8_sva_dfm_2_25_22_rsp_1,
          act_regs_data_1_9_sva_8_24_22, act_regs_data_2_8_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_7_sva_25 <= 1'b0;
      act_regs_data_2_7_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2603_enex5 ) begin
      act_regs_data_2_7_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_2_7_sva_dfm_2_25_22_rsp_0,
          act_regs_data_1_8_sva_8_25, act_regs_data_2_7_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_2_7_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_2_7_sva_dfm_2_25_22_rsp_1,
          act_regs_data_1_8_sva_8_24_22, act_regs_data_2_7_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_6_sva_25 <= 1'b0;
      act_regs_data_2_6_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2606_enex5 ) begin
      act_regs_data_2_6_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_2_6_sva_dfm_2_25_22_rsp_0,
          act_regs_data_1_7_sva_8_25, act_regs_data_2_6_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_2_6_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_2_6_sva_dfm_2_25_22_rsp_1,
          act_regs_data_1_7_sva_8_24_22, act_regs_data_2_6_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_5_sva_25 <= 1'b0;
      act_regs_data_2_5_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2609_enex5 ) begin
      act_regs_data_2_5_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_2_5_sva_dfm_2_25_22_rsp_0,
          act_regs_data_1_6_sva_8_25, act_regs_data_2_5_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_2_5_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_2_5_sva_dfm_2_25_22_rsp_1,
          act_regs_data_1_6_sva_8_24_22, act_regs_data_2_5_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_4_sva_25 <= 1'b0;
      act_regs_data_2_4_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2612_enex5 ) begin
      act_regs_data_2_4_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_2_4_sva_dfm_2_25_22_rsp_0,
          act_regs_data_1_5_sva_8_25, act_regs_data_2_4_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_2_4_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_2_4_sva_dfm_2_25_22_rsp_1,
          act_regs_data_1_5_sva_8_24_22, act_regs_data_2_4_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_3_sva_25 <= 1'b0;
      act_regs_data_2_3_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2615_enex5 ) begin
      act_regs_data_2_3_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_2_3_sva_dfm_2_25_22_rsp_0,
          act_regs_data_1_4_sva_8_25, act_regs_data_2_3_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_2_3_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_2_3_sva_dfm_2_25_22_rsp_1,
          act_regs_data_1_4_sva_8_24_22, act_regs_data_2_3_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_2_sva_25 <= 1'b0;
      act_regs_data_2_2_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2618_enex5 ) begin
      act_regs_data_2_2_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_2_2_sva_dfm_2_25_22_rsp_0,
          act_regs_data_1_3_sva_8_25, act_regs_data_2_2_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_2_2_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_2_2_sva_dfm_2_25_22_rsp_1,
          act_regs_data_1_3_sva_8_24_22, act_regs_data_2_2_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_1_sva_25 <= 1'b0;
      act_regs_data_2_1_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2621_enex5 ) begin
      act_regs_data_2_1_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_2_1_sva_dfm_2_25_22_rsp_0,
          act_regs_data_1_10_sva_8_25, act_regs_data_2_1_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_2_1_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_2_1_sva_dfm_2_25_22_rsp_1,
          act_regs_data_1_10_sva_8_24_22, act_regs_data_2_1_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_2_0_sva_25 <= 1'b0;
      act_regs_data_2_0_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2624_enex5 ) begin
      act_regs_data_2_0_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_2_0_sva_dfm_2_25_22_rsp_0,
          act_regs_data_1_1_sva_8_25, act_regs_data_2_0_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_2_0_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_2_0_sva_dfm_2_25_22_rsp_1,
          act_regs_data_1_1_sva_8_24_22, act_regs_data_2_0_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_15_sva_25 <= 1'b0;
      act_regs_data_1_15_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2627_enex5 ) begin
      act_regs_data_1_15_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_1_15_sva_dfm_2_25_22_rsp_0,
          act_regs_data_0_2_sva_8_25, act_regs_data_1_15_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_1_15_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_1_15_sva_dfm_2_25_22_rsp_1,
          act_regs_data_0_2_sva_8_24_22, act_regs_data_1_15_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_14_sva_25 <= 1'b0;
      act_regs_data_1_14_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2630_enex5 ) begin
      act_regs_data_1_14_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_1_14_sva_dfm_2_25_22_rsp_0,
          act_regs_data_0_15_sva_8_25, act_regs_data_1_14_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_1_14_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_1_14_sva_dfm_2_25_22_rsp_1,
          act_regs_data_0_15_sva_8_24_22, act_regs_data_1_14_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_13_sva_25 <= 1'b0;
      act_regs_data_1_13_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2633_enex5 ) begin
      act_regs_data_1_13_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_1_13_sva_dfm_2_25_22_rsp_0,
          act_regs_data_0_14_sva_8_25, act_regs_data_1_13_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_1_13_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_1_13_sva_dfm_2_25_22_rsp_1,
          act_regs_data_0_14_sva_8_24_22, act_regs_data_1_13_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_12_sva_25 <= 1'b0;
      act_regs_data_1_12_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2636_enex5 ) begin
      act_regs_data_1_12_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_1_12_sva_dfm_2_25_22_rsp_0,
          act_regs_data_0_13_sva_8_25, act_regs_data_1_12_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_1_12_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_1_12_sva_dfm_2_25_22_rsp_1,
          act_regs_data_0_13_sva_8_24_22, act_regs_data_1_12_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_11_sva_25 <= 1'b0;
      act_regs_data_1_11_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2639_enex5 ) begin
      act_regs_data_1_11_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_1_11_sva_dfm_2_25_22_rsp_0,
          act_regs_data_0_12_sva_8_25, act_regs_data_1_11_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_1_11_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_1_11_sva_dfm_2_25_22_rsp_1,
          act_regs_data_0_12_sva_8_24_22, act_regs_data_1_11_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_10_sva_25 <= 1'b0;
      act_regs_data_1_10_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2642_enex5 ) begin
      act_regs_data_1_10_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_1_10_sva_dfm_2_25_22_rsp_0,
          act_regs_data_0_11_sva_8_25, act_regs_data_1_10_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_1_10_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_1_10_sva_dfm_2_25_22_rsp_1,
          act_regs_data_0_11_sva_8_24_22, act_regs_data_1_10_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_9_sva_25 <= 1'b0;
      act_regs_data_1_9_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2645_enex5 ) begin
      act_regs_data_1_9_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_1_9_sva_dfm_2_25_22_rsp_0,
          act_regs_data_1_0_sva_8_25, act_regs_data_1_9_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_1_9_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_1_9_sva_dfm_2_25_22_rsp_1,
          act_regs_data_1_0_sva_8_24_22, act_regs_data_1_9_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_8_sva_25 <= 1'b0;
      act_regs_data_1_8_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2648_enex5 ) begin
      act_regs_data_1_8_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_1_8_sva_dfm_2_25_22_rsp_0,
          act_regs_data_0_9_sva_8_25, act_regs_data_1_8_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_1_8_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_1_8_sva_dfm_2_25_22_rsp_1,
          act_regs_data_0_9_sva_8_24_22, act_regs_data_1_8_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_7_sva_25 <= 1'b0;
      act_regs_data_1_7_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2651_enex5 ) begin
      act_regs_data_1_7_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_1_7_sva_dfm_2_25_22_rsp_0,
          act_regs_data_0_8_sva_8_25, act_regs_data_1_7_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_1_7_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_1_7_sva_dfm_2_25_22_rsp_1,
          act_regs_data_0_8_sva_8_24_22, act_regs_data_1_7_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_6_sva_25 <= 1'b0;
      act_regs_data_1_6_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2654_enex5 ) begin
      act_regs_data_1_6_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_1_6_sva_dfm_2_25_22_rsp_0,
          act_regs_data_0_7_sva_8_25, act_regs_data_1_6_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_1_6_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_1_6_sva_dfm_2_25_22_rsp_1,
          act_regs_data_0_7_sva_8_24_22, act_regs_data_1_6_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_5_sva_25 <= 1'b0;
      act_regs_data_1_5_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2657_enex5 ) begin
      act_regs_data_1_5_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_1_5_sva_dfm_2_25_22_rsp_0,
          act_regs_data_0_6_sva_8_25, act_regs_data_1_5_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_1_5_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_1_5_sva_dfm_2_25_22_rsp_1,
          act_regs_data_0_6_sva_8_24_22, act_regs_data_1_5_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_4_sva_25 <= 1'b0;
      act_regs_data_1_4_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2660_enex5 ) begin
      act_regs_data_1_4_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_1_4_sva_dfm_2_25_22_rsp_0,
          act_regs_data_0_5_sva_8_25, act_regs_data_1_4_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_1_4_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_1_4_sva_dfm_2_25_22_rsp_1,
          act_regs_data_0_5_sva_8_24_22, act_regs_data_1_4_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_3_sva_25 <= 1'b0;
      act_regs_data_1_3_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2663_enex5 ) begin
      act_regs_data_1_3_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_1_3_sva_dfm_2_25_22_rsp_0,
          act_regs_data_0_4_sva_8_25, act_regs_data_1_3_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_1_3_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_1_3_sva_dfm_2_25_22_rsp_1,
          act_regs_data_0_4_sva_8_24_22, act_regs_data_1_3_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_2_sva_25 <= 1'b0;
      act_regs_data_1_2_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2666_enex5 ) begin
      act_regs_data_1_2_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_1_2_sva_dfm_2_25_22_rsp_0,
          act_regs_data_0_3_sva_8_25, act_regs_data_1_2_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_1_2_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_1_2_sva_dfm_2_25_22_rsp_1,
          act_regs_data_0_3_sva_8_24_22, act_regs_data_1_2_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_1_sva_25 <= 1'b0;
      act_regs_data_1_1_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2669_enex5 ) begin
      act_regs_data_1_1_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_1_1_sva_dfm_2_25_22_rsp_0,
          act_regs_data_0_10_sva_8_25, act_regs_data_1_1_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_1_1_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_1_1_sva_dfm_2_25_22_rsp_1,
          act_regs_data_0_10_sva_8_24_22, act_regs_data_1_1_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_1_0_sva_25 <= 1'b0;
      act_regs_data_1_0_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2672_enex5 ) begin
      act_regs_data_1_0_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_1_0_sva_dfm_2_25_22_rsp_0,
          act_regs_data_0_1_sva_8_25, act_regs_data_1_0_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_1_0_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_1_0_sva_dfm_2_25_22_rsp_1,
          act_regs_data_0_1_sva_8_24_22, act_regs_data_1_0_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_15_sva_25 <= 1'b0;
      act_regs_data_0_15_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2675_enex5 ) begin
      act_regs_data_0_15_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_0_15_sva_dfm_2_25_22_rsp_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_1_25, act_regs_data_0_15_sva_8_25,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_0_15_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_0_15_sva_dfm_2_25_22_rsp_1,
          ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_1_24_22, act_regs_data_0_15_sva_8_24_22,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_14_sva_25 <= 1'b0;
      act_regs_data_0_14_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2678_enex5 ) begin
      act_regs_data_0_14_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_0_14_sva_dfm_2_25_22_rsp_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_1_25, act_regs_data_0_14_sva_8_25,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_0_14_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_0_14_sva_dfm_2_25_22_rsp_1,
          ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_1_24_22, act_regs_data_0_14_sva_8_24_22,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_9_sva_25 <= 1'b0;
      act_regs_data_0_9_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2681_enex5 ) begin
      act_regs_data_0_9_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_0_9_sva_dfm_2_25_22_rsp_0,
          act_regs_data_0_0_sva_8_25, act_regs_data_0_9_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_0_9_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_0_9_sva_dfm_2_25_22_rsp_1,
          act_regs_data_0_0_sva_8_24_22, act_regs_data_0_9_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_8_sva_25 <= 1'b0;
      act_regs_data_0_8_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2684_enex5 ) begin
      act_regs_data_0_8_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_0_8_sva_dfm_2_25_22_rsp_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_1_25, act_regs_data_0_8_sva_8_25,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_0_8_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_0_8_sva_dfm_2_25_22_rsp_1,
          ActUnit_PushOutput_if_output_port_reg_data_data_9_sva_1_24_22, act_regs_data_0_8_sva_8_24_22,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_7_sva_25 <= 1'b0;
      act_regs_data_0_7_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2687_enex5 ) begin
      act_regs_data_0_7_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_0_7_sva_dfm_2_25_22_rsp_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_1_25, act_regs_data_0_7_sva_8_25,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_0_7_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_0_7_sva_dfm_2_25_22_rsp_1,
          ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_1_24_22, act_regs_data_0_7_sva_8_24_22,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_6_sva_25 <= 1'b0;
      act_regs_data_0_6_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2690_enex5 ) begin
      act_regs_data_0_6_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_0_6_sva_dfm_2_25_22_rsp_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_1_25, act_regs_data_0_6_sva_8_25,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_0_6_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_0_6_sva_dfm_2_25_22_rsp_1,
          ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_1_24_22, act_regs_data_0_6_sva_8_24_22,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_5_sva_25 <= 1'b0;
      act_regs_data_0_5_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2693_enex5 ) begin
      act_regs_data_0_5_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_0_5_sva_dfm_2_25_22_rsp_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_1_25, act_regs_data_0_5_sva_8_25,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_0_5_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_0_5_sva_dfm_2_25_22_rsp_1,
          ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_1_24_22, act_regs_data_0_5_sva_8_24_22,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_4_sva_25 <= 1'b0;
      act_regs_data_0_4_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2696_enex5 ) begin
      act_regs_data_0_4_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_0_4_sva_dfm_2_25_22_rsp_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_1_25, act_regs_data_0_4_sva_8_25,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_0_4_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_0_4_sva_dfm_2_25_22_rsp_1,
          ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_1_24_22, act_regs_data_0_4_sva_8_24_22,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_3_sva_25 <= 1'b0;
      act_regs_data_0_3_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2699_enex5 ) begin
      act_regs_data_0_3_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_0_3_sva_dfm_2_25_22_rsp_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_1_25, act_regs_data_0_3_sva_8_25,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_0_3_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_0_3_sva_dfm_2_25_22_rsp_1,
          ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_1_24_22, act_regs_data_0_3_sva_8_24_22,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_0_2_sva_25 <= 1'b0;
      act_regs_data_0_2_sva_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2702_enex5 ) begin
      act_regs_data_0_2_sva_25 <= MUX1HOT_s_1_3_2(act_regs_data_0_2_sva_dfm_2_25_22_rsp_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_1_25, act_regs_data_0_2_sva_8_25,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      act_regs_data_0_2_sva_24_22 <= MUX1HOT_v_3_3_2(act_regs_data_0_2_sva_dfm_2_25_22_rsp_1,
          ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_1_24_22, act_regs_data_0_2_sva_8_24_22,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22
          <= 3'b000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_38_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25
          <= MUX_s_1_4_2(act_regs_data_0_15_sva_25, act_regs_data_1_15_sva_25, act_regs_data_2_15_sva_25,
          act_regs_data_3_15_sva_25, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22
          <= MUX_v_3_4_2(act_regs_data_0_15_sva_24_22, act_regs_data_1_15_sva_24_22,
          act_regs_data_2_15_sva_24_22, act_regs_data_3_15_sva_24_22, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22
          <= 3'b000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_41_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25
          <= MUX_s_1_4_2(act_regs_data_0_14_sva_25, act_regs_data_1_14_sva_25, act_regs_data_2_14_sva_25,
          act_regs_data_3_14_sva_25, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22
          <= MUX_v_3_4_2(act_regs_data_0_14_sva_24_22, act_regs_data_1_14_sva_24_22,
          act_regs_data_2_14_sva_24_22, act_regs_data_3_14_sva_24_22, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22
          <= 3'b000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_44_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25
          <= MUX_s_1_4_2(reg_act_regs_data_0_13_ftd_2_3, act_regs_data_1_13_sva_25,
          act_regs_data_2_13_sva_25, act_regs_data_3_13_sva_25, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22
          <= MUX_v_3_4_2(reg_act_regs_data_0_13_ftd_2_2_0, act_regs_data_1_13_sva_24_22,
          act_regs_data_2_13_sva_24_22, act_regs_data_3_13_sva_24_22, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22
          <= 3'b000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_47_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25
          <= MUX_s_1_4_2(reg_act_regs_data_0_12_ftd_2_3, act_regs_data_1_12_sva_25,
          act_regs_data_2_12_sva_25, act_regs_data_3_12_sva_25, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22
          <= MUX_v_3_4_2(reg_act_regs_data_0_12_ftd_2_2_0, act_regs_data_1_12_sva_24_22,
          act_regs_data_2_12_sva_24_22, act_regs_data_3_12_sva_24_22, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22
          <= 3'b000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_50_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25
          <= MUX_s_1_4_2(reg_act_regs_data_0_11_ftd_2_3, act_regs_data_1_11_sva_25,
          act_regs_data_2_11_sva_25, act_regs_data_3_11_sva_25, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22
          <= MUX_v_3_4_2(reg_act_regs_data_0_11_ftd_2_2_0, act_regs_data_1_11_sva_24_22,
          act_regs_data_2_11_sva_24_22, act_regs_data_3_11_sva_24_22, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22
          <= 3'b000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_53_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25
          <= MUX_s_1_4_2(reg_act_regs_data_0_10_ftd_2_3, act_regs_data_1_10_sva_25,
          act_regs_data_2_10_sva_25, act_regs_data_3_10_sva_25, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22
          <= MUX_v_3_4_2(reg_act_regs_data_0_10_ftd_2_2_0, act_regs_data_1_10_sva_24_22,
          act_regs_data_2_10_sva_24_22, act_regs_data_3_10_sva_24_22, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22
          <= 3'b000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_56_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25
          <= MUX_s_1_4_2(act_regs_data_0_9_sva_25, act_regs_data_1_9_sva_25, act_regs_data_2_9_sva_25,
          act_regs_data_3_9_sva_25, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22
          <= MUX_v_3_4_2(act_regs_data_0_9_sva_24_22, act_regs_data_1_9_sva_24_22,
          act_regs_data_2_9_sva_24_22, act_regs_data_3_9_sva_24_22, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22
          <= 3'b000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_59_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25
          <= MUX_s_1_4_2(act_regs_data_0_8_sva_25, act_regs_data_1_8_sva_25, act_regs_data_2_8_sva_25,
          act_regs_data_3_8_sva_25, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22
          <= MUX_v_3_4_2(act_regs_data_0_8_sva_24_22, act_regs_data_1_8_sva_24_22,
          act_regs_data_2_8_sva_24_22, act_regs_data_3_8_sva_24_22, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22
          <= 3'b000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_62_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25
          <= MUX_s_1_4_2(act_regs_data_0_7_sva_25, act_regs_data_1_7_sva_25, act_regs_data_2_7_sva_25,
          act_regs_data_3_7_sva_25, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22
          <= MUX_v_3_4_2(act_regs_data_0_7_sva_24_22, act_regs_data_1_7_sva_24_22,
          act_regs_data_2_7_sva_24_22, act_regs_data_3_7_sva_24_22, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22
          <= 3'b000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_65_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25
          <= MUX_s_1_4_2(act_regs_data_0_6_sva_25, act_regs_data_1_6_sva_25, act_regs_data_2_6_sva_25,
          act_regs_data_3_6_sva_25, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22
          <= MUX_v_3_4_2(act_regs_data_0_6_sva_24_22, act_regs_data_1_6_sva_24_22,
          act_regs_data_2_6_sva_24_22, act_regs_data_3_6_sva_24_22, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22
          <= 3'b000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_68_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25
          <= MUX_s_1_4_2(act_regs_data_0_5_sva_25, act_regs_data_1_5_sva_25, act_regs_data_2_5_sva_25,
          act_regs_data_3_5_sva_25, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22
          <= MUX_v_3_4_2(act_regs_data_0_5_sva_24_22, act_regs_data_1_5_sva_24_22,
          act_regs_data_2_5_sva_24_22, act_regs_data_3_5_sva_24_22, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22
          <= 3'b000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_71_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25
          <= MUX_s_1_4_2(act_regs_data_0_4_sva_25, act_regs_data_1_4_sva_25, act_regs_data_2_4_sva_25,
          act_regs_data_3_4_sva_25, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22
          <= MUX_v_3_4_2(act_regs_data_0_4_sva_24_22, act_regs_data_1_4_sva_24_22,
          act_regs_data_2_4_sva_24_22, act_regs_data_3_4_sva_24_22, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22
          <= 3'b000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_74_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25
          <= MUX_s_1_4_2(act_regs_data_0_3_sva_25, act_regs_data_1_3_sva_25, act_regs_data_2_3_sva_25,
          act_regs_data_3_3_sva_25, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22
          <= MUX_v_3_4_2(act_regs_data_0_3_sva_24_22, act_regs_data_1_3_sva_24_22,
          act_regs_data_2_3_sva_24_22, act_regs_data_3_3_sva_24_22, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22
          <= 3'b000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_77_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25
          <= MUX_s_1_4_2(act_regs_data_0_2_sva_25, act_regs_data_1_2_sva_25, act_regs_data_2_2_sva_25,
          act_regs_data_3_2_sva_25, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22
          <= MUX_v_3_4_2(act_regs_data_0_2_sva_24_22, act_regs_data_1_2_sva_24_22,
          act_regs_data_2_2_sva_24_22, act_regs_data_3_2_sva_24_22, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22
          <= 3'b000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_80_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25
          <= MUX_s_1_4_2(reg_act_regs_data_0_1_ftd_2_3, act_regs_data_1_1_sva_25,
          act_regs_data_2_1_sva_25, act_regs_data_3_1_sva_25, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22
          <= MUX_v_3_4_2(reg_act_regs_data_0_1_ftd_2_2_0, act_regs_data_1_1_sva_24_22,
          act_regs_data_2_1_sva_24_22, act_regs_data_3_1_sva_24_22, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25
          <= 1'b0;
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22
          <= 3'b000;
    end
    else if ( nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_and_83_enex5
        ) begin
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_25
          <= MUX_s_1_4_2(reg_act_regs_data_0_0_ftd_2_3, act_regs_data_1_0_sva_25,
          act_regs_data_2_0_sva_25, act_regs_data_3_0_sva_25, act_config_in_InstFetch_mux_tmp[1:0]);
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_24_22
          <= MUX_v_3_4_2(reg_act_regs_data_0_0_ftd_2_2_0, act_regs_data_1_0_sva_24_22,
          act_regs_data_2_0_sva_24_22, act_regs_data_3_0_sva_24_22, act_config_in_InstFetch_mux_tmp[1:0]);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_RunInst_case_15_nv_scvector_cctor_data_0_ftd_rsp_0 <= 1'b0;
      reg_ActUnit_RunInst_case_15_nv_scvector_cctor_data_0_ftd_rsp_1 <= 3'b000;
    end
    else if ( ActUnit_RunInst_switch_lp_and_813_enex5 ) begin
      reg_ActUnit_RunInst_case_15_nv_scvector_cctor_data_0_ftd_rsp_0 <= nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
      reg_ActUnit_RunInst_case_15_nv_scvector_cctor_data_0_ftd_rsp_1 <= nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_2_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
          <= 1'b0;
      reg_nv_scvector_cctor_nv_scvector_6_for_2_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
          <= 3'b000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_2_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
          <= nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
      reg_nv_scvector_cctor_nv_scvector_6_for_2_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
          <= nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_3_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
          <= 1'b0;
      reg_nv_scvector_cctor_nv_scvector_6_for_3_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
          <= 3'b000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_17_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_3_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
          <= nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
      reg_nv_scvector_cctor_nv_scvector_6_for_3_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
          <= nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_4_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
          <= 1'b0;
      reg_nv_scvector_cctor_nv_scvector_6_for_4_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
          <= 3'b000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_20_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_4_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
          <= nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
      reg_nv_scvector_cctor_nv_scvector_6_for_4_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
          <= nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_5_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
          <= 1'b0;
      reg_nv_scvector_cctor_nv_scvector_6_for_5_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
          <= 3'b000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_23_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_5_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
          <= nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
      reg_nv_scvector_cctor_nv_scvector_6_for_5_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
          <= nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_6_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
          <= 1'b0;
      reg_nv_scvector_cctor_nv_scvector_6_for_6_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
          <= 3'b000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_26_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_6_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
          <= nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
      reg_nv_scvector_cctor_nv_scvector_6_for_6_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
          <= nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_7_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
          <= 1'b0;
      reg_nv_scvector_cctor_nv_scvector_6_for_7_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
          <= 3'b000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_29_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_7_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
          <= nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
      reg_nv_scvector_cctor_nv_scvector_6_for_7_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
          <= nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_8_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
          <= 1'b0;
      reg_nv_scvector_cctor_nv_scvector_6_for_8_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
          <= 3'b000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_32_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_8_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
          <= nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
      reg_nv_scvector_cctor_nv_scvector_6_for_8_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
          <= nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_9_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
          <= 1'b0;
      reg_nv_scvector_cctor_nv_scvector_6_for_9_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
          <= 3'b000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_35_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_9_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
          <= nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
      reg_nv_scvector_cctor_nv_scvector_6_for_9_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
          <= nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_10_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
          <= 1'b0;
      reg_nv_scvector_cctor_nv_scvector_6_for_10_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
          <= 3'b000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_38_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_10_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
          <= nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
      reg_nv_scvector_cctor_nv_scvector_6_for_10_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
          <= nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_11_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
          <= 1'b0;
      reg_nv_scvector_cctor_nv_scvector_6_for_11_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
          <= 3'b000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_41_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_11_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
          <= nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
      reg_nv_scvector_cctor_nv_scvector_6_for_11_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
          <= nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_12_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
          <= 1'b0;
      reg_nv_scvector_cctor_nv_scvector_6_for_12_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
          <= 3'b000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_44_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_12_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
          <= nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
      reg_nv_scvector_cctor_nv_scvector_6_for_12_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
          <= nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_13_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
          <= 1'b0;
      reg_nv_scvector_cctor_nv_scvector_6_for_13_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
          <= 3'b000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_47_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_13_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
          <= nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
      reg_nv_scvector_cctor_nv_scvector_6_for_13_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
          <= nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_14_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
          <= 1'b0;
      reg_nv_scvector_cctor_nv_scvector_6_for_14_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
          <= 3'b000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_50_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_14_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
          <= nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
      reg_nv_scvector_cctor_nv_scvector_6_for_14_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
          <= nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_15_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
          <= 1'b0;
      reg_nv_scvector_cctor_nv_scvector_6_for_15_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
          <= 3'b000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_53_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_15_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
          <= nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
      reg_nv_scvector_cctor_nv_scvector_6_for_15_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
          <= nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_16_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
          <= 1'b0;
      reg_nv_scvector_cctor_nv_scvector_6_for_16_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
          <= 3'b000;
    end
    else if ( nv_scvector_cctor_nv_scvector_6_for_and_56_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_6_for_16_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0
          <= nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
      reg_nv_scvector_cctor_nv_scvector_6_for_16_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1
          <= nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_15_sva_8_25 <= 1'b0;
      act_regs_data_3_15_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2705_enex5 ) begin
      act_regs_data_3_15_sva_8_25 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_3_15_sva_dfm_2_25_22_rsp_0, or_dcpl_850);
      act_regs_data_3_15_sva_8_24_22 <= MUX_v_3_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_3_15_sva_dfm_2_25_22_rsp_1, or_dcpl_850);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_14_sva_8_25 <= 1'b0;
      act_regs_data_3_14_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2708_enex5 ) begin
      act_regs_data_3_14_sva_8_25 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_3_14_sva_dfm_2_25_22_rsp_0, or_dcpl_852);
      act_regs_data_3_14_sva_8_24_22 <= MUX_v_3_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_3_14_sva_dfm_2_25_22_rsp_1, or_dcpl_852);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_13_sva_8_25 <= 1'b0;
      act_regs_data_3_13_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2711_enex5 ) begin
      act_regs_data_3_13_sva_8_25 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_3_13_sva_dfm_2_25_22_rsp_0, or_dcpl_855);
      act_regs_data_3_13_sva_8_24_22 <= MUX_v_3_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_3_13_sva_dfm_2_25_22_rsp_1, or_dcpl_855);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_12_sva_8_25 <= 1'b0;
      act_regs_data_3_12_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2714_enex5 ) begin
      act_regs_data_3_12_sva_8_25 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_3_12_sva_dfm_2_25_22_rsp_0, or_dcpl_857);
      act_regs_data_3_12_sva_8_24_22 <= MUX_v_3_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_3_12_sva_dfm_2_25_22_rsp_1, or_dcpl_857);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_11_sva_8_25 <= 1'b0;
      act_regs_data_3_11_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2717_enex5 ) begin
      act_regs_data_3_11_sva_8_25 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_3_11_sva_dfm_2_25_22_rsp_0, or_dcpl_860);
      act_regs_data_3_11_sva_8_24_22 <= MUX_v_3_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_3_11_sva_dfm_2_25_22_rsp_1, or_dcpl_860);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_10_sva_8_25 <= 1'b0;
      act_regs_data_3_10_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2720_enex5 ) begin
      act_regs_data_3_10_sva_8_25 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_3_10_sva_dfm_2_25_22_rsp_0, or_dcpl_862);
      act_regs_data_3_10_sva_8_24_22 <= MUX_v_3_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_3_10_sva_dfm_2_25_22_rsp_1, or_dcpl_862);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_9_sva_8_25 <= 1'b0;
      act_regs_data_3_9_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2723_enex5 ) begin
      act_regs_data_3_9_sva_8_25 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_3_9_sva_dfm_2_25_22_rsp_0, or_dcpl_865);
      act_regs_data_3_9_sva_8_24_22 <= MUX_v_3_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_3_9_sva_dfm_2_25_22_rsp_1, or_dcpl_865);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_8_sva_8_25 <= 1'b0;
      act_regs_data_3_8_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2726_enex5 ) begin
      act_regs_data_3_8_sva_8_25 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_3_8_sva_dfm_2_25_22_rsp_0, or_dcpl_867);
      act_regs_data_3_8_sva_8_24_22 <= MUX_v_3_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_3_8_sva_dfm_2_25_22_rsp_1, or_dcpl_867);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_7_sva_8_25 <= 1'b0;
      act_regs_data_3_7_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2729_enex5 ) begin
      act_regs_data_3_7_sva_8_25 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_3_7_sva_dfm_2_25_22_rsp_0, or_dcpl_869);
      act_regs_data_3_7_sva_8_24_22 <= MUX_v_3_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_3_7_sva_dfm_2_25_22_rsp_1, or_dcpl_869);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_6_sva_8_25 <= 1'b0;
      act_regs_data_3_6_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2732_enex5 ) begin
      act_regs_data_3_6_sva_8_25 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_3_6_sva_dfm_2_25_22_rsp_0, or_dcpl_870);
      act_regs_data_3_6_sva_8_24_22 <= MUX_v_3_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_3_6_sva_dfm_2_25_22_rsp_1, or_dcpl_870);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_5_sva_8_25 <= 1'b0;
      act_regs_data_3_5_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2735_enex5 ) begin
      act_regs_data_3_5_sva_8_25 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_3_5_sva_dfm_2_25_22_rsp_0, or_dcpl_871);
      act_regs_data_3_5_sva_8_24_22 <= MUX_v_3_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_3_5_sva_dfm_2_25_22_rsp_1, or_dcpl_871);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_4_sva_8_25 <= 1'b0;
      act_regs_data_3_4_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2738_enex5 ) begin
      act_regs_data_3_4_sva_8_25 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_3_4_sva_dfm_2_25_22_rsp_0, or_dcpl_872);
      act_regs_data_3_4_sva_8_24_22 <= MUX_v_3_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_3_4_sva_dfm_2_25_22_rsp_1, or_dcpl_872);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_3_sva_8_25 <= 1'b0;
      act_regs_data_3_3_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2741_enex5 ) begin
      act_regs_data_3_3_sva_8_25 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_3_3_sva_dfm_2_25_22_rsp_0, or_dcpl_873);
      act_regs_data_3_3_sva_8_24_22 <= MUX_v_3_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_3_3_sva_dfm_2_25_22_rsp_1, or_dcpl_873);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_2_sva_8_25 <= 1'b0;
      act_regs_data_3_2_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2744_enex5 ) begin
      act_regs_data_3_2_sva_8_25 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_3_2_sva_dfm_2_25_22_rsp_0, or_dcpl_874);
      act_regs_data_3_2_sva_8_24_22 <= MUX_v_3_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_3_2_sva_dfm_2_25_22_rsp_1, or_dcpl_874);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_regs_data_3_1_sva_8_25 <= 1'b0;
      act_regs_data_3_1_sva_8_24_22 <= 3'b000;
    end
    else if ( act_regs_data_and_2747_enex5 ) begin
      act_regs_data_3_1_sva_8_25 <= MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[25]),
          act_regs_data_3_1_sva_dfm_2_25_22_rsp_0, or_dcpl_875);
      act_regs_data_3_1_sva_8_24_22 <= MUX_v_3_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[24:22]),
          act_regs_data_3_1_sva_dfm_2_25_22_rsp_1, or_dcpl_875);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_1_25 <= 1'b0;
      ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_1_24_22 <= 3'b000;
    end
    else if ( and_1881_tmp ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_1_25 <= ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_9_nl
          & (~ or_dcpl);
      ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_1_24_22 <= MUX_v_3_2_2(3'b000,
          ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_191_nl, not_8895_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_1_25 <= 1'b0;
      ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_1_24_22 <= 3'b000;
    end
    else if ( and_1883_tmp ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_1_25 <= ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_14_nl
          & (~ or_dcpl);
      ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_1_24_22 <= MUX_v_3_2_2(3'b000,
          ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_190_nl, not_8894_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_1_25 <= 1'b0;
      ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_1_24_22 <= 3'b000;
    end
    else if ( and_1885_tmp ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_1_25 <= ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_19_nl
          & (~ or_dcpl);
      ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_1_24_22 <= MUX_v_3_2_2(3'b000,
          ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_189_nl, not_8893_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_1_25 <= 1'b0;
      ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_1_24_22 <= 3'b000;
    end
    else if ( and_1887_tmp ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_1_25 <= ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_24_nl
          & (~ or_dcpl);
      ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_1_24_22 <= MUX_v_3_2_2(3'b000,
          ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_188_nl, not_8892_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_1_25 <= 1'b0;
      ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_1_24_22 <= 3'b000;
    end
    else if ( and_1889_tmp ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_1_25 <= ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_29_nl
          & (~ or_dcpl);
      ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_1_24_22 <= MUX_v_3_2_2(3'b000,
          ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_187_nl, not_8891_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_1_25 <= 1'b0;
      ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_1_24_22 <= 3'b000;
    end
    else if ( and_1891_tmp ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_1_25 <= ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_34_nl
          & (~ or_dcpl);
      ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_1_24_22 <= MUX_v_3_2_2(3'b000,
          ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_198_nl, not_8903_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_1_25 <= 1'b0;
      ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_1_24_22 <= 3'b000;
    end
    else if ( and_1893_tmp ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_1_25 <= ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_39_nl
          & (~ or_dcpl);
      ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_1_24_22 <= MUX_v_3_2_2(3'b000,
          ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_197_nl, not_8902_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_1_25 <= 1'b0;
      ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_1_24_22 <= 3'b000;
    end
    else if ( and_1895_tmp ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_1_25 <= ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_44_nl
          & (~ or_dcpl);
      ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_1_24_22 <= MUX_v_3_2_2(3'b000,
          ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_196_nl, not_8901_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_1_25 <= 1'b0;
      ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_1_24_22 <= 3'b000;
    end
    else if ( and_1897_tmp ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_1_25 <= ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_49_nl
          & (~ or_dcpl);
      ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_1_24_22 <= MUX_v_3_2_2(3'b000,
          ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_195_nl, not_8900_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_1_25 <= 1'b0;
      ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_1_24_22 <= 3'b000;
    end
    else if ( and_1899_tmp ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_1_25 <= ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_54_nl
          & (~ or_dcpl);
      ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_1_24_22 <= MUX_v_3_2_2(3'b000,
          ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_194_nl, not_8899_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_1_25 <= 1'b0;
      ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_1_24_22 <= 3'b000;
    end
    else if ( and_1901_tmp ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_1_25 <= ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_59_nl
          & (~ or_dcpl);
      ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_1_24_22 <= MUX_v_3_2_2(3'b000,
          ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_193_nl, not_8898_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_1_25 <= 1'b0;
      ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_1_24_22 <= 3'b000;
    end
    else if ( and_1903_tmp ) begin
      ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_1_25 <= ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_64_nl
          & (~ or_dcpl);
      ActUnit_PushOutput_if_output_port_reg_data_data_8_sva_1_24_22 <= MUX_v_3_2_2(3'b000,
          ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_192_nl, not_8897_nl);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_13_ftd_2_3 <= 1'b0;
      reg_act_regs_data_0_13_ftd_2_2_0 <= 3'b000;
    end
    else if ( act_regs_data_and_2750_enex5 ) begin
      reg_act_regs_data_0_13_ftd_2_3 <= MUX1HOT_s_1_3_2(act_regs_data_0_13_sva_dfm_2_25_22_rsp_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_1_25, act_regs_data_0_13_sva_8_25,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      reg_act_regs_data_0_13_ftd_2_2_0 <= MUX1HOT_v_3_3_2(act_regs_data_0_13_sva_dfm_2_25_22_rsp_1,
          ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_1_24_22, act_regs_data_0_13_sva_8_24_22,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_12_ftd_2_3 <= 1'b0;
      reg_act_regs_data_0_12_ftd_2_2_0 <= 3'b000;
    end
    else if ( act_regs_data_and_2753_enex5 ) begin
      reg_act_regs_data_0_12_ftd_2_3 <= MUX1HOT_s_1_3_2(act_regs_data_0_12_sva_dfm_2_25_22_rsp_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_1_25, act_regs_data_0_12_sva_8_25,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      reg_act_regs_data_0_12_ftd_2_2_0 <= MUX1HOT_v_3_3_2(act_regs_data_0_12_sva_dfm_2_25_22_rsp_1,
          ActUnit_PushOutput_if_output_port_reg_data_data_12_sva_1_24_22, act_regs_data_0_12_sva_8_24_22,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_11_ftd_2_3 <= 1'b0;
      reg_act_regs_data_0_11_ftd_2_2_0 <= 3'b000;
    end
    else if ( act_regs_data_and_2756_enex5 ) begin
      reg_act_regs_data_0_11_ftd_2_3 <= MUX1HOT_s_1_3_2(act_regs_data_0_11_sva_dfm_2_25_22_rsp_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_1_25, act_regs_data_0_11_sva_8_25,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      reg_act_regs_data_0_11_ftd_2_2_0 <= MUX1HOT_v_3_3_2(act_regs_data_0_11_sva_dfm_2_25_22_rsp_1,
          ActUnit_PushOutput_if_output_port_reg_data_data_11_sva_1_24_22, act_regs_data_0_11_sva_8_24_22,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_10_ftd_2_3 <= 1'b0;
      reg_act_regs_data_0_10_ftd_2_2_0 <= 3'b000;
    end
    else if ( act_regs_data_and_2759_enex5 ) begin
      reg_act_regs_data_0_10_ftd_2_3 <= MUX1HOT_s_1_3_2(act_regs_data_0_10_sva_dfm_2_25_22_rsp_0,
          ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_1_25, act_regs_data_0_10_sva_8_25,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      reg_act_regs_data_0_10_ftd_2_2_0 <= MUX1HOT_v_3_3_2(act_regs_data_0_10_sva_dfm_2_25_22_rsp_1,
          ActUnit_PushOutput_if_output_port_reg_data_data_10_sva_1_24_22, act_regs_data_0_10_sva_8_24_22,
          {while_nand_ssc_1 , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_1_ftd_2_3 <= 1'b0;
      reg_act_regs_data_0_1_ftd_2_2_0 <= 3'b000;
    end
    else if ( act_regs_data_and_2762_enex5 ) begin
      reg_act_regs_data_0_1_ftd_2_3 <= MUX1HOT_s_1_3_2(act_regs_data_0_1_sva_dfm_2_25_22_rsp_0,
          rva_out_reg_data_39_32_sva_dfm_6_3, act_regs_data_0_1_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      reg_act_regs_data_0_1_ftd_2_2_0 <= MUX1HOT_v_3_3_2(act_regs_data_0_1_sva_dfm_2_25_22_rsp_1,
          rva_out_reg_data_39_32_sva_dfm_6_2_0, act_regs_data_0_1_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_regs_data_0_0_ftd_2_3 <= 1'b0;
      reg_act_regs_data_0_0_ftd_2_2_0 <= 3'b000;
    end
    else if ( act_regs_data_and_2765_enex5 ) begin
      reg_act_regs_data_0_0_ftd_2_3 <= MUX1HOT_s_1_3_2(act_regs_data_0_0_sva_dfm_2_25_22_rsp_0,
          rva_out_reg_data_29_24_sva_dfm_6_3, act_regs_data_0_0_sva_8_25, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
      reg_act_regs_data_0_0_ftd_2_2_0 <= MUX1HOT_v_3_3_2(act_regs_data_0_0_sva_dfm_2_25_22_rsp_1,
          rva_out_reg_data_29_24_sva_dfm_6_2_0, act_regs_data_0_0_sva_8_24_22, {while_nand_ssc_1
          , ActUnit_RunLoad_and_ssc_1 , ActUnit_RunLoad_and_1_ssc_1});
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_ActUnit_RunInst_case_14_nv_scvector_cctor_data_0_1_ftd_rsp_0 <= 1'b0;
      reg_ActUnit_RunInst_case_14_nv_scvector_cctor_data_0_1_ftd_rsp_1 <= 3'b000;
    end
    else if ( ActUnit_RunInst_switch_lp_and_816_enex5 ) begin
      reg_ActUnit_RunInst_case_14_nv_scvector_cctor_data_0_1_ftd_rsp_0 <= nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
      reg_ActUnit_RunInst_case_14_nv_scvector_cctor_data_0_1_ftd_rsp_1 <= nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_2_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          <= 1'b0;
      reg_nv_scvector_cctor_nv_scvector_5_for_2_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          <= 3'b000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_2_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          <= nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
      reg_nv_scvector_cctor_nv_scvector_5_for_2_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          <= nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          <= 1'b0;
      reg_nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          <= 3'b000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_17_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          <= nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
      reg_nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          <= nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          <= 1'b0;
      reg_nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          <= 3'b000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_20_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          <= nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
      reg_nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          <= nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          <= 1'b0;
      reg_nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          <= 3'b000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_23_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          <= nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
      reg_nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          <= nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          <= 1'b0;
      reg_nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          <= 3'b000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_26_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          <= nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
      reg_nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          <= nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          <= 1'b0;
      reg_nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          <= 3'b000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_29_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          <= nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
      reg_nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          <= nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          <= 1'b0;
      reg_nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          <= 3'b000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_32_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          <= nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
      reg_nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          <= nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          <= 1'b0;
      reg_nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          <= 3'b000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_35_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          <= nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
      reg_nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          <= nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          <= 1'b0;
      reg_nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          <= 3'b000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_38_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          <= nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
      reg_nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          <= nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          <= 1'b0;
      reg_nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          <= 3'b000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_41_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          <= nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
      reg_nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          <= nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          <= 1'b0;
      reg_nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          <= 3'b000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_44_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          <= nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
      reg_nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          <= nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          <= 1'b0;
      reg_nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          <= 3'b000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_47_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          <= nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
      reg_nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          <= nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          <= 1'b0;
      reg_nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          <= 3'b000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_50_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          <= nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
      reg_nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          <= nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          <= 1'b0;
      reg_nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          <= 3'b000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_53_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          <= nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
      reg_nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          <= nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          <= 1'b0;
      reg_nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          <= 3'b000;
    end
    else if ( nv_scvector_cctor_nv_scvector_5_for_and_56_enex5 ) begin
      reg_nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
          <= nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_3;
      reg_nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1
          <= nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_2_itm_2_0;
    end
  end
  assign ActUnit_DecodeAxiRead_else_mux_3_nl = MUX_s_1_2_2(ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0,
      ActUnit_DecodeAxiWrite_else_unequal_tmp, or_dcpl_469);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_7_nl = (~ ActUnit_DecodeAxiRead_else_mux_3_nl)
      & ActUnit_DecodeAxiRead_unequal_tmp_1 & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & rva_in_PopNB_mioi_return_rsc_z_mxwt;
  assign and_1122_nl = and_dcpl_1077 & (fsm_output[3]) & while_asn_262_itm;
  assign while_else_1_while_else_1_nand_1_nl = ~(act_config_InstIncr_if_act_config_InstIncr_if_if_nor_tmp
      & act_config_InstIncr_act_config_InstIncr_if_and_svs_1 & is_incr_lpi_1_dfm_1);
  assign Silu_for_else_Silu_for_else_mux1h_2_nl = MUX1HOT_v_5_3_2((signext_5_1(Silu_for_y_3_sva_1_22_0_1[22])),
      (signext_5_1(Silu_for_3_else_else_if_acc_itm[1])), reg_nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26,
      {(~ Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_4_ssc_1 , Silu_for_else_else_else_and_5_ssc_1});
  assign Silu_for_else_nor_5_nl = ~(Silu_for_else_and_34_ssc_1 | Silu_for_else_else_else_and_4_ssc_1);
  assign Silu_for_Silu_for_and_22_nl = Silu_for_else_Silu_for_else_mux1h_2_nl & (signext_5_1(Silu_for_else_nor_5_nl))
      & ({{4{Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs}},
      Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs});
  assign mux1h_1_nl = MUX1HOT_v_5_3_2(Silu_for_Silu_for_and_22_nl, ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_30_26_2,
      act_regs_data_0_1_sva_dfm_2_30_26, {and_dcpl_1112 , and_dcpl_1393 , and_1720_cse});
  assign not_2610_nl = ~ or_dcpl_1012;
  assign and_1716_nl = MUX_v_5_2_2(5'b00000, mux1h_1_nl, not_2610_nl);
  assign act_config_InstIncr_if_not_9_nl = ~ act_config_InstIncr_if_act_config_InstIncr_if_if_nor_mdf_sva;
  assign act_config_InstIncr_if_act_config_InstIncr_if_and_1_nl = MUX_v_4_2_2(4'b0000,
      (operator_8_false_acc_sdt[7:4]), act_config_InstIncr_if_not_9_nl);
  assign act_config_InstIncr_if_act_config_InstIncr_if_and_2_nl = (operator_8_false_acc_sdt[3])
      & (~ act_config_InstIncr_if_act_config_InstIncr_if_if_nor_mdf_sva);
  assign act_config_InstIncr_if_not_10_nl = ~ act_config_InstIncr_if_act_config_InstIncr_if_if_nor_mdf_sva;
  assign act_config_InstIncr_if_act_config_InstIncr_if_and_3_nl = MUX_v_3_2_2(3'b000,
      (operator_8_false_acc_sdt[2:0]), act_config_InstIncr_if_not_10_nl);
  assign nl_operator_5_false_acc_nl = act_config_inst_counter_sva_dfm_3 + 5'b00001;
  assign operator_5_false_acc_nl = nl_operator_5_false_acc_nl[4:0];
  assign act_config_InstIncr_if_not_7_nl = ~ act_config_InstIncr_act_config_InstIncr_if_and_svs_1;
  assign act_config_InstIncr_act_config_InstIncr_and_1_nl = MUX_v_5_2_2(5'b00000,
      operator_5_false_acc_nl, act_config_InstIncr_if_not_7_nl);
  assign nl_Silu_for_1_else_else_if_acc_itm  = ({reg_ActUnit_RunInst_case_14_nv_scvector_cctor_data_0_1_ftd_rsp_0
      , (reg_ActUnit_RunInst_case_14_nv_scvector_cctor_data_0_1_ftd_rsp_1[2])}) +
      2'b01;
  assign nl_Silu_for_2_else_else_if_acc_itm  = ({reg_nv_scvector_cctor_nv_scvector_5_for_2_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , (reg_nv_scvector_cctor_nv_scvector_5_for_2_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1[2])})
      + 2'b01;
  assign nl_Silu_for_3_else_else_if_acc_itm  = ({reg_nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , (reg_nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1[2])})
      + 2'b01;
  assign nl_Silu_for_4_else_else_if_acc_itm  = ({reg_nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , (reg_nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1[2])})
      + 2'b01;
  assign nl_Silu_for_5_else_else_if_acc_itm  = ({reg_nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , (reg_nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1[2])})
      + 2'b01;
  assign nl_Silu_for_6_else_else_if_acc_itm  = ({reg_nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , (reg_nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1[2])})
      + 2'b01;
  assign nl_Silu_for_7_else_else_if_acc_itm  = ({reg_nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , (reg_nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1[2])})
      + 2'b01;
  assign nl_Silu_for_8_else_else_if_acc_itm  = ({reg_nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , (reg_nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1[2])})
      + 2'b01;
  assign nl_Silu_for_9_else_else_if_acc_itm  = ({reg_nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , (reg_nv_scvector_cctor_nv_scvector_5_for_9_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1[2])})
      + 2'b01;
  assign nl_Silu_for_10_else_else_if_acc_itm  = ({reg_nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , (reg_nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1[2])})
      + 2'b01;
  assign nl_Silu_for_11_else_else_if_acc_itm  = ({reg_nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , (reg_nv_scvector_cctor_nv_scvector_5_for_11_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1[2])})
      + 2'b01;
  assign nl_Silu_for_12_else_else_if_acc_itm  = ({reg_nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , (reg_nv_scvector_cctor_nv_scvector_5_for_12_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1[2])})
      + 2'b01;
  assign nl_Silu_for_13_else_else_if_acc_itm  = ({reg_nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , (reg_nv_scvector_cctor_nv_scvector_5_for_13_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1[2])})
      + 2'b01;
  assign nl_Silu_for_14_else_else_if_acc_itm  = ({reg_nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , (reg_nv_scvector_cctor_nv_scvector_5_for_14_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1[2])})
      + 2'b01;
  assign nl_Silu_for_15_else_else_if_acc_itm  = ({reg_nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , (reg_nv_scvector_cctor_nv_scvector_5_for_15_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1[2])})
      + 2'b01;
  assign nl_Silu_for_16_else_else_if_acc_itm  = ({reg_nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , (reg_nv_scvector_cctor_nv_scvector_5_for_16_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1[2])})
      + 2'b01;
  assign and_1276_nl = nor_222_cse & and_dcpl_1233;
  assign nor_1408_nl = ~((act_config_inst_regs_0_sva_dfm_5[7:4]!=4'b0010));
  assign nor_1409_nl = ~((act_config_inst_regs_1_sva_dfm_5[7:4]!=4'b0010));
  assign mux_617_nl = MUX_s_1_2_2(nor_1408_nl, nor_1409_nl, act_config_inst_counter_sva[0]);
  assign nor_1410_nl = ~((act_config_inst_regs_2_sva_dfm_5[7:4]!=4'b0010));
  assign nor_1411_nl = ~((act_config_inst_regs_3_sva_dfm_5[7:4]!=4'b0010));
  assign mux_616_nl = MUX_s_1_2_2(nor_1410_nl, nor_1411_nl, act_config_inst_counter_sva[0]);
  assign mux_618_nl = MUX_s_1_2_2(mux_617_nl, mux_616_nl, act_config_inst_counter_sva[1]);
  assign nor_1412_nl = ~((act_config_inst_regs_4_sva_dfm_5[7:4]!=4'b0010));
  assign nor_1413_nl = ~((act_config_inst_regs_5_sva_dfm_5[7:4]!=4'b0010));
  assign mux_614_nl = MUX_s_1_2_2(nor_1412_nl, nor_1413_nl, act_config_inst_counter_sva[0]);
  assign nor_1414_nl = ~((act_config_inst_regs_6_sva_dfm_5[7:4]!=4'b0010));
  assign nor_1415_nl = ~((act_config_inst_regs_7_sva_dfm_5[7:4]!=4'b0010));
  assign mux_613_nl = MUX_s_1_2_2(nor_1414_nl, nor_1415_nl, act_config_inst_counter_sva[0]);
  assign mux_615_nl = MUX_s_1_2_2(mux_614_nl, mux_613_nl, act_config_inst_counter_sva[1]);
  assign mux_619_nl = MUX_s_1_2_2(mux_618_nl, mux_615_nl, act_config_inst_counter_sva[2]);
  assign nor_1416_nl = ~((act_config_inst_regs_8_sva_dfm_5[7:4]!=4'b0010));
  assign nor_1417_nl = ~((act_config_inst_regs_9_sva_dfm_5[7:4]!=4'b0010));
  assign mux_610_nl = MUX_s_1_2_2(nor_1416_nl, nor_1417_nl, act_config_inst_counter_sva[0]);
  assign nor_1418_nl = ~((act_config_inst_regs_10_sva_dfm_5[7:4]!=4'b0010));
  assign nor_1419_nl = ~((act_config_inst_regs_11_sva_dfm_5[7:4]!=4'b0010));
  assign mux_609_nl = MUX_s_1_2_2(nor_1418_nl, nor_1419_nl, act_config_inst_counter_sva[0]);
  assign mux_611_nl = MUX_s_1_2_2(mux_610_nl, mux_609_nl, act_config_inst_counter_sva[1]);
  assign nor_1420_nl = ~((act_config_inst_regs_12_sva_dfm_5[7:4]!=4'b0010));
  assign nor_1421_nl = ~((act_config_inst_regs_13_sva_dfm_5[7:4]!=4'b0010));
  assign mux_607_nl = MUX_s_1_2_2(nor_1420_nl, nor_1421_nl, act_config_inst_counter_sva[0]);
  assign nor_1422_nl = ~((act_config_inst_regs_14_sva_dfm_5[7:4]!=4'b0010));
  assign nor_1423_nl = ~((act_config_inst_regs_15_sva_dfm_5[7:4]!=4'b0010));
  assign mux_606_nl = MUX_s_1_2_2(nor_1422_nl, nor_1423_nl, act_config_inst_counter_sva[0]);
  assign mux_608_nl = MUX_s_1_2_2(mux_607_nl, mux_606_nl, act_config_inst_counter_sva[1]);
  assign mux_612_nl = MUX_s_1_2_2(mux_611_nl, mux_608_nl, act_config_inst_counter_sva[2]);
  assign mux_620_nl = MUX_s_1_2_2(mux_619_nl, mux_612_nl, act_config_inst_counter_sva[3]);
  assign nor_1424_nl = ~((act_config_inst_regs_16_sva_dfm_6[7:4]!=4'b0010));
  assign nor_1425_nl = ~((act_config_inst_regs_17_sva_dfm_6[7:4]!=4'b0010));
  assign mux_602_nl = MUX_s_1_2_2(nor_1424_nl, nor_1425_nl, act_config_inst_counter_sva[0]);
  assign nor_1426_nl = ~((act_config_inst_regs_18_sva_dfm_6[7:4]!=4'b0010));
  assign nor_1427_nl = ~((act_config_inst_regs_19_sva_dfm_6[7:4]!=4'b0010));
  assign mux_601_nl = MUX_s_1_2_2(nor_1426_nl, nor_1427_nl, act_config_inst_counter_sva[0]);
  assign mux_603_nl = MUX_s_1_2_2(mux_602_nl, mux_601_nl, act_config_inst_counter_sva[1]);
  assign nor_1428_nl = ~((act_config_inst_regs_20_sva_dfm_6[7:4]!=4'b0010));
  assign nor_1429_nl = ~((act_config_inst_regs_21_sva_dfm_6[7:4]!=4'b0010));
  assign mux_599_nl = MUX_s_1_2_2(nor_1428_nl, nor_1429_nl, act_config_inst_counter_sva[0]);
  assign nor_1430_nl = ~((act_config_inst_regs_22_sva_dfm_6[7:4]!=4'b0010));
  assign nor_1431_nl = ~((act_config_inst_regs_23_sva_dfm_6[7:4]!=4'b0010));
  assign mux_598_nl = MUX_s_1_2_2(nor_1430_nl, nor_1431_nl, act_config_inst_counter_sva[0]);
  assign mux_600_nl = MUX_s_1_2_2(mux_599_nl, mux_598_nl, act_config_inst_counter_sva[1]);
  assign mux_604_nl = MUX_s_1_2_2(mux_603_nl, mux_600_nl, act_config_inst_counter_sva[2]);
  assign nor_1432_nl = ~((act_config_inst_regs_24_sva_dfm_6[7:4]!=4'b0010));
  assign nor_1433_nl = ~((act_config_inst_regs_25_sva_dfm_6[7:4]!=4'b0010));
  assign mux_595_nl = MUX_s_1_2_2(nor_1432_nl, nor_1433_nl, act_config_inst_counter_sva[0]);
  assign nor_1434_nl = ~((act_config_inst_regs_26_sva_dfm_6[7:4]!=4'b0010));
  assign nor_1435_nl = ~((act_config_inst_regs_27_sva_dfm_6[7:4]!=4'b0010));
  assign mux_594_nl = MUX_s_1_2_2(nor_1434_nl, nor_1435_nl, act_config_inst_counter_sva[0]);
  assign mux_596_nl = MUX_s_1_2_2(mux_595_nl, mux_594_nl, act_config_inst_counter_sva[1]);
  assign nor_1436_nl = ~((act_config_inst_regs_28_sva_dfm_6[7:4]!=4'b0010));
  assign nor_1437_nl = ~((act_config_inst_regs_29_sva_dfm_6[7:4]!=4'b0010));
  assign mux_592_nl = MUX_s_1_2_2(nor_1436_nl, nor_1437_nl, act_config_inst_counter_sva[0]);
  assign nor_1438_nl = ~((act_config_inst_regs_30_sva_dfm_6[7:4]!=4'b0010));
  assign nor_1439_nl = ~((act_config_inst_regs_31_sva_dfm_6[7:4]!=4'b0010));
  assign mux_591_nl = MUX_s_1_2_2(nor_1438_nl, nor_1439_nl, act_config_inst_counter_sva[0]);
  assign mux_593_nl = MUX_s_1_2_2(mux_592_nl, mux_591_nl, act_config_inst_counter_sva[1]);
  assign mux_597_nl = MUX_s_1_2_2(mux_596_nl, mux_593_nl, act_config_inst_counter_sva[2]);
  assign mux_605_nl = MUX_s_1_2_2(mux_604_nl, mux_597_nl, act_config_inst_counter_sva[3]);
  assign mux_621_nl = MUX_s_1_2_2(mux_620_nl, mux_605_nl, act_config_inst_counter_sva[4]);
  assign and_2331_nl = is_start_sva & mux_621_nl;
  assign nor_1440_nl = ~(is_start_sva | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11:9]!=3'b100)
      | (~(rva_in_PopNB_mioi_return_rsc_z_mxwt & rva_in_PopNB_mioi_data_rw_rsc_z_mxwt
      & (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[8]))));
  assign mux_622_nl = MUX_s_1_2_2(and_2331_nl, nor_1440_nl, fsm_output[1]);
  assign Silu_for_else_Silu_for_else_mux1h_1_nl = MUX1HOT_v_5_3_2((signext_5_1(Silu_for_y_2_sva_1_22_0_1[22])),
      (signext_5_1(Silu_for_2_else_else_if_acc_itm[1])), reg_nv_scvector_cctor_nv_scvector_5_for_2_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26,
      {(~ Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_2_ssc_1 , Silu_for_else_else_else_and_3_ssc_1});
  assign Silu_for_else_nor_3_nl = ~(Silu_for_else_and_33_ssc_1 | Silu_for_else_else_else_and_2_ssc_1);
  assign Silu_for_Silu_for_and_19_nl = Silu_for_else_Silu_for_else_mux1h_1_nl & (signext_5_1(Silu_for_else_nor_3_nl))
      & ({{4{Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs}},
      Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs});
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_121_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_0_0_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_291);
  assign ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_13_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      rva_out_reg_data_159_128_sva_dfm_3, ActUnit_DecodeAxiRead_unequal_tmp_1);
  assign ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_12_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      rva_out_reg_data_191_160_sva_dfm_3, ActUnit_DecodeAxiRead_unequal_tmp_1);
  assign ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_11_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      rva_out_reg_data_223_192_sva_dfm_3, ActUnit_DecodeAxiRead_unequal_tmp_1);
  assign ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_10_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      rva_out_reg_data_255_224_sva_dfm_3, ActUnit_DecodeAxiRead_unequal_tmp_1);
  assign ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_9_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      rva_out_reg_data_287_256_sva_dfm_3, ActUnit_DecodeAxiRead_unequal_tmp_1);
  assign ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_8_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      rva_out_reg_data_319_288_sva_dfm_3, ActUnit_DecodeAxiRead_unequal_tmp_1);
  assign ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_7_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      rva_out_reg_data_351_320_sva_dfm_3, ActUnit_DecodeAxiRead_unequal_tmp_1);
  assign ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_6_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      rva_out_reg_data_383_352_sva_dfm_3, ActUnit_DecodeAxiRead_unequal_tmp_1);
  assign ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_5_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      rva_out_reg_data_415_384_sva_dfm_3, ActUnit_DecodeAxiRead_unequal_tmp_1);
  assign ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_4_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      rva_out_reg_data_447_416_sva_dfm_3, ActUnit_DecodeAxiRead_unequal_tmp_1);
  assign ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_3_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      rva_out_reg_data_479_448_sva_dfm_3, ActUnit_DecodeAxiRead_unequal_tmp_1);
  assign ActUnit_DecodeAxiRead_ActUnit_DecodeAxiRead_and_nl = MUX_v_32_2_2(32'b00000000000000000000000000000000,
      rva_out_reg_data_511_480_sva_dfm_3, ActUnit_DecodeAxiRead_unequal_tmp_1);
  assign mux_572_nl = MUX_v_2_2_2((act_config_inst_regs_19_sva_dfm_6[7:6]), (act_config_inst_regs_3_sva_dfm_5[7:6]),
      and_dcpl_1257);
  assign not_2612_nl = ~ or_dcpl_1013;
  assign and_1721_nl = MUX_v_2_2_2(2'b00, mux_572_nl, not_2612_nl);
  assign mux_573_nl = MUX_v_8_2_2(act_config_inst_regs_28_sva_dfm_6, act_config_inst_regs_12_sva_dfm_5,
      and_dcpl_1257);
  assign not_2614_nl = ~ or_dcpl_1013;
  assign and_1723_nl = MUX_v_8_2_2(8'b00000000, mux_573_nl, not_2614_nl);
  assign mux_574_nl = MUX_v_8_2_2(act_config_inst_regs_29_sva_dfm_6, act_config_inst_regs_13_sva_dfm_5,
      and_dcpl_1257);
  assign not_2616_nl = ~ or_dcpl_1013;
  assign and_1725_nl = MUX_v_8_2_2(8'b00000000, mux_574_nl, not_2616_nl);
  assign mux_575_nl = MUX_v_8_2_2(act_config_inst_regs_30_sva_dfm_6, act_config_inst_regs_14_sva_dfm_5,
      and_dcpl_1257);
  assign not_2618_nl = ~ or_dcpl_1013;
  assign and_1727_nl = MUX_v_8_2_2(8'b00000000, mux_575_nl, not_2618_nl);
  assign mux_576_nl = MUX_v_8_2_2(act_config_inst_regs_31_sva_dfm_6, act_config_inst_regs_15_sva_dfm_5,
      and_dcpl_1257);
  assign not_2620_nl = ~ or_dcpl_1013;
  assign and_1729_nl = MUX_v_8_2_2(8'b00000000, mux_576_nl, not_2620_nl);
  assign mux_577_nl = MUX_v_8_2_2(act_config_inst_regs_18_sva_dfm_6, act_config_inst_regs_2_sva_dfm_5,
      and_dcpl_1257);
  assign not_2622_nl = ~ or_dcpl_1013;
  assign and_1731_nl = MUX_v_8_2_2(8'b00000000, mux_577_nl, not_2622_nl);
  assign mux_578_nl = MUX_v_8_2_2(act_config_inst_regs_21_sva_dfm_6, act_config_inst_regs_5_sva_dfm_5,
      and_dcpl_1257);
  assign not_2624_nl = ~ or_dcpl_1013;
  assign and_1733_nl = MUX_v_8_2_2(8'b00000000, mux_578_nl, not_2624_nl);
  assign mux_579_nl = MUX_v_8_2_2(act_config_inst_regs_23_sva_dfm_6, act_config_inst_regs_7_sva_dfm_5,
      and_dcpl_1257);
  assign not_2626_nl = ~ or_dcpl_1013;
  assign and_1735_nl = MUX_v_8_2_2(8'b00000000, mux_579_nl, not_2626_nl);
  assign mux_580_nl = MUX_v_8_2_2(act_config_inst_regs_25_sva_dfm_6, act_config_inst_regs_9_sva_dfm_5,
      and_dcpl_1257);
  assign not_2628_nl = ~ or_dcpl_1013;
  assign and_1737_nl = MUX_v_8_2_2(8'b00000000, mux_580_nl, not_2628_nl);
  assign mux_581_nl = MUX_v_8_2_2(act_config_inst_regs_26_sva_dfm_6, act_config_inst_regs_10_sva_dfm_5,
      and_dcpl_1257);
  assign not_2630_nl = ~ or_dcpl_1013;
  assign and_1739_nl = MUX_v_8_2_2(8'b00000000, mux_581_nl, not_2630_nl);
  assign mux_582_nl = MUX_v_8_2_2(act_config_inst_regs_27_sva_dfm_6, act_config_inst_regs_11_sva_dfm_5,
      and_dcpl_1257);
  assign not_2632_nl = ~ or_dcpl_1013;
  assign and_1741_nl = MUX_v_8_2_2(8'b00000000, mux_582_nl, not_2632_nl);
  assign mux_583_nl = MUX_v_7_2_2((act_config_inst_regs_17_sva_dfm_6[7:1]), (act_config_inst_regs_1_sva_dfm_5[7:1]),
      and_dcpl_1257);
  assign not_2634_nl = ~ or_dcpl_1013;
  assign and_1743_nl = MUX_v_7_2_2(7'b0000000, mux_583_nl, not_2634_nl);
  assign mux_584_nl = MUX_v_7_2_2((act_config_inst_regs_16_sva_dfm_6[7:1]), (act_config_inst_regs_0_sva_dfm_5[7:1]),
      and_dcpl_1257);
  assign not_2636_nl = ~ or_dcpl_1013;
  assign and_1745_nl = MUX_v_7_2_2(7'b0000000, mux_584_nl, not_2636_nl);
  assign mux_585_nl = MUX_v_3_2_2((act_config_inst_regs_22_sva_dfm_6[7:5]), (act_config_inst_regs_6_sva_dfm_5[7:5]),
      and_dcpl_1257);
  assign not_2638_nl = ~ or_dcpl_1013;
  assign and_1747_nl = MUX_v_3_2_2(3'b000, mux_585_nl, not_2638_nl);
  assign ActUnit_RunInst_switch_lp_mux_3_nl = MUX_s_1_2_2(ActUnit_RunInst_switch_lp_equal_tmp_1_mx0w0,
      ActUnit_RunInst_switch_lp_and_32_tmp, and_dcpl_849);
  assign ActUnit_RunInst_switch_lp_mux_4_nl = MUX_s_1_2_2(ActUnit_RunInst_switch_lp_equal_tmp_2_mx0w0,
      ActUnit_RunInst_switch_lp_equal_tmp_2, or_dcpl_823);
  assign ActUnit_RunInst_switch_lp_mux_6_nl = MUX_s_1_2_2(ActUnit_RunInst_switch_lp_equal_tmp_3_mx0w0,
      ActUnit_RunInst_switch_lp_equal_tmp_3, or_dcpl_823);
  assign ActUnit_RunInst_switch_lp_mux_8_nl = MUX_s_1_2_2(ActUnit_RunInst_switch_lp_equal_tmp_4_mx0w0,
      ActUnit_RunInst_switch_lp_equal_tmp_4, or_dcpl_823);
  assign ActUnit_RunInst_switch_lp_mux_10_nl = MUX_s_1_2_2(ActUnit_RunInst_switch_lp_equal_tmp_5_mx0w0,
      ActUnit_RunInst_switch_lp_equal_tmp_5, or_dcpl_823);
  assign ActUnit_RunInst_switch_lp_mux_12_nl = MUX_s_1_2_2(ActUnit_RunInst_switch_lp_equal_tmp_6_mx0w0,
      ActUnit_RunInst_switch_lp_equal_tmp_6, or_dcpl_823);
  assign ActUnit_RunInst_switch_lp_mux_14_nl = MUX_s_1_2_2(ActUnit_RunInst_switch_lp_equal_tmp_7_mx0w0,
      ActUnit_RunInst_switch_lp_equal_tmp_7, or_dcpl_823);
  assign ActUnit_RunInst_switch_lp_mux_16_nl = MUX_s_1_2_2(ActUnit_RunInst_switch_lp_equal_tmp_8_mx0w0,
      ActUnit_RunInst_switch_lp_equal_tmp_8, or_dcpl_823);
  assign mux_444_nl = MUX_s_1_2_2((fsm_output[1]), (~ and_2371_cse), fsm_output[2]);
  assign Tanh_for_or_2_nl = Tanh_for_and_79_ssc | Tanh_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
  assign Tanh_for_nor_1_nl = ~(Tanh_for_and_79_ssc | Tanh_for_16_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1);
  assign Tanh_for_or_3_nl = Tanh_for_and_77_ssc | Tanh_for_15_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
  assign Tanh_for_nor_2_nl = ~(Tanh_for_and_77_ssc | Tanh_for_15_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1);
  assign Tanh_for_or_4_nl = Tanh_for_and_75_ssc | Tanh_for_14_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
  assign Tanh_for_nor_3_nl = ~(Tanh_for_and_75_ssc | Tanh_for_14_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1);
  assign Tanh_for_or_5_nl = Tanh_for_and_73_ssc | Tanh_for_13_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
  assign Tanh_for_nor_4_nl = ~(Tanh_for_and_73_ssc | Tanh_for_13_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1);
  assign Tanh_for_or_6_nl = Tanh_for_and_71_ssc | Tanh_for_12_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
  assign Tanh_for_nor_5_nl = ~(Tanh_for_and_71_ssc | Tanh_for_12_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1);
  assign Tanh_for_or_7_nl = Tanh_for_and_69_ssc | Tanh_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
  assign Tanh_for_nor_6_nl = ~(Tanh_for_and_69_ssc | Tanh_for_11_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1);
  assign Tanh_for_or_8_nl = Tanh_for_and_67_ssc | Tanh_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
  assign Tanh_for_nor_7_nl = ~(Tanh_for_and_67_ssc | Tanh_for_10_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1);
  assign Tanh_for_or_9_nl = Tanh_for_and_65_ssc | Tanh_for_9_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
  assign Tanh_for_nor_8_nl = ~(Tanh_for_and_65_ssc | Tanh_for_9_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1);
  assign Tanh_for_or_10_nl = Tanh_for_and_63_ssc | Tanh_for_8_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
  assign Tanh_for_nor_9_nl = ~(Tanh_for_and_63_ssc | Tanh_for_8_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1);
  assign Tanh_for_or_11_nl = Tanh_for_and_61_ssc | Tanh_for_7_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
  assign Tanh_for_nor_10_nl = ~(Tanh_for_and_61_ssc | Tanh_for_7_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1);
  assign Tanh_for_or_12_nl = Tanh_for_and_59_ssc | Tanh_for_6_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
  assign Tanh_for_nor_11_nl = ~(Tanh_for_and_59_ssc | Tanh_for_6_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1);
  assign Tanh_for_or_13_nl = Tanh_for_and_57_ssc | Tanh_for_5_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
  assign Tanh_for_nor_12_nl = ~(Tanh_for_and_57_ssc | Tanh_for_5_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1);
  assign Tanh_for_or_14_nl = Tanh_for_and_55_ssc | Tanh_for_4_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
  assign Tanh_for_nor_13_nl = ~(Tanh_for_and_55_ssc | Tanh_for_4_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1);
  assign Tanh_for_or_15_nl = Tanh_for_and_53_ssc | Tanh_for_3_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
  assign Tanh_for_nor_14_nl = ~(Tanh_for_and_53_ssc | Tanh_for_3_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1);
  assign Tanh_for_or_16_nl = Tanh_for_and_51_ssc | Tanh_for_2_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
  assign Tanh_for_nor_15_nl = ~(Tanh_for_and_51_ssc | Tanh_for_2_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1);
  assign Tanh_for_or_17_nl = Tanh_for_and_49_ssc | Tanh_for_1_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1;
  assign Tanh_for_nor_16_nl = ~(Tanh_for_and_49_ssc | Tanh_for_1_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_8_svs_1);
  assign nv_scvector_cctor_nv_scvector_4_for_not_43_nl = ~ nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign nv_scvector_cctor_nv_scvector_4_for_not_59_nl = ~ nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign nv_scvector_cctor_nv_scvector_4_for_not_14_nl = ~ nv_scvector_cctor_nv_scvector_3_for_16_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign nv_scvector_cctor_nv_scvector_4_for_not_41_nl = ~ nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign nv_scvector_cctor_nv_scvector_4_for_not_58_nl = ~ nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign nv_scvector_cctor_nv_scvector_4_for_not_13_nl = ~ nv_scvector_cctor_nv_scvector_3_for_15_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign nv_scvector_cctor_nv_scvector_4_for_not_39_nl = ~ nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign nv_scvector_cctor_nv_scvector_4_for_not_57_nl = ~ nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign nv_scvector_cctor_nv_scvector_4_for_not_12_nl = ~ nv_scvector_cctor_nv_scvector_3_for_14_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign nv_scvector_cctor_nv_scvector_4_for_not_37_nl = ~ nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign nv_scvector_cctor_nv_scvector_4_for_not_56_nl = ~ nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign nv_scvector_cctor_nv_scvector_4_for_not_11_nl = ~ nv_scvector_cctor_nv_scvector_3_for_13_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign nv_scvector_cctor_nv_scvector_4_for_not_35_nl = ~ nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign nv_scvector_cctor_nv_scvector_4_for_not_55_nl = ~ nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign nv_scvector_cctor_nv_scvector_4_for_not_10_nl = ~ nv_scvector_cctor_nv_scvector_3_for_12_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign nv_scvector_cctor_nv_scvector_4_for_not_33_nl = ~ nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign nv_scvector_cctor_nv_scvector_4_for_not_54_nl = ~ nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign nv_scvector_cctor_nv_scvector_4_for_not_9_nl = ~ nv_scvector_cctor_nv_scvector_3_for_11_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign nv_scvector_cctor_nv_scvector_4_for_not_31_nl = ~ nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign nv_scvector_cctor_nv_scvector_4_for_not_53_nl = ~ nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign nv_scvector_cctor_nv_scvector_4_for_not_8_nl = ~ nv_scvector_cctor_nv_scvector_3_for_10_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign nv_scvector_cctor_nv_scvector_4_for_not_29_nl = ~ nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign nv_scvector_cctor_nv_scvector_4_for_not_52_nl = ~ nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign nv_scvector_cctor_nv_scvector_4_for_not_7_nl = ~ nv_scvector_cctor_nv_scvector_3_for_9_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign nv_scvector_cctor_nv_scvector_4_for_not_27_nl = ~ nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign nv_scvector_cctor_nv_scvector_4_for_not_51_nl = ~ nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign nv_scvector_cctor_nv_scvector_4_for_not_6_nl = ~ nv_scvector_cctor_nv_scvector_3_for_8_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign nv_scvector_cctor_nv_scvector_4_for_not_25_nl = ~ nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign nv_scvector_cctor_nv_scvector_4_for_not_50_nl = ~ nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign nv_scvector_cctor_nv_scvector_4_for_not_5_nl = ~ nv_scvector_cctor_nv_scvector_3_for_7_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign nv_scvector_cctor_nv_scvector_4_for_not_23_nl = ~ nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign nv_scvector_cctor_nv_scvector_4_for_not_49_nl = ~ nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign nv_scvector_cctor_nv_scvector_4_for_not_4_nl = ~ nv_scvector_cctor_nv_scvector_3_for_6_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign nv_scvector_cctor_nv_scvector_4_for_not_21_nl = ~ nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign nv_scvector_cctor_nv_scvector_4_for_not_48_nl = ~ nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign nv_scvector_cctor_nv_scvector_4_for_not_3_nl = ~ nv_scvector_cctor_nv_scvector_3_for_5_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign nv_scvector_cctor_nv_scvector_4_for_not_19_nl = ~ nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign nv_scvector_cctor_nv_scvector_4_for_not_47_nl = ~ nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign nv_scvector_cctor_nv_scvector_4_for_not_2_nl = ~ nv_scvector_cctor_nv_scvector_3_for_4_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign nv_scvector_cctor_nv_scvector_4_for_not_17_nl = ~ nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign nv_scvector_cctor_nv_scvector_4_for_not_46_nl = ~ nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign nv_scvector_cctor_nv_scvector_4_for_not_1_nl = ~ nv_scvector_cctor_nv_scvector_3_for_3_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign nv_scvector_cctor_nv_scvector_4_for_not_15_nl = ~ nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign nv_scvector_cctor_nv_scvector_4_for_not_45_nl = ~ nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign nv_scvector_cctor_nv_scvector_4_for_not_nl = ~ nv_scvector_cctor_nv_scvector_3_for_2_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign ActUnit_RunInst_switch_lp_not_10_nl = ~ nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign ActUnit_RunInst_switch_lp_not_12_nl = ~ nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign ActUnit_RunInst_switch_lp_not_1_nl = ~ nv_scvector_cctor_nv_scvector_3_for_1_nv_scvector_cctor_nv_scvector_3_for_nv_scvector_cctor_nv_scvector_3_for_mux_itm;
  assign ActUnit_RunInst_case_2_for_ActUnit_RunInst_case_2_for_and_1_nl = MUX_v_5_2_2(5'b00000,
      ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_30_26, ActUnit_RunInst_case_2_for_and_27_seb);
  assign ActUnit_RunInst_case_2_for_ActUnit_RunInst_case_2_for_and_2_nl = ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_25
      & ActUnit_RunInst_case_2_for_and_27_seb;
  assign ActUnit_RunInst_case_2_for_ActUnit_RunInst_case_2_for_and_4_nl = MUX_v_3_2_2(3'b000,
      ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_24_22, ActUnit_RunInst_case_2_for_and_27_seb);
  assign ActUnit_RunInst_case_2_for_ActUnit_RunInst_case_2_for_and_3_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_21_0, ActUnit_RunInst_case_2_for_and_27_seb);
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_nl = MUX_v_5_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_30_26,
      nv_scvector_cctor_nv_scvector_6_for_15_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26,
      act_write_data_data_and_96_cse);
  assign not_3249_nl = ~ and_dcpl_847;
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_1_nl = MUX_s_1_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_25,
      reg_nv_scvector_cctor_nv_scvector_6_for_15_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0,
      act_write_data_data_and_96_cse);
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_42_nl =
      MUX_v_3_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_24_22,
      reg_nv_scvector_cctor_nv_scvector_6_for_15_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1,
      act_write_data_data_and_96_cse);
  assign not_8967_nl = ~ and_dcpl_847;
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_2_nl = MUX_v_22_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_21_0,
      reg_nv_scvector_cctor_nv_scvector_6_for_15_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1,
      act_write_data_data_and_96_cse);
  assign not_2573_nl = ~ and_dcpl_847;
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_3_nl = MUX_v_5_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_30_26,
      nv_scvector_cctor_nv_scvector_6_for_10_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26,
      act_write_data_data_and_96_cse);
  assign not_3247_nl = ~ and_dcpl_847;
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_4_nl = MUX_s_1_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_25,
      reg_nv_scvector_cctor_nv_scvector_6_for_10_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0,
      act_write_data_data_and_96_cse);
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_43_nl =
      MUX_v_3_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_24_22,
      reg_nv_scvector_cctor_nv_scvector_6_for_10_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1,
      act_write_data_data_and_96_cse);
  assign not_8966_nl = ~ and_dcpl_847;
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_5_nl = MUX_v_22_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_21_0,
      reg_nv_scvector_cctor_nv_scvector_6_for_10_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1,
      act_write_data_data_and_96_cse);
  assign not_2571_nl = ~ and_dcpl_847;
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_6_nl = MUX_v_5_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_30_26,
      nv_scvector_cctor_nv_scvector_6_for_14_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26,
      act_write_data_data_and_96_cse);
  assign not_3245_nl = ~ and_dcpl_847;
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_7_nl = MUX_s_1_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_25,
      reg_nv_scvector_cctor_nv_scvector_6_for_14_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0,
      act_write_data_data_and_96_cse);
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_44_nl =
      MUX_v_3_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_24_22,
      reg_nv_scvector_cctor_nv_scvector_6_for_14_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1,
      act_write_data_data_and_96_cse);
  assign not_8965_nl = ~ and_dcpl_847;
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_8_nl = MUX_v_22_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_21_0,
      reg_nv_scvector_cctor_nv_scvector_6_for_14_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1,
      act_write_data_data_and_96_cse);
  assign not_2569_nl = ~ and_dcpl_847;
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_9_nl = MUX_v_5_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_30_26,
      nv_scvector_cctor_nv_scvector_6_for_2_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26,
      act_write_data_data_and_96_cse);
  assign not_3243_nl = ~ and_dcpl_847;
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_10_nl =
      MUX_s_1_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_25,
      reg_nv_scvector_cctor_nv_scvector_6_for_2_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0,
      act_write_data_data_and_96_cse);
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_45_nl =
      MUX_v_3_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_24_22,
      reg_nv_scvector_cctor_nv_scvector_6_for_2_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1,
      act_write_data_data_and_96_cse);
  assign not_8964_nl = ~ and_dcpl_847;
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_11_nl =
      MUX_v_22_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_21_0,
      reg_nv_scvector_cctor_nv_scvector_6_for_2_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1,
      act_write_data_data_and_96_cse);
  assign not_2567_nl = ~ and_dcpl_847;
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_12_nl =
      MUX_v_5_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_30_26,
      nv_scvector_cctor_nv_scvector_6_for_13_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26,
      act_write_data_data_and_96_cse);
  assign not_3241_nl = ~ and_dcpl_847;
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_13_nl =
      MUX_s_1_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_25,
      reg_nv_scvector_cctor_nv_scvector_6_for_13_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0,
      act_write_data_data_and_96_cse);
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_46_nl =
      MUX_v_3_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_24_22,
      reg_nv_scvector_cctor_nv_scvector_6_for_13_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1,
      act_write_data_data_and_96_cse);
  assign not_8963_nl = ~ and_dcpl_847;
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_14_nl =
      MUX_v_22_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_21_0,
      reg_nv_scvector_cctor_nv_scvector_6_for_13_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1,
      act_write_data_data_and_96_cse);
  assign not_2565_nl = ~ and_dcpl_847;
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_15_nl =
      MUX_v_5_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_30_26,
      nv_scvector_cctor_nv_scvector_6_for_3_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26,
      act_write_data_data_and_96_cse);
  assign not_3239_nl = ~ and_dcpl_847;
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_16_nl =
      MUX_s_1_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_25,
      reg_nv_scvector_cctor_nv_scvector_6_for_3_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0,
      act_write_data_data_and_96_cse);
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_47_nl =
      MUX_v_3_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_24_22,
      reg_nv_scvector_cctor_nv_scvector_6_for_3_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1,
      act_write_data_data_and_96_cse);
  assign not_8962_nl = ~ and_dcpl_847;
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_17_nl =
      MUX_v_22_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_21_0,
      reg_nv_scvector_cctor_nv_scvector_6_for_3_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1,
      act_write_data_data_and_96_cse);
  assign not_2563_nl = ~ and_dcpl_847;
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_18_nl =
      MUX_v_5_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_30_26,
      nv_scvector_cctor_nv_scvector_6_for_12_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26,
      act_write_data_data_and_96_cse);
  assign not_3237_nl = ~ and_dcpl_847;
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_19_nl =
      MUX_s_1_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_25,
      reg_nv_scvector_cctor_nv_scvector_6_for_12_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0,
      act_write_data_data_and_96_cse);
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_48_nl =
      MUX_v_3_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_24_22,
      reg_nv_scvector_cctor_nv_scvector_6_for_12_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1,
      act_write_data_data_and_96_cse);
  assign not_8961_nl = ~ and_dcpl_847;
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_20_nl =
      MUX_v_22_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_21_0,
      reg_nv_scvector_cctor_nv_scvector_6_for_12_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1,
      act_write_data_data_and_96_cse);
  assign not_2561_nl = ~ and_dcpl_847;
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_21_nl =
      MUX_v_5_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_30_26,
      nv_scvector_cctor_nv_scvector_6_for_4_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26,
      act_write_data_data_and_96_cse);
  assign not_3235_nl = ~ and_dcpl_847;
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_22_nl =
      MUX_s_1_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_25,
      reg_nv_scvector_cctor_nv_scvector_6_for_4_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0,
      act_write_data_data_and_96_cse);
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_49_nl =
      MUX_v_3_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_24_22,
      reg_nv_scvector_cctor_nv_scvector_6_for_4_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1,
      act_write_data_data_and_96_cse);
  assign not_8960_nl = ~ and_dcpl_847;
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_23_nl =
      MUX_v_22_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_21_0,
      reg_nv_scvector_cctor_nv_scvector_6_for_4_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1,
      act_write_data_data_and_96_cse);
  assign not_2559_nl = ~ and_dcpl_847;
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_24_nl =
      MUX_v_5_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_30_26,
      nv_scvector_cctor_nv_scvector_6_for_11_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26,
      act_write_data_data_and_96_cse);
  assign not_3233_nl = ~ and_dcpl_847;
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_25_nl =
      MUX_s_1_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_25,
      reg_nv_scvector_cctor_nv_scvector_6_for_11_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0,
      act_write_data_data_and_96_cse);
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_50_nl =
      MUX_v_3_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_24_22,
      reg_nv_scvector_cctor_nv_scvector_6_for_11_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1,
      act_write_data_data_and_96_cse);
  assign not_8959_nl = ~ and_dcpl_847;
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_26_nl =
      MUX_v_22_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_21_0,
      reg_nv_scvector_cctor_nv_scvector_6_for_11_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1,
      act_write_data_data_and_96_cse);
  assign not_2557_nl = ~ and_dcpl_847;
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_27_nl =
      MUX_v_5_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_30_26,
      nv_scvector_cctor_nv_scvector_6_for_5_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26,
      act_write_data_data_and_96_cse);
  assign not_3231_nl = ~ and_dcpl_847;
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_28_nl =
      MUX_s_1_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_25,
      reg_nv_scvector_cctor_nv_scvector_6_for_5_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0,
      act_write_data_data_and_96_cse);
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_51_nl =
      MUX_v_3_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_24_22,
      reg_nv_scvector_cctor_nv_scvector_6_for_5_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1,
      act_write_data_data_and_96_cse);
  assign not_8958_nl = ~ and_dcpl_847;
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_29_nl =
      MUX_v_22_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_21_0,
      reg_nv_scvector_cctor_nv_scvector_6_for_5_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1,
      act_write_data_data_and_96_cse);
  assign not_2555_nl = ~ and_dcpl_847;
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_30_nl =
      MUX_v_5_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_30_26,
      nv_scvector_cctor_nv_scvector_6_for_9_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26,
      act_write_data_data_and_96_cse);
  assign not_3229_nl = ~ and_dcpl_847;
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_31_nl =
      MUX_s_1_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_25,
      reg_nv_scvector_cctor_nv_scvector_6_for_9_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0,
      act_write_data_data_and_96_cse);
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_52_nl =
      MUX_v_3_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_24_22,
      reg_nv_scvector_cctor_nv_scvector_6_for_9_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1,
      act_write_data_data_and_96_cse);
  assign not_8957_nl = ~ and_dcpl_847;
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_32_nl =
      MUX_v_22_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_21_0,
      reg_nv_scvector_cctor_nv_scvector_6_for_9_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1,
      act_write_data_data_and_96_cse);
  assign not_2553_nl = ~ and_dcpl_847;
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_33_nl =
      MUX_v_5_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_30_26,
      nv_scvector_cctor_nv_scvector_6_for_6_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26,
      act_write_data_data_and_96_cse);
  assign not_3227_nl = ~ and_dcpl_847;
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_34_nl =
      MUX_s_1_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_25,
      reg_nv_scvector_cctor_nv_scvector_6_for_6_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0,
      act_write_data_data_and_96_cse);
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_53_nl =
      MUX_v_3_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_24_22,
      reg_nv_scvector_cctor_nv_scvector_6_for_6_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1,
      act_write_data_data_and_96_cse);
  assign not_8956_nl = ~ and_dcpl_847;
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_35_nl =
      MUX_v_22_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_21_0,
      reg_nv_scvector_cctor_nv_scvector_6_for_6_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1,
      act_write_data_data_and_96_cse);
  assign not_2551_nl = ~ and_dcpl_847;
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_36_nl =
      MUX_v_5_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_30_26,
      nv_scvector_cctor_nv_scvector_6_for_8_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26,
      act_write_data_data_and_96_cse);
  assign not_3225_nl = ~ and_dcpl_847;
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_37_nl =
      MUX_s_1_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_25,
      reg_nv_scvector_cctor_nv_scvector_6_for_8_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0,
      act_write_data_data_and_96_cse);
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_54_nl =
      MUX_v_3_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_24_22,
      reg_nv_scvector_cctor_nv_scvector_6_for_8_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1,
      act_write_data_data_and_96_cse);
  assign not_8955_nl = ~ and_dcpl_847;
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_38_nl =
      MUX_v_22_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_21_0,
      reg_nv_scvector_cctor_nv_scvector_6_for_8_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1,
      act_write_data_data_and_96_cse);
  assign not_2549_nl = ~ and_dcpl_847;
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_39_nl =
      MUX_v_5_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_30_26,
      nv_scvector_cctor_nv_scvector_6_for_7_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_sva_30_26,
      act_write_data_data_and_96_cse);
  assign not_3223_nl = ~ and_dcpl_847;
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_40_nl =
      MUX_s_1_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_25,
      reg_nv_scvector_cctor_nv_scvector_6_for_7_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_0,
      act_write_data_data_and_96_cse);
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_55_nl =
      MUX_v_3_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_24_22,
      reg_nv_scvector_cctor_nv_scvector_6_for_7_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_rsp_1,
      act_write_data_data_and_96_cse);
  assign not_8954_nl = ~ and_dcpl_847;
  assign act_write_data_data_act_write_data_data_act_write_data_data_mux_41_nl =
      MUX_v_22_2_2(ActUnit_RunInst_case_2_for_slc_act_regs_data_32_31_0_2_ctmp_sva_1_21_0,
      reg_nv_scvector_cctor_nv_scvector_6_for_7_nv_scvector_cctor_nv_scvector_6_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1,
      act_write_data_data_and_96_cse);
  assign not_2547_nl = ~ and_dcpl_847;
  assign ActUnit_CheckStart_if_ActUnit_CheckStart_if_and_nl = ActUnit_CheckStart_start_reg_sva
      & act_config_is_valid_sva & ActUnit_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva;
  assign ActUnit_RunInst_switch_lp_or_1_nl = ActUnit_CheckStart_Connections_InBlocking_bool_Connections_SYN_PORT_PopNB_return_sva_mx0c4
      | and_dcpl_1246;
  assign mux_445_nl = MUX_s_1_2_2(and_dcpl_848, or_tmp_484, fsm_output[2]);
  assign ActUnit_PushOutput_if_for_i_not_nl = ~ ActUnit_PushOutput_if_for_i_4_0_sva_3_0_mx0c0;
  assign Silu_for_else_Silu_for_else_mux1h_nl = MUX1HOT_v_5_3_2((signext_5_1(Silu_for_y_1_sva_1_22_0_1[22])),
      (signext_5_1(Silu_for_1_else_else_if_acc_itm[1])), reg_ActUnit_RunInst_case_14_nv_scvector_cctor_data_0_ftd_1_30_26,
      {(~ Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_ssc_1 , Silu_for_else_else_else_and_1_ssc_1});
  assign Silu_for_else_nor_1_nl = ~(Silu_for_else_and_32_ssc_1 | Silu_for_else_else_else_and_ssc_1);
  assign Silu_for_Silu_for_and_16_nl = Silu_for_else_Silu_for_else_mux1h_nl & (signext_5_1(Silu_for_else_nor_1_nl))
      & ({{4{Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs}},
      Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs});
  assign ActUnit_DecodeAxiRead_else_mux_1_nl = MUX_s_1_2_2(ActUnit_DecodeAxiRead_else_unequal_tmp_mx0w0,
      ActUnit_DecodeAxiRead_else_unequal_tmp, or_dcpl_466);
  assign ActUnit_DecodeAxi_ActUnit_DecodeAxi_and_5_nl = (~ ActUnit_DecodeAxiRead_else_mux_1_nl)
      & ActUnit_DecodeAxiRead_unequal_tmp_1 & (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt)
      & rva_in_PopNB_mioi_return_rsc_z_mxwt;
  assign act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_24_nl
      = act_config_inst_regs_16_sva_0 & act_config_ActConfigRead_else_else_not_21;
  assign act_config_ActConfigRead_else_mux_19_nl = MUX_s_1_2_2(act_config_inst_regs_0_sva_0,
      act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_24_nl,
      act_config_ActConfigRead_else_unequal_tmp_1);
  assign act_config_ActConfigRead_mux_19_nl = MUX_s_1_2_2(act_config_is_valid_sva,
      act_config_ActConfigRead_else_mux_19_nl, act_config_ActConfigRead_unequal_tmp_1);
  assign ActUnit_DecodeAxiRead_mux_33_nl = MUX_s_1_2_2(act_config_ActConfigRead_mux_19_nl,
      ActUnit_PushOutput_if_for_and_stg_2_7_sva, ActUnit_DecodeAxiRead_unequal_tmp_1);
  assign ActUnit_DecodeAxi_if_mux_91_nl = MUX_s_1_2_2(ActUnit_DecodeAxiRead_mux_33_nl,
      ActUnit_PushOutput_if_for_and_stg_2_7_sva, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt);
  assign ActUnit_DecodeAxi_mux_93_nl = MUX_s_1_2_2(ActUnit_PushOutput_if_for_and_stg_2_7_sva,
      ActUnit_DecodeAxi_if_mux_91_nl, rva_in_PopNB_mioi_return_rsc_z_mxwt);
  assign act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_18_nl
      = act_config_inst_regs_17_sva_0 & act_config_ActConfigRead_else_else_not_21;
  assign act_config_ActConfigRead_else_mux_17_nl = MUX_s_1_2_2(act_config_inst_regs_1_sva_0,
      act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_18_nl,
      act_config_ActConfigRead_else_unequal_tmp_1);
  assign act_config_ActConfigRead_mux_17_nl = MUX_s_1_2_2(act_config_is_zero_first_sva,
      act_config_ActConfigRead_else_mux_17_nl, act_config_ActConfigRead_unequal_tmp_1);
  assign ActUnit_DecodeAxiRead_mux_31_nl = MUX_s_1_2_2(act_config_ActConfigRead_mux_17_nl,
      Gelu_for_and_2_cse_sva, ActUnit_DecodeAxiRead_unequal_tmp_1);
  assign ActUnit_DecodeAxi_if_mux_89_nl = MUX_s_1_2_2(ActUnit_DecodeAxiRead_mux_31_nl,
      Gelu_for_and_2_cse_sva, rva_in_PopNB_mioi_data_rw_rsc_z_mxwt);
  assign ActUnit_DecodeAxi_mux_94_nl = MUX_s_1_2_2(Gelu_for_and_2_cse_sva, ActUnit_DecodeAxi_if_mux_89_nl,
      rva_in_PopNB_mioi_return_rsc_z_mxwt);
  assign act_config_ActConfigRead_else_else_act_config_ActConfigRead_else_else_and_22_nl
      = MUX_v_5_2_2(5'b00000, (act_config_inst_regs_22_sva_dfm_6[4:0]), act_config_ActConfigRead_else_else_not_21);
  assign act_config_ActConfigWrite_mux_1_nl = MUX_s_1_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[8]),
      act_config_is_zero_first_sva, act_config_ActConfigRead_unequal_tmp_1);
  assign ActUnit_DecodeAxiWrite_mux_4_nl = MUX_s_1_2_2(act_config_ActConfigWrite_mux_1_nl,
      act_config_is_zero_first_sva, ActUnit_DecodeAxiRead_unequal_tmp_1);
  assign mux_1495_nl = MUX_v_22_2_2(ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_21_0_mx0w1,
      act_regs_data_0_7_sva_dfm_2_21_0, and_1751_cse);
  assign not_2640_nl = ~ or_dcpl_1015;
  assign and_1749_nl = MUX_v_22_2_2(22'b0000000000000000000000, mux_1495_nl, not_2640_nl);
  assign and_1452_nl = and_dcpl_1235 & and_dcpl_1402 & and_dcpl_1395;
  assign mux1h_3_nl = MUX1HOT_v_22_3_2((Silu_for_1_else_if_Silu_for_else_if_mul_cmp_1_z[44:23]),
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_21_0_mx0w1,
      act_regs_data_0_14_sva_dfm_2_21_0, {and_dcpl_1112 , and_1452_nl , and_1720_cse});
  assign not_2642_nl = ~ or_dcpl_1012;
  assign and_1752_nl = MUX_v_22_2_2(22'b0000000000000000000000, mux1h_3_nl, not_2642_nl);
  assign mux_1496_nl = MUX_v_22_2_2(ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_21_0_mx0w1,
      act_regs_data_0_15_sva_dfm_2_21_0, and_1751_cse);
  assign not_2644_nl = ~ or_dcpl_1015;
  assign and_1756_nl = MUX_v_22_2_2(22'b0000000000000000000000, mux_1496_nl, not_2644_nl);
  assign mux_1497_nl = MUX_v_22_2_2(ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_21_0_mx0w1,
      act_regs_data_0_2_sva_dfm_2_21_0, and_1751_cse);
  assign not_2646_nl = ~ or_dcpl_1015;
  assign and_1759_nl = MUX_v_22_2_2(22'b0000000000000000000000, mux_1497_nl, not_2646_nl);
  assign mux_1498_nl = MUX_v_22_2_2(ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_21_0_mx0w1,
      act_regs_data_0_3_sva_dfm_2_21_0, and_1751_cse);
  assign not_2648_nl = ~ or_dcpl_1015;
  assign and_1762_nl = MUX_v_22_2_2(22'b0000000000000000000000, mux_1498_nl, not_2648_nl);
  assign mux_1499_nl = MUX_v_22_2_2(ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_21_0_mx0w1,
      act_regs_data_0_4_sva_dfm_2_21_0, and_1751_cse);
  assign not_2650_nl = ~ or_dcpl_1015;
  assign and_1765_nl = MUX_v_22_2_2(22'b0000000000000000000000, mux_1499_nl, not_2650_nl);
  assign mux_1500_nl = MUX_v_22_2_2(ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_21_0_mx0w1,
      act_regs_data_0_5_sva_dfm_2_21_0, and_1751_cse);
  assign not_2652_nl = ~ or_dcpl_1015;
  assign and_1768_nl = MUX_v_22_2_2(22'b0000000000000000000000, mux_1500_nl, not_2652_nl);
  assign mux_1501_nl = MUX_v_22_2_2(ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_21_0_mx0w1,
      act_regs_data_0_8_sva_dfm_2_21_0, and_1751_cse);
  assign not_2654_nl = ~ or_dcpl_1015;
  assign and_1771_nl = MUX_v_22_2_2(22'b0000000000000000000000, mux_1501_nl, not_2654_nl);
  assign mux_1502_nl = MUX_v_22_2_2(ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_21_0_mx0w1,
      act_regs_data_0_6_sva_dfm_2_21_0, and_1751_cse);
  assign not_2656_nl = ~ or_dcpl_1015;
  assign and_1774_nl = MUX_v_22_2_2(22'b0000000000000000000000, mux_1502_nl, not_2656_nl);
  assign and_1577_nl = Gelu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
      & operator_32_8_true_AC_TRN_AC_WRAP_6_less_15_tmp & Gelu_for_1_else_slc_32_svs
      & Gelu_for_1_slc_32_1_svs;
  assign mux_125_nl = MUX_s_1_2_2(mux_tmp_108, or_tmp_158, and_1577_nl);
  assign and_1578_nl = Gelu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
      & Gelu_for_1_else_slc_32_svs & Gelu_for_1_slc_32_1_svs;
  assign mux_126_nl = MUX_s_1_2_2(mux_tmp_108, or_tmp_158, and_1578_nl);
  assign and_1579_nl = Gelu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
      & operator_32_8_true_AC_TRN_AC_WRAP_6_less_14_tmp & Gelu_for_2_else_slc_32_svs
      & Gelu_for_2_slc_32_1_svs;
  assign mux_127_nl = MUX_s_1_2_2(mux_tmp_108, or_tmp_158, and_1579_nl);
  assign and_1580_nl = Gelu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
      & Gelu_for_2_else_slc_32_svs & Gelu_for_2_slc_32_1_svs;
  assign mux_128_nl = MUX_s_1_2_2(mux_tmp_108, or_tmp_158, and_1580_nl);
  assign and_1581_nl = Gelu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
      & operator_32_8_true_AC_TRN_AC_WRAP_6_less_13_tmp & Gelu_for_3_else_slc_32_svs
      & Gelu_for_3_slc_32_1_svs;
  assign mux_129_nl = MUX_s_1_2_2(mux_tmp_108, or_tmp_158, and_1581_nl);
  assign and_1582_nl = Gelu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
      & Gelu_for_3_else_slc_32_svs & Gelu_for_3_slc_32_1_svs;
  assign mux_130_nl = MUX_s_1_2_2(mux_tmp_108, or_tmp_158, and_1582_nl);
  assign and_1583_nl = Gelu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
      & operator_32_8_true_AC_TRN_AC_WRAP_6_less_12_tmp & Gelu_for_4_else_slc_32_svs
      & Gelu_for_4_slc_32_1_svs;
  assign mux_131_nl = MUX_s_1_2_2(mux_tmp_108, or_tmp_158, and_1583_nl);
  assign and_1584_nl = Gelu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
      & Gelu_for_4_else_slc_32_svs & Gelu_for_4_slc_32_1_svs;
  assign mux_132_nl = MUX_s_1_2_2(mux_tmp_108, or_tmp_158, and_1584_nl);
  assign and_1585_nl = Gelu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
      & operator_32_8_true_AC_TRN_AC_WRAP_6_less_11_tmp & Gelu_for_5_else_slc_32_svs
      & Gelu_for_5_slc_32_1_svs;
  assign mux_133_nl = MUX_s_1_2_2(mux_tmp_108, or_tmp_158, and_1585_nl);
  assign and_1586_nl = Gelu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
      & Gelu_for_5_else_slc_32_svs & Gelu_for_5_slc_32_1_svs;
  assign mux_134_nl = MUX_s_1_2_2(mux_tmp_108, or_tmp_158, and_1586_nl);
  assign and_1587_nl = Gelu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
      & operator_32_8_true_AC_TRN_AC_WRAP_6_less_10_tmp & Gelu_for_6_else_slc_32_svs
      & Gelu_for_6_slc_32_1_svs;
  assign mux_135_nl = MUX_s_1_2_2(mux_tmp_108, or_tmp_158, and_1587_nl);
  assign and_1588_nl = Gelu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
      & Gelu_for_6_else_slc_32_svs & Gelu_for_6_slc_32_1_svs;
  assign mux_136_nl = MUX_s_1_2_2(mux_tmp_108, or_tmp_158, and_1588_nl);
  assign and_1589_nl = Gelu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
      & operator_32_8_true_AC_TRN_AC_WRAP_6_less_9_tmp & Gelu_for_7_else_slc_32_svs
      & Gelu_for_7_slc_32_1_svs;
  assign mux_137_nl = MUX_s_1_2_2(mux_tmp_108, or_tmp_158, and_1589_nl);
  assign and_1590_nl = Gelu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
      & Gelu_for_7_else_slc_32_svs & Gelu_for_7_slc_32_1_svs;
  assign mux_138_nl = MUX_s_1_2_2(mux_tmp_108, or_tmp_158, and_1590_nl);
  assign and_1591_nl = Gelu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
      & operator_32_8_true_AC_TRN_AC_WRAP_6_less_8_tmp & Gelu_for_8_else_slc_32_svs
      & Gelu_for_8_slc_32_1_svs;
  assign mux_139_nl = MUX_s_1_2_2(mux_tmp_108, or_tmp_158, and_1591_nl);
  assign and_1592_nl = Gelu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_5_slc_operator_32_8_true_AC_TRN_AC_WRAP_5_acc_32_svs
      & Gelu_for_8_else_slc_32_svs & Gelu_for_8_slc_32_1_svs;
  assign mux_140_nl = MUX_s_1_2_2(mux_tmp_108, or_tmp_158, and_1592_nl);
  assign and_1593_nl = Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & operator_32_8_true_AC_TRN_AC_WRAP_6_less_7_tmp & Gelu_for_9_else_slc_32_svs
      & Gelu_for_9_slc_32_1_svs;
  assign mux_141_nl = MUX_s_1_2_2(mux_tmp_108, or_tmp_158, and_1593_nl);
  assign and_1594_nl = Silu_for_9_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & Gelu_for_9_else_slc_32_svs & Gelu_for_9_slc_32_1_svs;
  assign mux_142_nl = MUX_s_1_2_2(mux_tmp_108, or_tmp_158, and_1594_nl);
  assign and_1595_nl = Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & operator_32_8_true_AC_TRN_AC_WRAP_6_less_6_tmp & Gelu_for_10_else_slc_32_svs
      & Gelu_for_10_slc_32_1_svs;
  assign mux_143_nl = MUX_s_1_2_2(mux_tmp_108, or_tmp_158, and_1595_nl);
  assign and_1596_nl = Silu_for_10_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & Gelu_for_10_else_slc_32_svs & Gelu_for_10_slc_32_1_svs;
  assign mux_144_nl = MUX_s_1_2_2(mux_tmp_108, or_tmp_158, and_1596_nl);
  assign and_1597_nl = Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & operator_32_8_true_AC_TRN_AC_WRAP_6_less_5_tmp & Gelu_for_11_else_slc_32_svs
      & Gelu_for_11_slc_32_1_svs;
  assign mux_145_nl = MUX_s_1_2_2(mux_tmp_108, or_tmp_158, and_1597_nl);
  assign and_1598_nl = Silu_for_11_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & Gelu_for_11_else_slc_32_svs & Gelu_for_11_slc_32_1_svs;
  assign mux_146_nl = MUX_s_1_2_2(mux_tmp_108, or_tmp_158, and_1598_nl);
  assign and_1599_nl = Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & operator_32_8_true_AC_TRN_AC_WRAP_6_less_4_tmp & Gelu_for_12_else_slc_32_svs
      & Gelu_for_12_slc_32_1_svs;
  assign mux_147_nl = MUX_s_1_2_2(mux_tmp_108, or_tmp_158, and_1599_nl);
  assign and_1600_nl = Silu_for_12_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & Gelu_for_12_else_slc_32_svs & Gelu_for_12_slc_32_1_svs;
  assign mux_148_nl = MUX_s_1_2_2(mux_tmp_108, or_tmp_158, and_1600_nl);
  assign and_1601_nl = Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & operator_32_8_true_AC_TRN_AC_WRAP_6_less_3_tmp & Gelu_for_13_else_slc_32_svs
      & Gelu_for_13_slc_32_1_svs;
  assign mux_149_nl = MUX_s_1_2_2(mux_tmp_108, or_tmp_158, and_1601_nl);
  assign and_1602_nl = Silu_for_13_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & Gelu_for_13_else_slc_32_svs & Gelu_for_13_slc_32_1_svs;
  assign mux_150_nl = MUX_s_1_2_2(mux_tmp_108, or_tmp_158, and_1602_nl);
  assign and_1603_nl = Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & operator_32_8_true_AC_TRN_AC_WRAP_6_less_2_tmp & Gelu_for_14_else_slc_32_svs
      & Gelu_for_14_slc_32_1_svs;
  assign mux_151_nl = MUX_s_1_2_2(mux_tmp_108, or_tmp_158, and_1603_nl);
  assign and_1604_nl = Silu_for_14_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & Gelu_for_14_else_slc_32_svs & Gelu_for_14_slc_32_1_svs;
  assign mux_152_nl = MUX_s_1_2_2(mux_tmp_108, or_tmp_158, and_1604_nl);
  assign and_1605_nl = Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & operator_32_8_true_AC_TRN_AC_WRAP_6_less_1_tmp & Gelu_for_15_else_slc_32_svs
      & Gelu_for_15_slc_32_1_svs;
  assign mux_153_nl = MUX_s_1_2_2(mux_tmp_108, or_tmp_158, and_1605_nl);
  assign and_1606_nl = Silu_for_15_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & Gelu_for_15_else_slc_32_svs & Gelu_for_15_slc_32_1_svs;
  assign mux_154_nl = MUX_s_1_2_2(mux_tmp_108, or_tmp_158, and_1606_nl);
  assign and_1607_nl = operator_32_8_true_AC_TRN_AC_WRAP_6_less_tmp & Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & Gelu_for_16_else_slc_32_svs & Gelu_for_16_slc_32_1_svs;
  assign mux_155_nl = MUX_s_1_2_2(mux_tmp_108, or_tmp_158, and_1607_nl);
  assign and_1608_nl = Silu_for_16_operator_32_8_true_AC_TRN_AC_WRAP_2_slc_operator_32_8_true_AC_TRN_AC_WRAP_2_acc_32_svs
      & Gelu_for_16_else_slc_32_svs & Gelu_for_16_slc_32_1_svs;
  assign mux_156_nl = MUX_s_1_2_2(mux_tmp_108, or_tmp_158, and_1608_nl);
  assign ActUnit_DecodeAxiWrite_if_mux_5_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[3:2]),
      (act_config_inst_regs_16_sva_dfm_6[3:2]), not_tmp_503);
  assign ActUnit_DecodeAxiWrite_if_mux_7_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[11:10]),
      (act_config_inst_regs_17_sva_dfm_6[3:2]), not_tmp_503);
  assign ActUnit_DecodeAxiWrite_if_mux_9_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[19:18]),
      (act_config_inst_regs_18_sva_dfm_6[3:2]), not_tmp_503);
  assign ActUnit_DecodeAxiWrite_if_mux_11_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[27:26]),
      (act_config_inst_regs_19_sva_dfm_6[3:2]), not_tmp_503);
  assign ActUnit_DecodeAxiWrite_if_mux_13_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[35:34]),
      (act_config_inst_regs_20_sva_dfm_6[3:2]), not_tmp_503);
  assign ActUnit_DecodeAxiWrite_if_mux_15_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[43:42]),
      (act_config_inst_regs_21_sva_dfm_6[3:2]), not_tmp_503);
  assign ActUnit_DecodeAxiWrite_if_mux_17_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[51:50]),
      (act_config_inst_regs_22_sva_dfm_6[3:2]), not_tmp_503);
  assign ActUnit_DecodeAxiWrite_if_mux_19_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[59:58]),
      (act_config_inst_regs_23_sva_dfm_6[3:2]), not_tmp_503);
  assign ActUnit_DecodeAxiWrite_if_mux_21_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[67:66]),
      (act_config_inst_regs_24_sva_dfm_6[3:2]), not_tmp_503);
  assign ActUnit_DecodeAxiWrite_if_mux_23_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[75:74]),
      (act_config_inst_regs_25_sva_dfm_6[3:2]), not_tmp_503);
  assign ActUnit_DecodeAxiWrite_if_mux_25_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[83:82]),
      (act_config_inst_regs_26_sva_dfm_6[3:2]), not_tmp_503);
  assign ActUnit_DecodeAxiWrite_if_mux_27_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[91:90]),
      (act_config_inst_regs_27_sva_dfm_6[3:2]), not_tmp_503);
  assign ActUnit_DecodeAxiWrite_if_mux_29_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[99:98]),
      (act_config_inst_regs_28_sva_dfm_6[3:2]), not_tmp_503);
  assign ActUnit_DecodeAxiWrite_if_mux_31_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[107:106]),
      (act_config_inst_regs_29_sva_dfm_6[3:2]), not_tmp_503);
  assign ActUnit_DecodeAxiWrite_if_mux_33_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[115:114]),
      (act_config_inst_regs_30_sva_dfm_6[3:2]), not_tmp_503);
  assign ActUnit_DecodeAxiWrite_if_mux_35_nl = MUX_v_2_2_2((rva_in_PopNB_mioi_data_data_rsc_z_mxwt[123:122]),
      (act_config_inst_regs_31_sva_dfm_6[3:2]), not_tmp_503);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_231_nl = act_regs_data_3_9_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_3_0_sva_dfm_2_31, and_dcpl_1270);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_229_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_3_9_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_230_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_3_9_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_69_nl = act_regs_data_3_9_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_338_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_3_9_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_291_nl = act_regs_data_3_14_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_4_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_2_15_sva_dfm_2_31, and_dcpl_1277);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_289_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_3_14_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_290_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_3_14_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_104_nl = act_regs_data_3_14_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_336_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_3_14_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_279_nl = act_regs_data_3_13_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_8_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_2_14_sva_dfm_2_31, and_dcpl_1280);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_277_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_3_13_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_278_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_3_13_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_97_nl = act_regs_data_3_13_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_334_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_3_13_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_267_nl = act_regs_data_3_12_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_12_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_2_13_sva_dfm_2_31, and_dcpl_1284);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_265_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_3_12_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_266_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_3_12_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_90_nl = act_regs_data_3_12_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_332_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_3_12_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_255_nl = act_regs_data_3_11_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_16_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_2_12_sva_dfm_2_31, and_dcpl_1287);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_253_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_3_11_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_254_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_3_11_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_83_nl = act_regs_data_3_11_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_330_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_3_11_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_243_nl = act_regs_data_3_10_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_20_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_2_11_sva_dfm_2_31, and_dcpl_1291);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_241_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_3_10_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_242_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_3_10_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_76_nl = act_regs_data_3_10_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_328_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_3_10_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_132_nl = act_regs_data_3_1_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_24_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_2_10_sva_dfm_2_31, and_dcpl_1294);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_130_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_3_1_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_131_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_3_1_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_12_nl = act_regs_data_3_1_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_326_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_3_1_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_219_nl = act_regs_data_3_8_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_28_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_2_9_sva_dfm_2_31, and_dcpl_1297);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_217_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_3_8_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_218_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_3_8_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_62_nl = act_regs_data_3_8_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_324_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_3_8_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_204_nl = act_regs_data_3_7_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_32_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_2_8_sva_dfm_2_31, and_dcpl_1299);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_202_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_3_7_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_203_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_3_7_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_54_nl = act_regs_data_3_7_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_322_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_3_7_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_192_nl = act_regs_data_3_6_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_36_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_2_7_sva_dfm_2_31, and_dcpl_1302);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_190_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_3_6_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_191_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_3_6_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_47_nl = act_regs_data_3_6_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_320_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_3_6_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_180_nl = act_regs_data_3_5_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_40_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_2_6_sva_dfm_2_31, and_dcpl_1304);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_178_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_3_5_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_179_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_3_5_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_40_nl = act_regs_data_3_5_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_318_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_3_5_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_168_nl = act_regs_data_3_4_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_44_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_2_5_sva_dfm_2_31, and_dcpl_1306);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_166_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_3_4_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_167_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_3_4_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_33_nl = act_regs_data_3_4_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_316_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_3_4_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_156_nl = act_regs_data_3_3_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_48_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_2_4_sva_dfm_2_31, and_dcpl_1308);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_154_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_3_3_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_155_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_3_3_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_26_nl = act_regs_data_3_3_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_314_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_3_3_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_144_nl = act_regs_data_3_2_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_52_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_2_3_sva_dfm_2_31, and_dcpl_1310);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_142_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_3_2_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_143_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_3_2_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_19_nl = act_regs_data_3_2_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_312_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_3_2_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_303_nl = act_regs_data_3_15_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_56_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_2_2_sva_dfm_2_31, and_dcpl_1312);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_301_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_3_15_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_302_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_3_15_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_111_nl = act_regs_data_3_15_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_310_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_3_15_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_120_nl = act_regs_data_3_0_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_60_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_2_1_sva_dfm_2_31, and_dcpl_1314);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_118_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_3_0_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_119_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_3_0_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_5_nl = act_regs_data_3_0_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_308_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_3_0_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_289);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_225_nl = act_regs_data_2_9_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_64_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_2_0_sva_dfm_2_31, and_dcpl_1316);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_223_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_2_9_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_224_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_2_9_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_67_nl = act_regs_data_2_9_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_306_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_2_9_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_285_nl = act_regs_data_2_14_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_68_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_1_15_sva_dfm_2_31, and_dcpl_1320);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_283_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_2_14_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_284_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_2_14_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_102_nl = act_regs_data_2_14_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_305_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_2_14_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_273_nl = act_regs_data_2_13_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_72_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_1_14_sva_dfm_2_31, and_dcpl_1322);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_271_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_2_13_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_272_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_2_13_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_95_nl = act_regs_data_2_13_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_307_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_2_13_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_261_nl = act_regs_data_2_12_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_76_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_1_13_sva_dfm_2_31, and_dcpl_1324);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_259_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_2_12_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_260_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_2_12_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_88_nl = act_regs_data_2_12_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_309_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_2_12_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_249_nl = act_regs_data_2_11_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_80_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_1_12_sva_dfm_2_31, and_dcpl_1326);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_247_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_2_11_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_248_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_2_11_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_81_nl = act_regs_data_2_11_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_311_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_2_11_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_237_nl = act_regs_data_2_10_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_84_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_1_11_sva_dfm_2_31, and_dcpl_1328);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_235_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_2_10_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_236_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_2_10_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_74_nl = act_regs_data_2_10_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_313_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_2_10_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_126_nl = act_regs_data_2_1_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_88_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_1_10_sva_dfm_2_31, and_dcpl_1330);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_124_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_2_1_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_125_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_2_1_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_10_nl = act_regs_data_2_1_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_315_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_2_1_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_213_nl = act_regs_data_2_8_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_92_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_1_9_sva_dfm_2_31, and_dcpl_1332);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_211_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_2_8_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_212_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_2_8_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_60_nl = act_regs_data_2_8_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_317_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_2_8_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_198_nl = act_regs_data_2_7_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_96_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_1_8_sva_dfm_2_31, and_dcpl_1334);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_196_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_2_7_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_197_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_2_7_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_52_nl = act_regs_data_2_7_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_319_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_2_7_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_186_nl = act_regs_data_2_6_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_100_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_1_7_sva_dfm_2_31, and_dcpl_1338);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_184_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_2_6_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_185_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_2_6_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_45_nl = act_regs_data_2_6_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_321_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_2_6_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_174_nl = act_regs_data_2_5_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_104_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_1_6_sva_dfm_2_31, and_dcpl_1340);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_172_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_2_5_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_173_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_2_5_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_38_nl = act_regs_data_2_5_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_323_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_2_5_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_162_nl = act_regs_data_2_4_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_108_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_1_5_sva_dfm_2_31, and_dcpl_1342);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_160_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_2_4_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_161_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_2_4_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_31_nl = act_regs_data_2_4_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_325_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_2_4_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_150_nl = act_regs_data_2_3_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_112_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_1_4_sva_dfm_2_31, and_dcpl_1344);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_148_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_2_3_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_149_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_2_3_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_24_nl = act_regs_data_2_3_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_327_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_2_3_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_138_nl = act_regs_data_2_2_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_116_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_1_3_sva_dfm_2_31, and_dcpl_1346);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_136_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_2_2_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_137_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_2_2_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_17_nl = act_regs_data_2_2_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_329_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_2_2_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_297_nl = act_regs_data_2_15_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_120_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_1_2_sva_dfm_2_31, and_dcpl_1348);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_295_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_2_15_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_296_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_2_15_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_109_nl = act_regs_data_2_15_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_331_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_2_15_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_114_nl = act_regs_data_2_0_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_124_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_1_1_sva_dfm_2_31, and_dcpl_1350);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_112_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_2_0_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_113_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_2_0_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_3_nl = act_regs_data_2_0_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_333_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_2_0_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_293);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_222_nl = act_regs_data_1_9_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_128_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_1_0_sva_dfm_2_31, and_dcpl_1352);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_220_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_1_9_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_221_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_1_9_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_66_nl = act_regs_data_1_9_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_335_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_1_9_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_282_nl = act_regs_data_1_14_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_132_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_0_15_sva_dfm_2_31, and_dcpl_1355);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_280_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_1_14_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_281_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_1_14_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_101_nl = act_regs_data_1_14_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_337_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_1_14_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_270_nl = act_regs_data_1_13_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_136_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_0_14_sva_dfm_2_31, and_dcpl_1357);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_268_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_1_13_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_269_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_1_13_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_94_nl = act_regs_data_1_13_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_339_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_1_13_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_258_nl = act_regs_data_1_12_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_140_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_0_13_sva_dfm_2_31, and_dcpl_1359);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_256_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_1_12_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_257_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_1_12_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_87_nl = act_regs_data_1_12_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_340_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_1_12_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_246_nl = act_regs_data_1_11_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_144_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_0_12_sva_dfm_2_31, and_dcpl_1361);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_244_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_1_11_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_245_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_1_11_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_80_nl = act_regs_data_1_11_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_341_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_1_11_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_234_nl = act_regs_data_1_10_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_148_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_0_11_sva_dfm_2_31, and_dcpl_1363);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_232_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_1_10_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_233_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_1_10_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_73_nl = act_regs_data_1_10_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_342_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_1_10_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_129_nl = act_regs_data_1_1_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_152_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_0_10_sva_dfm_2_31, and_dcpl_1365);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_127_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_1_1_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_128_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_1_1_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_11_nl = act_regs_data_1_1_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_343_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_1_1_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_210_nl = act_regs_data_1_8_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_156_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_0_9_sva_dfm_2_31, and_dcpl_1367);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_208_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_1_8_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_209_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_1_8_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_59_nl = act_regs_data_1_8_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_344_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_1_8_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_201_nl = act_regs_data_1_7_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_160_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_0_8_sva_dfm_2_31, and_dcpl_1369);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_199_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_1_7_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_200_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_1_7_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_53_nl = act_regs_data_1_7_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_345_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_1_7_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_189_nl = act_regs_data_1_6_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_164_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_0_7_sva_dfm_2_31, and_dcpl_1372);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_187_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_1_6_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_188_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_1_6_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_46_nl = act_regs_data_1_6_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_346_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_1_6_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_177_nl = act_regs_data_1_5_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_168_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_0_6_sva_dfm_2_31, and_dcpl_1374);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_175_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_1_5_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_176_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_1_5_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_39_nl = act_regs_data_1_5_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_347_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_1_5_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_165_nl = act_regs_data_1_4_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_172_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_0_5_sva_dfm_2_31, and_dcpl_1376);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_163_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_1_4_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_164_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_1_4_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_32_nl = act_regs_data_1_4_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_348_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_1_4_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_153_nl = act_regs_data_1_3_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_176_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_0_4_sva_dfm_2_31, and_dcpl_1378);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_151_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_1_3_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_152_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_1_3_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_25_nl = act_regs_data_1_3_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_349_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_1_3_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_141_nl = act_regs_data_1_2_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_180_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_0_3_sva_dfm_2_31, and_dcpl_1380);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_139_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_1_2_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_140_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_1_2_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_18_nl = act_regs_data_1_2_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_350_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_1_2_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_294_nl = act_regs_data_1_15_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_184_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_0_2_sva_dfm_2_31, and_dcpl_1382);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_292_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_1_15_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_293_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_1_15_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_108_nl = act_regs_data_1_15_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_351_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_1_15_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_117_nl = act_regs_data_1_0_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_188_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_0_1_sva_dfm_2_31, and_dcpl_1384);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_115_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_1_0_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_116_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_1_0_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_4_nl = act_regs_data_1_0_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_352_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_1_0_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_295);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_228_nl = act_regs_data_0_9_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_291;
  assign ActUnit_RunLoad_if_else_for_ActUnit_RunLoad_if_else_for_mux_192_nl = MUX_s_1_2_2((ActUnit_RunLoad_if_else_for_slc_act_port_read_out_data_32_31_0_2_ctmp_sva_1[31]),
      act_regs_data_0_0_sva_dfm_2_31, and_dcpl_1386);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_226_nl = MUX_v_5_2_2(5'b00000,
      act_regs_data_0_9_sva_dfm_2_30_26, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_291);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_227_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_0_9_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_291);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_68_nl = act_regs_data_0_9_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_291;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_353_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_0_9_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_291);
  assign while_and_64_nl = act_config_InstIncr_act_config_InstIncr_if_and_svs_1 &
      is_incr_lpi_1_dfm_1 & is_start_sva;
  assign or_1426_nl = (fsm_output[2:0]!=3'b001);
  assign mux_451_nl = MUX_s_1_2_2(not_tmp_620, or_1426_nl, fsm_output[3]);
  assign Silu_for_else_mux_32_nl = MUX_s_1_2_2((Silu_for_y_8_sva_1_22_0_1[22]), (Silu_for_8_else_else_if_acc_itm[1]),
      Silu_for_else_and_14_ssc_1);
  assign Silu_for_else_Silu_for_else_mux1h_39_nl = MUX1HOT_v_2_4_2((Silu_for_y_8_sva_1_22_0_1[21:20]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1[1:0]),
      (Silu_for_y_8_sva_3_21_0[21:20]), (reg_nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:20]),
      {(~ Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_14_ssc_1 , Silu_for_else_and_39_ssc_1 , Silu_for_else_or_7_itm});
  assign Silu_for_else_Silu_for_else_mux1h_48_nl = MUX1HOT_v_20_4_2((Silu_for_y_8_sva_1_22_0_1[19:0]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:2]),
      (Silu_for_y_8_sva_3_21_0[19:0]), (reg_nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[19:0]),
      {(~ Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_14_ssc_1 , Silu_for_else_and_39_ssc_1 , Silu_for_else_or_7_itm});
  assign Silu_for_else_mux_33_nl = MUX_s_1_2_2((Silu_for_y_7_sva_1_22_0_1[22]), (Silu_for_7_else_else_if_acc_itm[1]),
      Silu_for_else_and_12_ssc_1);
  assign Silu_for_else_Silu_for_else_mux1h_38_nl = MUX1HOT_v_2_4_2((Silu_for_y_7_sva_1_22_0_1[21:20]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1[1:0]),
      (Silu_for_7_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0[21:20]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:20]),
      {(~ Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_12_ssc_1 , Silu_for_else_and_38_ssc_1 , Silu_for_else_or_6_itm});
  assign Silu_for_else_Silu_for_else_mux1h_50_nl = MUX1HOT_v_20_4_2((Silu_for_y_7_sva_1_22_0_1[19:0]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:2]),
      (Silu_for_7_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0[19:0]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[19:0]),
      {(~ Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_12_ssc_1 , Silu_for_else_and_38_ssc_1 , Silu_for_else_or_6_itm});
  assign Silu_for_else_mux_34_nl = MUX_s_1_2_2((Silu_for_y_6_sva_1_22_0_1[22]), (Silu_for_6_else_else_if_acc_itm[1]),
      Silu_for_else_and_10_ssc_1);
  assign Silu_for_else_Silu_for_else_mux1h_37_nl = MUX1HOT_v_2_4_2((Silu_for_y_6_sva_1_22_0_1[21:20]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1[1:0]),
      (Silu_for_6_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0[21:20]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:20]),
      {(~ Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_10_ssc_1 , Silu_for_else_and_37_ssc_1 , Silu_for_else_or_5_itm});
  assign Silu_for_else_Silu_for_else_mux1h_52_nl = MUX1HOT_v_20_4_2((Silu_for_y_6_sva_1_22_0_1[19:0]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:2]),
      (Silu_for_6_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0[19:0]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[19:0]),
      {(~ Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_10_ssc_1 , Silu_for_else_and_37_ssc_1 , Silu_for_else_or_5_itm});
  assign Silu_for_else_mux_35_nl = MUX_s_1_2_2((Silu_for_y_5_sva_1_22_0_1[22]), (Silu_for_5_else_else_if_acc_itm[1]),
      Silu_for_else_and_8_ssc_1);
  assign Silu_for_else_Silu_for_else_mux1h_36_nl = MUX1HOT_v_2_4_2((Silu_for_y_5_sva_1_22_0_1[21:20]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1[1:0]),
      (Silu_for_5_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0[21:20]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:20]),
      {(~ Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_8_ssc_1 , Silu_for_else_and_36_ssc_1 , Silu_for_else_or_4_itm});
  assign Silu_for_else_Silu_for_else_mux1h_54_nl = MUX1HOT_v_20_4_2((Silu_for_y_5_sva_1_22_0_1[19:0]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:2]),
      (Silu_for_5_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0[19:0]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[19:0]),
      {(~ Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_8_ssc_1 , Silu_for_else_and_36_ssc_1 , Silu_for_else_or_4_itm});
  assign Silu_for_else_mux_36_nl = MUX_s_1_2_2((Silu_for_y_4_sva_1_22_0_1[22]), (Silu_for_4_else_else_if_acc_itm[1]),
      Silu_for_else_and_6_ssc_1);
  assign Silu_for_else_Silu_for_else_mux1h_35_nl = MUX1HOT_v_2_4_2((Silu_for_y_4_sva_1_22_0_1[21:20]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1[1:0]),
      (Silu_for_4_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0[21:20]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:20]),
      {(~ Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_6_ssc_1 , Silu_for_else_and_35_ssc_1 , Silu_for_else_or_3_itm});
  assign Silu_for_else_Silu_for_else_mux1h_56_nl = MUX1HOT_v_20_4_2((Silu_for_y_4_sva_1_22_0_1[19:0]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:2]),
      (Silu_for_4_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0[19:0]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[19:0]),
      {(~ Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_6_ssc_1 , Silu_for_else_and_35_ssc_1 , Silu_for_else_or_3_itm});
  assign Silu_for_else_mux_37_nl = MUX_s_1_2_2((Silu_for_y_3_sva_1_22_0_1[22]), (Silu_for_3_else_else_if_acc_itm[1]),
      Silu_for_else_and_4_ssc_1);
  assign Silu_for_else_Silu_for_else_mux1h_34_nl = MUX1HOT_v_2_4_2((Silu_for_y_3_sva_1_22_0_1[21:20]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1[1:0]),
      (Silu_for_3_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0[21:20]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:20]),
      {(~ Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_4_ssc_1 , Silu_for_else_and_34_ssc_1 , Silu_for_else_or_2_itm});
  assign Silu_for_else_Silu_for_else_mux1h_58_nl = MUX1HOT_v_20_4_2((Silu_for_y_3_sva_1_22_0_1[19:0]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:2]),
      (Silu_for_3_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0[19:0]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[19:0]),
      {(~ Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_4_ssc_1 , Silu_for_else_and_34_ssc_1 , Silu_for_else_or_2_itm});
  assign Silu_for_else_mux_38_nl = MUX_s_1_2_2((Silu_for_y_2_sva_1_22_0_1[22]), (Silu_for_2_else_else_if_acc_itm[1]),
      Silu_for_else_and_2_ssc_1);
  assign Silu_for_else_Silu_for_else_mux1h_33_nl = MUX1HOT_v_2_4_2((Silu_for_y_2_sva_1_22_0_1[21:20]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_2_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1[1:0]),
      (Silu_for_2_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0[21:20]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_2_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:20]),
      {(~ Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_2_ssc_1 , Silu_for_else_and_33_ssc_1 , Silu_for_else_or_1_itm});
  assign Silu_for_else_Silu_for_else_mux1h_60_nl = MUX1HOT_v_20_4_2((Silu_for_y_2_sva_1_22_0_1[19:0]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_2_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[21:2]),
      (Silu_for_2_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_21_0[19:0]),
      (reg_nv_scvector_cctor_nv_scvector_5_for_2_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_1[19:0]),
      {(~ Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_2_ssc_1 , Silu_for_else_and_33_ssc_1 , Silu_for_else_or_1_itm});
  assign Silu_for_else_mux_39_nl = MUX_s_1_2_2((Silu_for_y_1_sva_1_22_0_1[22]), (Silu_for_1_else_else_if_acc_itm[1]),
      Silu_for_else_and_ssc_1);
  assign Silu_for_else_Silu_for_else_mux1h_32_nl = MUX1HOT_v_2_4_2((Silu_for_y_1_sva_1_22_0_1[21:20]),
      (reg_ActUnit_RunInst_case_14_nv_scvector_cctor_data_0_1_ftd_rsp_1[1:0]), (Silu_for_y_1_sva_3_21_0[21:20]),
      (reg_ActUnit_RunInst_case_14_nv_scvector_cctor_data_0_1_ftd_1[21:20]), {(~
      Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_ssc_1 , Silu_for_else_and_32_ssc_1 , Silu_for_else_or_itm});
  assign Silu_for_else_Silu_for_else_mux1h_62_nl = MUX1HOT_v_20_4_2((Silu_for_y_1_sva_1_22_0_1[19:0]),
      (reg_ActUnit_RunInst_case_14_nv_scvector_cctor_data_0_1_ftd_1[21:2]), (Silu_for_y_1_sva_3_21_0[19:0]),
      (reg_ActUnit_RunInst_case_14_nv_scvector_cctor_data_0_1_ftd_1[19:0]), {(~ Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_ssc_1 , Silu_for_else_and_32_ssc_1 , Silu_for_else_or_itm});
  assign Silu_for_else_Silu_for_else_mux1h_23_nl = MUX1HOT_s_1_4_2((Silu_for_y_8_sva_1_22_0_1[22]),
      (Silu_for_8_else_else_if_acc_itm[1]), ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_1_25,
      reg_nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0,
      {(~ Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_14_ssc_1 , Silu_for_else_else_else_and_14_ssc_1 , Silu_for_else_else_else_and_15_ssc_1});
  assign Silu_for_else_Silu_for_else_mux1h_49_nl = MUX1HOT_v_3_5_2((signext_3_1(Silu_for_y_8_sva_1_22_0_1[22])),
      ({{1{Silu_for_8_else_else_if_acc_itm[1]}}, Silu_for_8_else_else_if_acc_itm}),
      Silu_for_y_8_sva_3_24_22, ActUnit_PushOutput_if_output_port_reg_data_data_7_sva_1_24_22,
      reg_nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1,
      {(~ Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_14_ssc_1 , Silu_for_else_and_39_ssc_1 , Silu_for_else_else_else_and_14_ssc_1
      , Silu_for_else_else_else_and_15_ssc_1});
  assign Silu_for_else_Silu_for_else_mux1h_22_nl = MUX1HOT_s_1_4_2((Silu_for_y_7_sva_1_22_0_1[22]),
      (Silu_for_7_else_else_if_acc_itm[1]), ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_1_25,
      reg_nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0,
      {(~ Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_12_ssc_1 , Silu_for_else_else_else_and_12_ssc_1 , Silu_for_else_else_else_and_13_ssc_1});
  assign Silu_for_else_Silu_for_else_mux1h_51_nl = MUX1HOT_v_3_5_2((signext_3_1(Silu_for_y_7_sva_1_22_0_1[22])),
      ({{1{Silu_for_7_else_else_if_acc_itm[1]}}, Silu_for_7_else_else_if_acc_itm}),
      Silu_for_7_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_24_22,
      ActUnit_PushOutput_if_output_port_reg_data_data_6_sva_1_24_22, reg_nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1,
      {(~ Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_12_ssc_1 , Silu_for_else_and_38_ssc_1 , Silu_for_else_else_else_and_12_ssc_1
      , Silu_for_else_else_else_and_13_ssc_1});
  assign Silu_for_else_Silu_for_else_mux1h_21_nl = MUX1HOT_s_1_4_2((Silu_for_y_6_sva_1_22_0_1[22]),
      (Silu_for_6_else_else_if_acc_itm[1]), ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_1_25,
      reg_nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0,
      {(~ Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_10_ssc_1 , Silu_for_else_else_else_and_10_ssc_1 , Silu_for_else_else_else_and_11_ssc_1});
  assign Silu_for_else_Silu_for_else_mux1h_53_nl = MUX1HOT_v_3_5_2((signext_3_1(Silu_for_y_6_sva_1_22_0_1[22])),
      ({{1{Silu_for_6_else_else_if_acc_itm[1]}}, Silu_for_6_else_else_if_acc_itm}),
      Silu_for_6_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_24_22,
      ActUnit_PushOutput_if_output_port_reg_data_data_5_sva_1_24_22, reg_nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1,
      {(~ Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_10_ssc_1 , Silu_for_else_and_37_ssc_1 , Silu_for_else_else_else_and_10_ssc_1
      , Silu_for_else_else_else_and_11_ssc_1});
  assign Silu_for_else_Silu_for_else_mux1h_20_nl = MUX1HOT_s_1_4_2((Silu_for_y_5_sva_1_22_0_1[22]),
      (Silu_for_5_else_else_if_acc_itm[1]), ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_1_25,
      reg_nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0,
      {(~ Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_8_ssc_1 , Silu_for_else_else_else_and_8_ssc_1 , Silu_for_else_else_else_and_9_ssc_1});
  assign Silu_for_else_Silu_for_else_mux1h_55_nl = MUX1HOT_v_3_5_2((signext_3_1(Silu_for_y_5_sva_1_22_0_1[22])),
      ({{1{Silu_for_5_else_else_if_acc_itm[1]}}, Silu_for_5_else_else_if_acc_itm}),
      Silu_for_5_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_24_22,
      ActUnit_PushOutput_if_output_port_reg_data_data_4_sva_1_24_22, reg_nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1,
      {(~ Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_8_ssc_1 , Silu_for_else_and_36_ssc_1 , Silu_for_else_else_else_and_8_ssc_1
      , Silu_for_else_else_else_and_9_ssc_1});
  assign Silu_for_else_Silu_for_else_mux1h_19_nl = MUX1HOT_s_1_4_2((Silu_for_y_4_sva_1_22_0_1[22]),
      (Silu_for_4_else_else_if_acc_itm[1]), ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_1_25,
      reg_nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0,
      {(~ Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_6_ssc_1 , Silu_for_else_else_else_and_6_ssc_1 , Silu_for_else_else_else_and_7_ssc_1});
  assign Silu_for_else_Silu_for_else_mux1h_57_nl = MUX1HOT_v_3_5_2((signext_3_1(Silu_for_y_4_sva_1_22_0_1[22])),
      ({{1{Silu_for_4_else_else_if_acc_itm[1]}}, Silu_for_4_else_else_if_acc_itm}),
      Silu_for_4_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_24_22,
      ActUnit_PushOutput_if_output_port_reg_data_data_3_sva_1_24_22, reg_nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1,
      {(~ Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_6_ssc_1 , Silu_for_else_and_35_ssc_1 , Silu_for_else_else_else_and_6_ssc_1
      , Silu_for_else_else_else_and_7_ssc_1});
  assign Silu_for_else_Silu_for_else_mux1h_18_nl = MUX1HOT_s_1_4_2((Silu_for_y_3_sva_1_22_0_1[22]),
      (Silu_for_3_else_else_if_acc_itm[1]), ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_1_25,
      reg_nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0,
      {(~ Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_4_ssc_1 , Silu_for_else_else_else_and_4_ssc_1 , Silu_for_else_else_else_and_5_ssc_1});
  assign Silu_for_else_Silu_for_else_mux1h_59_nl = MUX1HOT_v_3_5_2((signext_3_1(Silu_for_y_3_sva_1_22_0_1[22])),
      ({{1{Silu_for_3_else_else_if_acc_itm[1]}}, Silu_for_3_else_else_if_acc_itm}),
      Silu_for_3_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_24_22,
      ActUnit_PushOutput_if_output_port_reg_data_data_2_sva_1_24_22, reg_nv_scvector_cctor_nv_scvector_5_for_3_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1,
      {(~ Silu_for_3_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_4_ssc_1 , Silu_for_else_and_34_ssc_1 , Silu_for_else_else_else_and_4_ssc_1
      , Silu_for_else_else_else_and_5_ssc_1});
  assign Silu_for_else_Silu_for_else_mux1h_17_nl = MUX1HOT_s_1_4_2((Silu_for_y_2_sva_1_22_0_1[22]),
      (Silu_for_2_else_else_if_acc_itm[1]), ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_1_25,
      reg_nv_scvector_cctor_nv_scvector_5_for_2_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0,
      {(~ Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_2_ssc_1 , Silu_for_else_else_else_and_2_ssc_1 , Silu_for_else_else_else_and_3_ssc_1});
  assign Silu_for_else_Silu_for_else_mux1h_61_nl = MUX1HOT_v_3_5_2((signext_3_1(Silu_for_y_2_sva_1_22_0_1[22])),
      ({{1{Silu_for_2_else_else_if_acc_itm[1]}}, Silu_for_2_else_else_if_acc_itm}),
      Silu_for_2_else_else_else_if_slc_Silu_for_else_else_else_if_acc_32_1_itm_24_22,
      ActUnit_PushOutput_if_output_port_reg_data_data_14_sva_1_24_22, reg_nv_scvector_cctor_nv_scvector_5_for_2_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1,
      {(~ Silu_for_2_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_2_ssc_1 , Silu_for_else_and_33_ssc_1 , Silu_for_else_else_else_and_2_ssc_1
      , Silu_for_else_else_else_and_3_ssc_1});
  assign Silu_for_else_Silu_for_else_mux1h_16_nl = MUX1HOT_s_1_4_2((Silu_for_y_1_sva_1_22_0_1[22]),
      (Silu_for_1_else_else_if_acc_itm[1]), ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_1_25,
      reg_ActUnit_RunInst_case_14_nv_scvector_cctor_data_0_1_ftd_rsp_0, {(~ Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_ssc_1 , Silu_for_else_else_else_and_ssc_1 , Silu_for_else_else_else_and_1_ssc_1});
  assign Silu_for_else_Silu_for_else_mux1h_63_nl = MUX1HOT_v_3_5_2((signext_3_1(Silu_for_y_1_sva_1_22_0_1[22])),
      ({{1{Silu_for_1_else_else_if_acc_itm[1]}}, Silu_for_1_else_else_if_acc_itm}),
      Silu_for_y_1_sva_3_24_22, ActUnit_PushOutput_if_output_port_reg_data_data_13_sva_1_24_22,
      reg_ActUnit_RunInst_case_14_nv_scvector_cctor_data_0_1_ftd_rsp_1, {(~ Silu_for_1_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_ssc_1 , Silu_for_else_and_32_ssc_1 , Silu_for_else_else_else_and_ssc_1
      , Silu_for_else_else_else_and_1_ssc_1});
  assign Silu_for_else_Silu_for_else_mux1h_3_nl = MUX1HOT_v_5_3_2((signext_5_1(Silu_for_y_4_sva_1_22_0_1[22])),
      (signext_5_1(Silu_for_4_else_else_if_acc_itm[1])), reg_nv_scvector_cctor_nv_scvector_5_for_4_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26,
      {(~ Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_6_ssc_1 , Silu_for_else_else_else_and_7_ssc_1});
  assign Silu_for_else_nor_7_nl = ~(Silu_for_else_and_35_ssc_1 | Silu_for_else_else_else_and_6_ssc_1);
  assign Silu_for_Silu_for_and_25_nl = Silu_for_else_Silu_for_else_mux1h_3_nl & (signext_5_1(Silu_for_else_nor_7_nl))
      & ({{4{Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs}},
      Silu_for_4_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs});
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_70_nl = MUX1HOT_v_5_3_2(Silu_for_Silu_for_and_25_nl,
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_30_26_2, act_regs_data_0_10_sva_dfm_2_30_26,
      {and_dcpl_1112 , and_dcpl_1235 , and_dcpl_1236});
  assign not_8877_nl = ~ or_dcpl;
  assign Silu_for_else_Silu_for_else_mux1h_4_nl = MUX1HOT_v_5_3_2((signext_5_1(Silu_for_y_5_sva_1_22_0_1[22])),
      (signext_5_1(Silu_for_5_else_else_if_acc_itm[1])), reg_nv_scvector_cctor_nv_scvector_5_for_5_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26,
      {(~ Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_8_ssc_1 , Silu_for_else_else_else_and_9_ssc_1});
  assign Silu_for_else_nor_9_nl = ~(Silu_for_else_and_36_ssc_1 | Silu_for_else_else_else_and_8_ssc_1);
  assign Silu_for_Silu_for_and_28_nl = Silu_for_else_Silu_for_else_mux1h_4_nl & (signext_5_1(Silu_for_else_nor_9_nl))
      & ({{4{Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs}},
      Silu_for_5_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs});
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_75_nl = MUX1HOT_v_5_3_2(Silu_for_Silu_for_and_28_nl,
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_30_26_2, act_regs_data_0_11_sva_dfm_2_30_26,
      {and_dcpl_1112 , and_dcpl_1235 , and_dcpl_1236});
  assign not_8878_nl = ~ or_dcpl;
  assign Silu_for_else_Silu_for_else_mux1h_5_nl = MUX1HOT_v_5_3_2((signext_5_1(Silu_for_y_6_sva_1_22_0_1[22])),
      (signext_5_1(Silu_for_6_else_else_if_acc_itm[1])), reg_nv_scvector_cctor_nv_scvector_5_for_6_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26,
      {(~ Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_10_ssc_1 , Silu_for_else_else_else_and_11_ssc_1});
  assign Silu_for_else_nor_11_nl = ~(Silu_for_else_and_37_ssc_1 | Silu_for_else_else_else_and_10_ssc_1);
  assign Silu_for_Silu_for_and_31_nl = Silu_for_else_Silu_for_else_mux1h_5_nl & (signext_5_1(Silu_for_else_nor_11_nl))
      & ({{4{Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs}},
      Silu_for_6_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs});
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_80_nl = MUX1HOT_v_5_3_2(Silu_for_Silu_for_and_31_nl,
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_30_26_2, act_regs_data_0_12_sva_dfm_2_30_26,
      {and_dcpl_1112 , and_dcpl_1235 , and_dcpl_1236});
  assign not_8879_nl = ~ or_dcpl;
  assign Silu_for_else_Silu_for_else_mux1h_6_nl = MUX1HOT_v_5_3_2((signext_5_1(Silu_for_y_7_sva_1_22_0_1[22])),
      (signext_5_1(Silu_for_7_else_else_if_acc_itm[1])), reg_nv_scvector_cctor_nv_scvector_5_for_7_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26,
      {(~ Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_12_ssc_1 , Silu_for_else_else_else_and_13_ssc_1});
  assign Silu_for_else_nor_13_nl = ~(Silu_for_else_and_38_ssc_1 | Silu_for_else_else_else_and_12_ssc_1);
  assign Silu_for_Silu_for_and_34_nl = Silu_for_else_Silu_for_else_mux1h_6_nl & (signext_5_1(Silu_for_else_nor_13_nl))
      & ({{4{Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs}},
      Silu_for_7_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs});
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_85_nl = MUX1HOT_v_5_3_2(Silu_for_Silu_for_and_34_nl,
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_30_26_2, act_regs_data_0_13_sva_dfm_2_30_26,
      {and_dcpl_1112 , and_dcpl_1235 , and_dcpl_1236});
  assign not_8880_nl = ~ or_dcpl;
  assign Silu_for_else_Silu_for_else_mux1h_7_nl = MUX1HOT_v_5_3_2((signext_5_1(Silu_for_y_8_sva_1_22_0_1[22])),
      (signext_5_1(Silu_for_8_else_else_if_acc_itm[1])), reg_nv_scvector_cctor_nv_scvector_5_for_8_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_ftd_1_30_26,
      {(~ Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_1_slc_operator_32_8_true_AC_TRN_AC_WRAP_1_acc_32_svs)
      , Silu_for_else_and_14_ssc_1 , Silu_for_else_else_else_and_15_ssc_1});
  assign Silu_for_else_nor_15_nl = ~(Silu_for_else_and_39_ssc_1 | Silu_for_else_else_else_and_14_ssc_1);
  assign Silu_for_Silu_for_and_37_nl = Silu_for_else_Silu_for_else_mux1h_7_nl & (signext_5_1(Silu_for_else_nor_15_nl))
      & ({{4{Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs}},
      Silu_for_8_operator_32_8_true_AC_TRN_AC_WRAP_slc_operator_32_8_true_AC_TRN_AC_WRAP_acc_32_svs});
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_90_nl = MUX1HOT_v_5_3_2(Silu_for_Silu_for_and_37_nl,
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_30_26_2, act_regs_data_0_14_sva_dfm_2_30_26,
      {and_dcpl_1112 , and_dcpl_1235 , and_dcpl_1236});
  assign not_8881_nl = ~ or_dcpl;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_123_nl = act_regs_data_0_0_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_291;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_288_nl = act_regs_data_0_14_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_291;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux_nl = MUX_s_1_2_2(ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_31_3,
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_288_nl, and_dcpl_1236);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_135_nl = act_regs_data_0_1_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_291;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux_1_nl = MUX_s_1_2_2(ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_31_3,
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_135_nl, and_dcpl_1236);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_276_nl = act_regs_data_0_13_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_291;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux_2_nl = MUX_s_1_2_2(ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_31_3,
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_276_nl, and_dcpl_1236);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_300_nl = act_regs_data_0_15_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_291;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux_3_nl = MUX_s_1_2_2(ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_31_3,
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_300_nl, and_dcpl_1236);
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux_4_nl = MUX_v_5_2_2(ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_30_26_2,
      act_regs_data_0_15_sva_dfm_2_30_26, and_dcpl_1236);
  assign not_8882_nl = ~ or_dcpl;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_264_nl = act_regs_data_0_12_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_291;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux_5_nl = MUX_s_1_2_2(ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_31_3,
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_264_nl, and_dcpl_1236);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_147_nl = act_regs_data_0_2_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_291;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux_6_nl = MUX_s_1_2_2(ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_31_3,
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_147_nl, and_dcpl_1236);
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux_7_nl = MUX_v_5_2_2(ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_30_26_2,
      act_regs_data_0_2_sva_dfm_2_30_26, and_dcpl_1236);
  assign not_8883_nl = ~ or_dcpl;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_252_nl = act_regs_data_0_11_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_291;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux_8_nl = MUX_s_1_2_2(ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_31_3,
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_252_nl, and_dcpl_1236);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_159_nl = act_regs_data_0_3_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_291;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux_9_nl = MUX_s_1_2_2(ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_31_3,
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_159_nl, and_dcpl_1236);
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux_10_nl = MUX_v_5_2_2(ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_30_26_2,
      act_regs_data_0_3_sva_dfm_2_30_26, and_dcpl_1236);
  assign not_8884_nl = ~ or_dcpl;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_240_nl = act_regs_data_0_10_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_291;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux_11_nl = MUX_s_1_2_2(ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_31_3,
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_240_nl, and_dcpl_1236);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_171_nl = act_regs_data_0_4_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_291;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux_12_nl = MUX_s_1_2_2(ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_31_3,
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_171_nl, and_dcpl_1236);
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux_13_nl = MUX_v_5_2_2(ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_30_26_2,
      act_regs_data_0_4_sva_dfm_2_30_26, and_dcpl_1236);
  assign not_8885_nl = ~ or_dcpl;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_216_nl = act_regs_data_0_8_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_291;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux_14_nl = MUX_s_1_2_2(ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_31_3,
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_216_nl, and_dcpl_1236);
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux_15_nl = MUX_v_5_2_2(ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_30_26_2,
      act_regs_data_0_8_sva_dfm_2_30_26, and_dcpl_1236);
  assign not_8886_nl = ~ or_dcpl;
  assign ActUnit_PushOutput_if_for_i_mux_nl = MUX_s_1_2_2(ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_25_22_mx0w2_3,
      act_regs_data_0_8_sva_dfm_2_25_22_rsp_0, and_dcpl_1236);
  assign ActUnit_PushOutput_if_for_i_mux_1_nl = MUX_v_3_2_2(ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_25_22_mx0w2_2_0,
      act_regs_data_0_8_sva_dfm_2_25_22_rsp_1, and_dcpl_1236);
  assign not_8896_nl = ~ or_dcpl;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_183_nl = act_regs_data_0_5_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_291;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux_16_nl = MUX_s_1_2_2(ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_31_3,
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_183_nl, and_dcpl_1236);
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux_17_nl = MUX_v_5_2_2(ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_30_26_2,
      act_regs_data_0_5_sva_dfm_2_30_26, and_dcpl_1236);
  assign not_8888_nl = ~ or_dcpl;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_207_nl = act_regs_data_0_7_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_291;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux_18_nl = MUX_s_1_2_2(ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_31_3,
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_207_nl, and_dcpl_1236);
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux_19_nl = MUX_v_5_2_2(ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_30_26_2,
      act_regs_data_0_7_sva_dfm_2_30_26, and_dcpl_1236);
  assign not_8889_nl = ~ or_dcpl;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_195_nl = act_regs_data_0_6_sva_dfm_2_31
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_291;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux_20_nl = MUX_s_1_2_2(ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_31_3,
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_195_nl, and_dcpl_1236);
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux_21_nl = MUX_v_5_2_2(ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_30_26_2,
      act_regs_data_0_6_sva_dfm_2_30_26, and_dcpl_1236);
  assign not_8890_nl = ~ or_dcpl;
  assign while_while_mux1h_150_nl = MUX1HOT_s_1_6_2(reg_act_regs_data_0_0_ftd, (ActUnit_RunInst_case_3_act_port_reg_data_sva[31]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_1_lpi_1_dfm_1_ftd, Silu_for_y_1_lpi_1_dfm_4_31, Gelu_for_y_1_lpi_1_dfm_4_31_1,
      {while_nand_64_ssc_1 , ActUnit_RunInst_switch_lp_and_704_ssc_1 , ActUnit_RunInst_switch_lp_and_65_ssc_1
      , ActUnit_RunInst_switch_lp_and_67_ssc_1 , ActUnit_RunInst_switch_lp_and_71_ssc_1
      , ActUnit_RunInst_switch_lp_and_73_ssc_1});
  assign while_and_213_nl = while_while_mux1h_150_nl & (~ ActUnit_RunInst_switch_lp_and_69_ssc_1);
  assign while_while_mux1h_153_nl = MUX1HOT_s_1_6_2(reg_act_regs_data_0_1_ftd, (ActUnit_RunInst_case_3_act_port_reg_data_sva[63]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_2_lpi_1_dfm_1_ftd, Silu_for_y_2_lpi_1_dfm_4_31, Gelu_for_y_2_lpi_1_dfm_4_31_1,
      {while_nand_64_ssc_1 , ActUnit_RunInst_switch_lp_and_704_ssc_1 , ActUnit_RunInst_switch_lp_and_65_ssc_1
      , ActUnit_RunInst_switch_lp_and_67_ssc_1 , ActUnit_RunInst_switch_lp_and_71_ssc_1
      , ActUnit_RunInst_switch_lp_and_73_ssc_1});
  assign while_and_214_nl = while_while_mux1h_153_nl & (~ ActUnit_RunInst_switch_lp_and_69_ssc_1);
  assign while_while_mux1h_156_nl = MUX1HOT_s_1_6_2(act_regs_data_0_2_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[95]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_3_lpi_1_dfm_1_ftd, Silu_for_y_3_lpi_1_dfm_4_31, Gelu_for_y_3_lpi_1_dfm_4_31_1,
      {while_nand_64_ssc_1 , ActUnit_RunInst_switch_lp_and_704_ssc_1 , ActUnit_RunInst_switch_lp_and_65_ssc_1
      , ActUnit_RunInst_switch_lp_and_67_ssc_1 , ActUnit_RunInst_switch_lp_and_71_ssc_1
      , ActUnit_RunInst_switch_lp_and_73_ssc_1});
  assign while_and_215_nl = while_while_mux1h_156_nl & (~ ActUnit_RunInst_switch_lp_and_69_ssc_1);
  assign while_while_mux1h_159_nl = MUX1HOT_s_1_6_2(act_regs_data_0_3_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[127]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_4_lpi_1_dfm_1_ftd, Silu_for_y_4_lpi_1_dfm_4_31, Gelu_for_y_4_lpi_1_dfm_4_31_1,
      {while_nand_64_ssc_1 , ActUnit_RunInst_switch_lp_and_704_ssc_1 , ActUnit_RunInst_switch_lp_and_65_ssc_1
      , ActUnit_RunInst_switch_lp_and_67_ssc_1 , ActUnit_RunInst_switch_lp_and_71_ssc_1
      , ActUnit_RunInst_switch_lp_and_73_ssc_1});
  assign while_and_216_nl = while_while_mux1h_159_nl & (~ ActUnit_RunInst_switch_lp_and_69_ssc_1);
  assign while_while_mux1h_162_nl = MUX1HOT_s_1_6_2(act_regs_data_0_4_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[159]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_5_lpi_1_dfm_1_ftd, Silu_for_y_5_lpi_1_dfm_4_31, Gelu_for_y_5_lpi_1_dfm_4_31_1,
      {while_nand_64_ssc_1 , ActUnit_RunInst_switch_lp_and_704_ssc_1 , ActUnit_RunInst_switch_lp_and_65_ssc_1
      , ActUnit_RunInst_switch_lp_and_67_ssc_1 , ActUnit_RunInst_switch_lp_and_71_ssc_1
      , ActUnit_RunInst_switch_lp_and_73_ssc_1});
  assign while_and_217_nl = while_while_mux1h_162_nl & (~ ActUnit_RunInst_switch_lp_and_69_ssc_1);
  assign while_while_mux1h_165_nl = MUX1HOT_s_1_6_2(act_regs_data_0_5_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[191]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_6_lpi_1_dfm_1_ftd, Silu_for_y_6_lpi_1_dfm_4_31, Gelu_for_y_6_lpi_1_dfm_4_31_1,
      {while_nand_64_ssc_1 , ActUnit_RunInst_switch_lp_and_704_ssc_1 , ActUnit_RunInst_switch_lp_and_65_ssc_1
      , ActUnit_RunInst_switch_lp_and_67_ssc_1 , ActUnit_RunInst_switch_lp_and_71_ssc_1
      , ActUnit_RunInst_switch_lp_and_73_ssc_1});
  assign while_and_218_nl = while_while_mux1h_165_nl & (~ ActUnit_RunInst_switch_lp_and_69_ssc_1);
  assign while_while_mux1h_168_nl = MUX1HOT_s_1_6_2(act_regs_data_0_6_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[223]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_7_lpi_1_dfm_1_ftd, Silu_for_y_7_lpi_1_dfm_4_31, Gelu_for_y_7_lpi_1_dfm_4_31_1,
      {while_nand_64_ssc_1 , ActUnit_RunInst_switch_lp_and_704_ssc_1 , ActUnit_RunInst_switch_lp_and_65_ssc_1
      , ActUnit_RunInst_switch_lp_and_67_ssc_1 , ActUnit_RunInst_switch_lp_and_71_ssc_1
      , ActUnit_RunInst_switch_lp_and_73_ssc_1});
  assign while_and_219_nl = while_while_mux1h_168_nl & (~ ActUnit_RunInst_switch_lp_and_69_ssc_1);
  assign while_while_mux1h_171_nl = MUX1HOT_s_1_6_2(act_regs_data_0_7_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[255]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_8_lpi_1_dfm_1_ftd, Silu_for_y_8_lpi_1_dfm_4_31, Gelu_for_y_8_lpi_1_dfm_4_31_1,
      {while_nand_64_ssc_1 , ActUnit_RunInst_switch_lp_and_704_ssc_1 , ActUnit_RunInst_switch_lp_and_65_ssc_1
      , ActUnit_RunInst_switch_lp_and_67_ssc_1 , ActUnit_RunInst_switch_lp_and_71_ssc_1
      , ActUnit_RunInst_switch_lp_and_73_ssc_1});
  assign while_and_220_nl = while_while_mux1h_171_nl & (~ ActUnit_RunInst_switch_lp_and_69_ssc_1);
  assign while_while_mux1h_174_nl = MUX1HOT_s_1_6_2(act_regs_data_0_8_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[287]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_9_lpi_1_dfm_1_ftd, Silu_for_y_9_lpi_1_dfm_4_31_1, Gelu_for_y_9_lpi_1_dfm_4_31_1,
      {while_nand_64_ssc_1 , ActUnit_RunInst_switch_lp_and_704_ssc_1 , ActUnit_RunInst_switch_lp_and_65_ssc_1
      , ActUnit_RunInst_switch_lp_and_67_ssc_1 , ActUnit_RunInst_switch_lp_and_71_ssc_1
      , ActUnit_RunInst_switch_lp_and_73_ssc_1});
  assign while_and_221_nl = while_while_mux1h_174_nl & (~ ActUnit_RunInst_switch_lp_and_69_ssc_1);
  assign while_while_mux1h_177_nl = MUX1HOT_s_1_6_2(act_regs_data_0_9_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[319]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_10_lpi_1_dfm_1_ftd, Silu_for_y_10_lpi_1_dfm_4_31_1, Gelu_for_y_10_lpi_1_dfm_4_31_1,
      {while_nand_64_ssc_1 , ActUnit_RunInst_switch_lp_and_704_ssc_1 , ActUnit_RunInst_switch_lp_and_65_ssc_1
      , ActUnit_RunInst_switch_lp_and_67_ssc_1 , ActUnit_RunInst_switch_lp_and_71_ssc_1
      , ActUnit_RunInst_switch_lp_and_73_ssc_1});
  assign while_and_222_nl = while_while_mux1h_177_nl & (~ ActUnit_RunInst_switch_lp_and_69_ssc_1);
  assign while_while_mux1h_180_nl = MUX1HOT_s_1_6_2(reg_act_regs_data_0_10_ftd, (ActUnit_RunInst_case_3_act_port_reg_data_sva[351]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_11_lpi_1_dfm_1_ftd, Silu_for_y_11_lpi_1_dfm_4_31_1, Gelu_for_y_11_lpi_1_dfm_4_31_1,
      {while_nand_64_ssc_1 , ActUnit_RunInst_switch_lp_and_704_ssc_1 , ActUnit_RunInst_switch_lp_and_65_ssc_1
      , ActUnit_RunInst_switch_lp_and_67_ssc_1 , ActUnit_RunInst_switch_lp_and_71_ssc_1
      , ActUnit_RunInst_switch_lp_and_73_ssc_1});
  assign while_and_223_nl = while_while_mux1h_180_nl & (~ ActUnit_RunInst_switch_lp_and_69_ssc_1);
  assign while_while_mux1h_183_nl = MUX1HOT_s_1_6_2(reg_act_regs_data_0_11_ftd, (ActUnit_RunInst_case_3_act_port_reg_data_sva[383]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_12_lpi_1_dfm_1_ftd, Silu_for_y_12_lpi_1_dfm_4_31_1, Gelu_for_y_12_lpi_1_dfm_4_31_1,
      {while_nand_64_ssc_1 , ActUnit_RunInst_switch_lp_and_704_ssc_1 , ActUnit_RunInst_switch_lp_and_65_ssc_1
      , ActUnit_RunInst_switch_lp_and_67_ssc_1 , ActUnit_RunInst_switch_lp_and_71_ssc_1
      , ActUnit_RunInst_switch_lp_and_73_ssc_1});
  assign while_and_224_nl = while_while_mux1h_183_nl & (~ ActUnit_RunInst_switch_lp_and_69_ssc_1);
  assign while_while_mux1h_186_nl = MUX1HOT_s_1_6_2(reg_act_regs_data_0_12_ftd, (ActUnit_RunInst_case_3_act_port_reg_data_sva[415]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_13_lpi_1_dfm_1_ftd, Silu_for_y_13_lpi_1_dfm_4_31_1, Gelu_for_y_13_lpi_1_dfm_4_31_1,
      {while_nand_64_ssc_1 , ActUnit_RunInst_switch_lp_and_704_ssc_1 , ActUnit_RunInst_switch_lp_and_65_ssc_1
      , ActUnit_RunInst_switch_lp_and_67_ssc_1 , ActUnit_RunInst_switch_lp_and_71_ssc_1
      , ActUnit_RunInst_switch_lp_and_73_ssc_1});
  assign while_and_225_nl = while_while_mux1h_186_nl & (~ ActUnit_RunInst_switch_lp_and_69_ssc_1);
  assign while_while_mux1h_189_nl = MUX1HOT_s_1_6_2(reg_act_regs_data_0_13_ftd, (ActUnit_RunInst_case_3_act_port_reg_data_sva[447]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_14_lpi_1_dfm_1_ftd, Silu_for_y_14_lpi_1_dfm_4_31_1, Gelu_for_y_14_lpi_1_dfm_4_31_1,
      {while_nand_64_ssc_1 , ActUnit_RunInst_switch_lp_and_704_ssc_1 , ActUnit_RunInst_switch_lp_and_65_ssc_1
      , ActUnit_RunInst_switch_lp_and_67_ssc_1 , ActUnit_RunInst_switch_lp_and_71_ssc_1
      , ActUnit_RunInst_switch_lp_and_73_ssc_1});
  assign while_and_226_nl = while_while_mux1h_189_nl & (~ ActUnit_RunInst_switch_lp_and_69_ssc_1);
  assign while_while_mux1h_192_nl = MUX1HOT_s_1_6_2(act_regs_data_0_14_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[479]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_15_lpi_1_dfm_1_ftd, Silu_for_y_15_lpi_1_dfm_4_31_1, Gelu_for_y_15_lpi_1_dfm_4_31_1,
      {while_nand_64_ssc_1 , ActUnit_RunInst_switch_lp_and_704_ssc_1 , ActUnit_RunInst_switch_lp_and_65_ssc_1
      , ActUnit_RunInst_switch_lp_and_67_ssc_1 , ActUnit_RunInst_switch_lp_and_71_ssc_1
      , ActUnit_RunInst_switch_lp_and_73_ssc_1});
  assign while_and_227_nl = while_while_mux1h_192_nl & (~ ActUnit_RunInst_switch_lp_and_69_ssc_1);
  assign while_while_mux1h_195_nl = MUX1HOT_s_1_6_2(act_regs_data_0_15_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[511]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_lpi_1_dfm_1_ftd, Silu_for_y_lpi_1_dfm_4_31_1, Gelu_for_y_lpi_1_dfm_4_31_1,
      {while_nand_64_ssc_1 , ActUnit_RunInst_switch_lp_and_704_ssc_1 , ActUnit_RunInst_switch_lp_and_65_ssc_1
      , ActUnit_RunInst_switch_lp_and_67_ssc_1 , ActUnit_RunInst_switch_lp_and_71_ssc_1
      , ActUnit_RunInst_switch_lp_and_73_ssc_1});
  assign while_and_228_nl = while_while_mux1h_195_nl & (~ ActUnit_RunInst_switch_lp_and_69_ssc_1);
  assign while_while_mux1h_198_nl = MUX1HOT_s_1_6_2(act_regs_data_1_0_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[31]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_1_lpi_1_dfm_1_ftd, Silu_for_y_1_lpi_1_dfm_4_31, Gelu_for_y_1_lpi_1_dfm_4_31_1,
      {while_nand_80_ssc_1 , ActUnit_RunInst_switch_lp_and_737_ssc_1 , ActUnit_RunInst_switch_lp_and_225_ssc_1
      , ActUnit_RunInst_switch_lp_and_227_ssc_1 , ActUnit_RunInst_switch_lp_and_231_ssc_1
      , ActUnit_RunInst_switch_lp_and_233_ssc_1});
  assign while_and_229_nl = while_while_mux1h_198_nl & (~ ActUnit_RunInst_switch_lp_and_229_ssc_1);
  assign while_while_mux1h_201_nl = MUX1HOT_s_1_6_2(act_regs_data_1_1_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[63]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_2_lpi_1_dfm_1_ftd, Silu_for_y_2_lpi_1_dfm_4_31, Gelu_for_y_2_lpi_1_dfm_4_31_1,
      {while_nand_80_ssc_1 , ActUnit_RunInst_switch_lp_and_737_ssc_1 , ActUnit_RunInst_switch_lp_and_225_ssc_1
      , ActUnit_RunInst_switch_lp_and_227_ssc_1 , ActUnit_RunInst_switch_lp_and_231_ssc_1
      , ActUnit_RunInst_switch_lp_and_233_ssc_1});
  assign while_and_230_nl = while_while_mux1h_201_nl & (~ ActUnit_RunInst_switch_lp_and_229_ssc_1);
  assign while_while_mux1h_204_nl = MUX1HOT_s_1_6_2(act_regs_data_1_2_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[95]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_3_lpi_1_dfm_1_ftd, Silu_for_y_3_lpi_1_dfm_4_31, Gelu_for_y_3_lpi_1_dfm_4_31_1,
      {while_nand_80_ssc_1 , ActUnit_RunInst_switch_lp_and_737_ssc_1 , ActUnit_RunInst_switch_lp_and_225_ssc_1
      , ActUnit_RunInst_switch_lp_and_227_ssc_1 , ActUnit_RunInst_switch_lp_and_231_ssc_1
      , ActUnit_RunInst_switch_lp_and_233_ssc_1});
  assign while_and_231_nl = while_while_mux1h_204_nl & (~ ActUnit_RunInst_switch_lp_and_229_ssc_1);
  assign while_while_mux1h_207_nl = MUX1HOT_s_1_6_2(act_regs_data_1_3_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[127]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_4_lpi_1_dfm_1_ftd, Silu_for_y_4_lpi_1_dfm_4_31, Gelu_for_y_4_lpi_1_dfm_4_31_1,
      {while_nand_80_ssc_1 , ActUnit_RunInst_switch_lp_and_737_ssc_1 , ActUnit_RunInst_switch_lp_and_225_ssc_1
      , ActUnit_RunInst_switch_lp_and_227_ssc_1 , ActUnit_RunInst_switch_lp_and_231_ssc_1
      , ActUnit_RunInst_switch_lp_and_233_ssc_1});
  assign while_and_232_nl = while_while_mux1h_207_nl & (~ ActUnit_RunInst_switch_lp_and_229_ssc_1);
  assign while_while_mux1h_210_nl = MUX1HOT_s_1_6_2(act_regs_data_1_4_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[159]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_5_lpi_1_dfm_1_ftd, Silu_for_y_5_lpi_1_dfm_4_31, Gelu_for_y_5_lpi_1_dfm_4_31_1,
      {while_nand_80_ssc_1 , ActUnit_RunInst_switch_lp_and_737_ssc_1 , ActUnit_RunInst_switch_lp_and_225_ssc_1
      , ActUnit_RunInst_switch_lp_and_227_ssc_1 , ActUnit_RunInst_switch_lp_and_231_ssc_1
      , ActUnit_RunInst_switch_lp_and_233_ssc_1});
  assign while_and_233_nl = while_while_mux1h_210_nl & (~ ActUnit_RunInst_switch_lp_and_229_ssc_1);
  assign while_while_mux1h_213_nl = MUX1HOT_s_1_6_2(act_regs_data_1_5_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[191]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_6_lpi_1_dfm_1_ftd, Silu_for_y_6_lpi_1_dfm_4_31, Gelu_for_y_6_lpi_1_dfm_4_31_1,
      {while_nand_80_ssc_1 , ActUnit_RunInst_switch_lp_and_737_ssc_1 , ActUnit_RunInst_switch_lp_and_225_ssc_1
      , ActUnit_RunInst_switch_lp_and_227_ssc_1 , ActUnit_RunInst_switch_lp_and_231_ssc_1
      , ActUnit_RunInst_switch_lp_and_233_ssc_1});
  assign while_and_234_nl = while_while_mux1h_213_nl & (~ ActUnit_RunInst_switch_lp_and_229_ssc_1);
  assign while_while_mux1h_216_nl = MUX1HOT_s_1_6_2(act_regs_data_1_6_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[223]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_7_lpi_1_dfm_1_ftd, Silu_for_y_7_lpi_1_dfm_4_31, Gelu_for_y_7_lpi_1_dfm_4_31_1,
      {while_nand_80_ssc_1 , ActUnit_RunInst_switch_lp_and_737_ssc_1 , ActUnit_RunInst_switch_lp_and_225_ssc_1
      , ActUnit_RunInst_switch_lp_and_227_ssc_1 , ActUnit_RunInst_switch_lp_and_231_ssc_1
      , ActUnit_RunInst_switch_lp_and_233_ssc_1});
  assign while_and_235_nl = while_while_mux1h_216_nl & (~ ActUnit_RunInst_switch_lp_and_229_ssc_1);
  assign while_while_mux1h_219_nl = MUX1HOT_s_1_6_2(act_regs_data_1_7_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[255]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_8_lpi_1_dfm_1_ftd, Silu_for_y_8_lpi_1_dfm_4_31, Gelu_for_y_8_lpi_1_dfm_4_31_1,
      {while_nand_80_ssc_1 , ActUnit_RunInst_switch_lp_and_737_ssc_1 , ActUnit_RunInst_switch_lp_and_225_ssc_1
      , ActUnit_RunInst_switch_lp_and_227_ssc_1 , ActUnit_RunInst_switch_lp_and_231_ssc_1
      , ActUnit_RunInst_switch_lp_and_233_ssc_1});
  assign while_and_236_nl = while_while_mux1h_219_nl & (~ ActUnit_RunInst_switch_lp_and_229_ssc_1);
  assign while_while_mux1h_222_nl = MUX1HOT_s_1_6_2(act_regs_data_1_8_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[287]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_9_lpi_1_dfm_1_ftd, Silu_for_y_9_lpi_1_dfm_4_31_1, Gelu_for_y_9_lpi_1_dfm_4_31_1,
      {while_nand_80_ssc_1 , ActUnit_RunInst_switch_lp_and_737_ssc_1 , ActUnit_RunInst_switch_lp_and_225_ssc_1
      , ActUnit_RunInst_switch_lp_and_227_ssc_1 , ActUnit_RunInst_switch_lp_and_231_ssc_1
      , ActUnit_RunInst_switch_lp_and_233_ssc_1});
  assign while_and_237_nl = while_while_mux1h_222_nl & (~ ActUnit_RunInst_switch_lp_and_229_ssc_1);
  assign while_while_mux1h_225_nl = MUX1HOT_s_1_6_2(act_regs_data_1_9_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[319]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_10_lpi_1_dfm_1_ftd, Silu_for_y_10_lpi_1_dfm_4_31_1, Gelu_for_y_10_lpi_1_dfm_4_31_1,
      {while_nand_80_ssc_1 , ActUnit_RunInst_switch_lp_and_737_ssc_1 , ActUnit_RunInst_switch_lp_and_225_ssc_1
      , ActUnit_RunInst_switch_lp_and_227_ssc_1 , ActUnit_RunInst_switch_lp_and_231_ssc_1
      , ActUnit_RunInst_switch_lp_and_233_ssc_1});
  assign while_and_238_nl = while_while_mux1h_225_nl & (~ ActUnit_RunInst_switch_lp_and_229_ssc_1);
  assign while_while_mux1h_228_nl = MUX1HOT_s_1_6_2(act_regs_data_1_10_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[351]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_11_lpi_1_dfm_1_ftd, Silu_for_y_11_lpi_1_dfm_4_31_1, Gelu_for_y_11_lpi_1_dfm_4_31_1,
      {while_nand_80_ssc_1 , ActUnit_RunInst_switch_lp_and_737_ssc_1 , ActUnit_RunInst_switch_lp_and_225_ssc_1
      , ActUnit_RunInst_switch_lp_and_227_ssc_1 , ActUnit_RunInst_switch_lp_and_231_ssc_1
      , ActUnit_RunInst_switch_lp_and_233_ssc_1});
  assign while_and_239_nl = while_while_mux1h_228_nl & (~ ActUnit_RunInst_switch_lp_and_229_ssc_1);
  assign while_while_mux1h_231_nl = MUX1HOT_s_1_6_2(act_regs_data_1_11_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[383]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_12_lpi_1_dfm_1_ftd, Silu_for_y_12_lpi_1_dfm_4_31_1, Gelu_for_y_12_lpi_1_dfm_4_31_1,
      {while_nand_80_ssc_1 , ActUnit_RunInst_switch_lp_and_737_ssc_1 , ActUnit_RunInst_switch_lp_and_225_ssc_1
      , ActUnit_RunInst_switch_lp_and_227_ssc_1 , ActUnit_RunInst_switch_lp_and_231_ssc_1
      , ActUnit_RunInst_switch_lp_and_233_ssc_1});
  assign while_and_240_nl = while_while_mux1h_231_nl & (~ ActUnit_RunInst_switch_lp_and_229_ssc_1);
  assign while_while_mux1h_234_nl = MUX1HOT_s_1_6_2(act_regs_data_1_12_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[415]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_13_lpi_1_dfm_1_ftd, Silu_for_y_13_lpi_1_dfm_4_31_1, Gelu_for_y_13_lpi_1_dfm_4_31_1,
      {while_nand_80_ssc_1 , ActUnit_RunInst_switch_lp_and_737_ssc_1 , ActUnit_RunInst_switch_lp_and_225_ssc_1
      , ActUnit_RunInst_switch_lp_and_227_ssc_1 , ActUnit_RunInst_switch_lp_and_231_ssc_1
      , ActUnit_RunInst_switch_lp_and_233_ssc_1});
  assign while_and_241_nl = while_while_mux1h_234_nl & (~ ActUnit_RunInst_switch_lp_and_229_ssc_1);
  assign while_while_mux1h_237_nl = MUX1HOT_s_1_6_2(act_regs_data_1_13_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[447]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_14_lpi_1_dfm_1_ftd, Silu_for_y_14_lpi_1_dfm_4_31_1, Gelu_for_y_14_lpi_1_dfm_4_31_1,
      {while_nand_80_ssc_1 , ActUnit_RunInst_switch_lp_and_737_ssc_1 , ActUnit_RunInst_switch_lp_and_225_ssc_1
      , ActUnit_RunInst_switch_lp_and_227_ssc_1 , ActUnit_RunInst_switch_lp_and_231_ssc_1
      , ActUnit_RunInst_switch_lp_and_233_ssc_1});
  assign while_and_242_nl = while_while_mux1h_237_nl & (~ ActUnit_RunInst_switch_lp_and_229_ssc_1);
  assign while_while_mux1h_240_nl = MUX1HOT_s_1_6_2(act_regs_data_1_14_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[479]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_15_lpi_1_dfm_1_ftd, Silu_for_y_15_lpi_1_dfm_4_31_1, Gelu_for_y_15_lpi_1_dfm_4_31_1,
      {while_nand_80_ssc_1 , ActUnit_RunInst_switch_lp_and_737_ssc_1 , ActUnit_RunInst_switch_lp_and_225_ssc_1
      , ActUnit_RunInst_switch_lp_and_227_ssc_1 , ActUnit_RunInst_switch_lp_and_231_ssc_1
      , ActUnit_RunInst_switch_lp_and_233_ssc_1});
  assign while_and_243_nl = while_while_mux1h_240_nl & (~ ActUnit_RunInst_switch_lp_and_229_ssc_1);
  assign while_while_mux1h_243_nl = MUX1HOT_s_1_6_2(act_regs_data_1_15_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[511]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_lpi_1_dfm_1_ftd, Silu_for_y_lpi_1_dfm_4_31_1, Gelu_for_y_lpi_1_dfm_4_31_1,
      {while_nand_80_ssc_1 , ActUnit_RunInst_switch_lp_and_737_ssc_1 , ActUnit_RunInst_switch_lp_and_225_ssc_1
      , ActUnit_RunInst_switch_lp_and_227_ssc_1 , ActUnit_RunInst_switch_lp_and_231_ssc_1
      , ActUnit_RunInst_switch_lp_and_233_ssc_1});
  assign while_and_244_nl = while_while_mux1h_243_nl & (~ ActUnit_RunInst_switch_lp_and_229_ssc_1);
  assign while_while_mux1h_246_nl = MUX1HOT_s_1_6_2(act_regs_data_2_0_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[31]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_1_lpi_1_dfm_1_ftd, Silu_for_y_1_lpi_1_dfm_4_31, Gelu_for_y_1_lpi_1_dfm_4_31_1,
      {while_nand_96_ssc_1 , ActUnit_RunInst_switch_lp_and_769_ssc_1 , ActUnit_RunInst_switch_lp_and_385_ssc_1
      , ActUnit_RunInst_switch_lp_and_387_ssc_1 , ActUnit_RunInst_switch_lp_and_391_ssc_1
      , ActUnit_RunInst_switch_lp_and_393_ssc_1});
  assign while_and_245_nl = while_while_mux1h_246_nl & (~ ActUnit_RunInst_switch_lp_and_389_ssc_1);
  assign while_while_mux1h_249_nl = MUX1HOT_s_1_6_2(act_regs_data_2_1_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[63]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_2_lpi_1_dfm_1_ftd, Silu_for_y_2_lpi_1_dfm_4_31, Gelu_for_y_2_lpi_1_dfm_4_31_1,
      {while_nand_96_ssc_1 , ActUnit_RunInst_switch_lp_and_769_ssc_1 , ActUnit_RunInst_switch_lp_and_385_ssc_1
      , ActUnit_RunInst_switch_lp_and_387_ssc_1 , ActUnit_RunInst_switch_lp_and_391_ssc_1
      , ActUnit_RunInst_switch_lp_and_393_ssc_1});
  assign while_and_246_nl = while_while_mux1h_249_nl & (~ ActUnit_RunInst_switch_lp_and_389_ssc_1);
  assign while_while_mux1h_252_nl = MUX1HOT_s_1_6_2(act_regs_data_2_2_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[95]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_3_lpi_1_dfm_1_ftd, Silu_for_y_3_lpi_1_dfm_4_31, Gelu_for_y_3_lpi_1_dfm_4_31_1,
      {while_nand_96_ssc_1 , ActUnit_RunInst_switch_lp_and_769_ssc_1 , ActUnit_RunInst_switch_lp_and_385_ssc_1
      , ActUnit_RunInst_switch_lp_and_387_ssc_1 , ActUnit_RunInst_switch_lp_and_391_ssc_1
      , ActUnit_RunInst_switch_lp_and_393_ssc_1});
  assign while_and_247_nl = while_while_mux1h_252_nl & (~ ActUnit_RunInst_switch_lp_and_389_ssc_1);
  assign while_while_mux1h_255_nl = MUX1HOT_s_1_6_2(act_regs_data_2_3_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[127]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_4_lpi_1_dfm_1_ftd, Silu_for_y_4_lpi_1_dfm_4_31, Gelu_for_y_4_lpi_1_dfm_4_31_1,
      {while_nand_96_ssc_1 , ActUnit_RunInst_switch_lp_and_769_ssc_1 , ActUnit_RunInst_switch_lp_and_385_ssc_1
      , ActUnit_RunInst_switch_lp_and_387_ssc_1 , ActUnit_RunInst_switch_lp_and_391_ssc_1
      , ActUnit_RunInst_switch_lp_and_393_ssc_1});
  assign while_and_248_nl = while_while_mux1h_255_nl & (~ ActUnit_RunInst_switch_lp_and_389_ssc_1);
  assign while_while_mux1h_258_nl = MUX1HOT_s_1_6_2(act_regs_data_2_4_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[159]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_5_lpi_1_dfm_1_ftd, Silu_for_y_5_lpi_1_dfm_4_31, Gelu_for_y_5_lpi_1_dfm_4_31_1,
      {while_nand_96_ssc_1 , ActUnit_RunInst_switch_lp_and_769_ssc_1 , ActUnit_RunInst_switch_lp_and_385_ssc_1
      , ActUnit_RunInst_switch_lp_and_387_ssc_1 , ActUnit_RunInst_switch_lp_and_391_ssc_1
      , ActUnit_RunInst_switch_lp_and_393_ssc_1});
  assign while_and_249_nl = while_while_mux1h_258_nl & (~ ActUnit_RunInst_switch_lp_and_389_ssc_1);
  assign while_while_mux1h_261_nl = MUX1HOT_s_1_6_2(act_regs_data_2_5_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[191]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_6_lpi_1_dfm_1_ftd, Silu_for_y_6_lpi_1_dfm_4_31, Gelu_for_y_6_lpi_1_dfm_4_31_1,
      {while_nand_96_ssc_1 , ActUnit_RunInst_switch_lp_and_769_ssc_1 , ActUnit_RunInst_switch_lp_and_385_ssc_1
      , ActUnit_RunInst_switch_lp_and_387_ssc_1 , ActUnit_RunInst_switch_lp_and_391_ssc_1
      , ActUnit_RunInst_switch_lp_and_393_ssc_1});
  assign while_and_250_nl = while_while_mux1h_261_nl & (~ ActUnit_RunInst_switch_lp_and_389_ssc_1);
  assign while_while_mux1h_264_nl = MUX1HOT_s_1_6_2(act_regs_data_2_6_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[223]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_7_lpi_1_dfm_1_ftd, Silu_for_y_7_lpi_1_dfm_4_31, Gelu_for_y_7_lpi_1_dfm_4_31_1,
      {while_nand_96_ssc_1 , ActUnit_RunInst_switch_lp_and_769_ssc_1 , ActUnit_RunInst_switch_lp_and_385_ssc_1
      , ActUnit_RunInst_switch_lp_and_387_ssc_1 , ActUnit_RunInst_switch_lp_and_391_ssc_1
      , ActUnit_RunInst_switch_lp_and_393_ssc_1});
  assign while_and_251_nl = while_while_mux1h_264_nl & (~ ActUnit_RunInst_switch_lp_and_389_ssc_1);
  assign while_while_mux1h_267_nl = MUX1HOT_s_1_6_2(act_regs_data_2_7_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[255]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_8_lpi_1_dfm_1_ftd, Silu_for_y_8_lpi_1_dfm_4_31, Gelu_for_y_8_lpi_1_dfm_4_31_1,
      {while_nand_96_ssc_1 , ActUnit_RunInst_switch_lp_and_769_ssc_1 , ActUnit_RunInst_switch_lp_and_385_ssc_1
      , ActUnit_RunInst_switch_lp_and_387_ssc_1 , ActUnit_RunInst_switch_lp_and_391_ssc_1
      , ActUnit_RunInst_switch_lp_and_393_ssc_1});
  assign while_and_252_nl = while_while_mux1h_267_nl & (~ ActUnit_RunInst_switch_lp_and_389_ssc_1);
  assign while_while_mux1h_270_nl = MUX1HOT_s_1_6_2(act_regs_data_2_8_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[287]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_9_lpi_1_dfm_1_ftd, Silu_for_y_9_lpi_1_dfm_4_31_1, Gelu_for_y_9_lpi_1_dfm_4_31_1,
      {while_nand_96_ssc_1 , ActUnit_RunInst_switch_lp_and_769_ssc_1 , ActUnit_RunInst_switch_lp_and_385_ssc_1
      , ActUnit_RunInst_switch_lp_and_387_ssc_1 , ActUnit_RunInst_switch_lp_and_391_ssc_1
      , ActUnit_RunInst_switch_lp_and_393_ssc_1});
  assign while_and_253_nl = while_while_mux1h_270_nl & (~ ActUnit_RunInst_switch_lp_and_389_ssc_1);
  assign while_while_mux1h_273_nl = MUX1HOT_s_1_6_2(act_regs_data_2_9_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[319]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_10_lpi_1_dfm_1_ftd, Silu_for_y_10_lpi_1_dfm_4_31_1, Gelu_for_y_10_lpi_1_dfm_4_31_1,
      {while_nand_96_ssc_1 , ActUnit_RunInst_switch_lp_and_769_ssc_1 , ActUnit_RunInst_switch_lp_and_385_ssc_1
      , ActUnit_RunInst_switch_lp_and_387_ssc_1 , ActUnit_RunInst_switch_lp_and_391_ssc_1
      , ActUnit_RunInst_switch_lp_and_393_ssc_1});
  assign while_and_254_nl = while_while_mux1h_273_nl & (~ ActUnit_RunInst_switch_lp_and_389_ssc_1);
  assign while_while_mux1h_276_nl = MUX1HOT_s_1_6_2(act_regs_data_2_10_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[351]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_11_lpi_1_dfm_1_ftd, Silu_for_y_11_lpi_1_dfm_4_31_1, Gelu_for_y_11_lpi_1_dfm_4_31_1,
      {while_nand_96_ssc_1 , ActUnit_RunInst_switch_lp_and_769_ssc_1 , ActUnit_RunInst_switch_lp_and_385_ssc_1
      , ActUnit_RunInst_switch_lp_and_387_ssc_1 , ActUnit_RunInst_switch_lp_and_391_ssc_1
      , ActUnit_RunInst_switch_lp_and_393_ssc_1});
  assign while_and_255_nl = while_while_mux1h_276_nl & (~ ActUnit_RunInst_switch_lp_and_389_ssc_1);
  assign while_while_mux1h_279_nl = MUX1HOT_s_1_6_2(act_regs_data_2_11_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[383]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_12_lpi_1_dfm_1_ftd, Silu_for_y_12_lpi_1_dfm_4_31_1, Gelu_for_y_12_lpi_1_dfm_4_31_1,
      {while_nand_96_ssc_1 , ActUnit_RunInst_switch_lp_and_769_ssc_1 , ActUnit_RunInst_switch_lp_and_385_ssc_1
      , ActUnit_RunInst_switch_lp_and_387_ssc_1 , ActUnit_RunInst_switch_lp_and_391_ssc_1
      , ActUnit_RunInst_switch_lp_and_393_ssc_1});
  assign while_and_256_nl = while_while_mux1h_279_nl & (~ ActUnit_RunInst_switch_lp_and_389_ssc_1);
  assign while_while_mux1h_282_nl = MUX1HOT_s_1_6_2(act_regs_data_2_12_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[415]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_13_lpi_1_dfm_1_ftd, Silu_for_y_13_lpi_1_dfm_4_31_1, Gelu_for_y_13_lpi_1_dfm_4_31_1,
      {while_nand_96_ssc_1 , ActUnit_RunInst_switch_lp_and_769_ssc_1 , ActUnit_RunInst_switch_lp_and_385_ssc_1
      , ActUnit_RunInst_switch_lp_and_387_ssc_1 , ActUnit_RunInst_switch_lp_and_391_ssc_1
      , ActUnit_RunInst_switch_lp_and_393_ssc_1});
  assign while_and_257_nl = while_while_mux1h_282_nl & (~ ActUnit_RunInst_switch_lp_and_389_ssc_1);
  assign while_while_mux1h_285_nl = MUX1HOT_s_1_6_2(act_regs_data_2_13_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[447]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_14_lpi_1_dfm_1_ftd, Silu_for_y_14_lpi_1_dfm_4_31_1, Gelu_for_y_14_lpi_1_dfm_4_31_1,
      {while_nand_96_ssc_1 , ActUnit_RunInst_switch_lp_and_769_ssc_1 , ActUnit_RunInst_switch_lp_and_385_ssc_1
      , ActUnit_RunInst_switch_lp_and_387_ssc_1 , ActUnit_RunInst_switch_lp_and_391_ssc_1
      , ActUnit_RunInst_switch_lp_and_393_ssc_1});
  assign while_and_258_nl = while_while_mux1h_285_nl & (~ ActUnit_RunInst_switch_lp_and_389_ssc_1);
  assign while_while_mux1h_288_nl = MUX1HOT_s_1_6_2(act_regs_data_2_14_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[479]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_15_lpi_1_dfm_1_ftd, Silu_for_y_15_lpi_1_dfm_4_31_1, Gelu_for_y_15_lpi_1_dfm_4_31_1,
      {while_nand_96_ssc_1 , ActUnit_RunInst_switch_lp_and_769_ssc_1 , ActUnit_RunInst_switch_lp_and_385_ssc_1
      , ActUnit_RunInst_switch_lp_and_387_ssc_1 , ActUnit_RunInst_switch_lp_and_391_ssc_1
      , ActUnit_RunInst_switch_lp_and_393_ssc_1});
  assign while_and_259_nl = while_while_mux1h_288_nl & (~ ActUnit_RunInst_switch_lp_and_389_ssc_1);
  assign while_while_mux1h_291_nl = MUX1HOT_s_1_6_2(act_regs_data_2_15_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[511]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_lpi_1_dfm_1_ftd, Silu_for_y_lpi_1_dfm_4_31_1, Gelu_for_y_lpi_1_dfm_4_31_1,
      {while_nand_96_ssc_1 , ActUnit_RunInst_switch_lp_and_769_ssc_1 , ActUnit_RunInst_switch_lp_and_385_ssc_1
      , ActUnit_RunInst_switch_lp_and_387_ssc_1 , ActUnit_RunInst_switch_lp_and_391_ssc_1
      , ActUnit_RunInst_switch_lp_and_393_ssc_1});
  assign while_and_260_nl = while_while_mux1h_291_nl & (~ ActUnit_RunInst_switch_lp_and_389_ssc_1);
  assign while_while_mux1h_294_nl = MUX1HOT_s_1_6_2(act_regs_data_3_0_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[31]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_1_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_1_lpi_1_dfm_1_ftd, Silu_for_y_1_lpi_1_dfm_4_31, Gelu_for_y_1_lpi_1_dfm_4_31_1,
      {while_nand_112_ssc_1 , ActUnit_RunInst_switch_lp_and_801_ssc_1 , ActUnit_RunInst_switch_lp_and_545_ssc_1
      , ActUnit_RunInst_switch_lp_and_547_ssc_1 , ActUnit_RunInst_switch_lp_and_551_ssc_1
      , ActUnit_RunInst_switch_lp_and_553_ssc_1});
  assign while_and_261_nl = while_while_mux1h_294_nl & (~ ActUnit_RunInst_switch_lp_and_549_ssc_1);
  assign while_while_mux1h_297_nl = MUX1HOT_s_1_6_2(act_regs_data_3_1_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[63]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_2_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_2_lpi_1_dfm_1_ftd, Silu_for_y_2_lpi_1_dfm_4_31, Gelu_for_y_2_lpi_1_dfm_4_31_1,
      {while_nand_112_ssc_1 , ActUnit_RunInst_switch_lp_and_801_ssc_1 , ActUnit_RunInst_switch_lp_and_545_ssc_1
      , ActUnit_RunInst_switch_lp_and_547_ssc_1 , ActUnit_RunInst_switch_lp_and_551_ssc_1
      , ActUnit_RunInst_switch_lp_and_553_ssc_1});
  assign while_and_262_nl = while_while_mux1h_297_nl & (~ ActUnit_RunInst_switch_lp_and_549_ssc_1);
  assign while_while_mux1h_300_nl = MUX1HOT_s_1_6_2(act_regs_data_3_2_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[95]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_3_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_3_lpi_1_dfm_1_ftd, Silu_for_y_3_lpi_1_dfm_4_31, Gelu_for_y_3_lpi_1_dfm_4_31_1,
      {while_nand_112_ssc_1 , ActUnit_RunInst_switch_lp_and_801_ssc_1 , ActUnit_RunInst_switch_lp_and_545_ssc_1
      , ActUnit_RunInst_switch_lp_and_547_ssc_1 , ActUnit_RunInst_switch_lp_and_551_ssc_1
      , ActUnit_RunInst_switch_lp_and_553_ssc_1});
  assign while_and_263_nl = while_while_mux1h_300_nl & (~ ActUnit_RunInst_switch_lp_and_549_ssc_1);
  assign while_while_mux1h_303_nl = MUX1HOT_s_1_6_2(act_regs_data_3_3_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[127]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_4_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_4_lpi_1_dfm_1_ftd, Silu_for_y_4_lpi_1_dfm_4_31, Gelu_for_y_4_lpi_1_dfm_4_31_1,
      {while_nand_112_ssc_1 , ActUnit_RunInst_switch_lp_and_801_ssc_1 , ActUnit_RunInst_switch_lp_and_545_ssc_1
      , ActUnit_RunInst_switch_lp_and_547_ssc_1 , ActUnit_RunInst_switch_lp_and_551_ssc_1
      , ActUnit_RunInst_switch_lp_and_553_ssc_1});
  assign while_and_264_nl = while_while_mux1h_303_nl & (~ ActUnit_RunInst_switch_lp_and_549_ssc_1);
  assign while_while_mux1h_306_nl = MUX1HOT_s_1_6_2(act_regs_data_3_4_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[159]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_5_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_5_lpi_1_dfm_1_ftd, Silu_for_y_5_lpi_1_dfm_4_31, Gelu_for_y_5_lpi_1_dfm_4_31_1,
      {while_nand_112_ssc_1 , ActUnit_RunInst_switch_lp_and_801_ssc_1 , ActUnit_RunInst_switch_lp_and_545_ssc_1
      , ActUnit_RunInst_switch_lp_and_547_ssc_1 , ActUnit_RunInst_switch_lp_and_551_ssc_1
      , ActUnit_RunInst_switch_lp_and_553_ssc_1});
  assign while_and_265_nl = while_while_mux1h_306_nl & (~ ActUnit_RunInst_switch_lp_and_549_ssc_1);
  assign while_while_mux1h_309_nl = MUX1HOT_s_1_6_2(act_regs_data_3_5_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[191]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_6_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_6_lpi_1_dfm_1_ftd, Silu_for_y_6_lpi_1_dfm_4_31, Gelu_for_y_6_lpi_1_dfm_4_31_1,
      {while_nand_112_ssc_1 , ActUnit_RunInst_switch_lp_and_801_ssc_1 , ActUnit_RunInst_switch_lp_and_545_ssc_1
      , ActUnit_RunInst_switch_lp_and_547_ssc_1 , ActUnit_RunInst_switch_lp_and_551_ssc_1
      , ActUnit_RunInst_switch_lp_and_553_ssc_1});
  assign while_and_266_nl = while_while_mux1h_309_nl & (~ ActUnit_RunInst_switch_lp_and_549_ssc_1);
  assign while_while_mux1h_312_nl = MUX1HOT_s_1_6_2(act_regs_data_3_6_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[223]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_7_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_7_lpi_1_dfm_1_ftd, Silu_for_y_7_lpi_1_dfm_4_31, Gelu_for_y_7_lpi_1_dfm_4_31_1,
      {while_nand_112_ssc_1 , ActUnit_RunInst_switch_lp_and_801_ssc_1 , ActUnit_RunInst_switch_lp_and_545_ssc_1
      , ActUnit_RunInst_switch_lp_and_547_ssc_1 , ActUnit_RunInst_switch_lp_and_551_ssc_1
      , ActUnit_RunInst_switch_lp_and_553_ssc_1});
  assign while_and_267_nl = while_while_mux1h_312_nl & (~ ActUnit_RunInst_switch_lp_and_549_ssc_1);
  assign while_while_mux1h_315_nl = MUX1HOT_s_1_6_2(act_regs_data_3_7_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[255]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_8_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_8_lpi_1_dfm_1_ftd, Silu_for_y_8_lpi_1_dfm_4_31, Gelu_for_y_8_lpi_1_dfm_4_31_1,
      {while_nand_112_ssc_1 , ActUnit_RunInst_switch_lp_and_801_ssc_1 , ActUnit_RunInst_switch_lp_and_545_ssc_1
      , ActUnit_RunInst_switch_lp_and_547_ssc_1 , ActUnit_RunInst_switch_lp_and_551_ssc_1
      , ActUnit_RunInst_switch_lp_and_553_ssc_1});
  assign while_and_268_nl = while_while_mux1h_315_nl & (~ ActUnit_RunInst_switch_lp_and_549_ssc_1);
  assign while_while_mux1h_318_nl = MUX1HOT_s_1_6_2(act_regs_data_3_8_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[287]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_9_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_9_lpi_1_dfm_1_ftd, Silu_for_y_9_lpi_1_dfm_4_31_1, Gelu_for_y_9_lpi_1_dfm_4_31_1,
      {while_nand_112_ssc_1 , ActUnit_RunInst_switch_lp_and_801_ssc_1 , ActUnit_RunInst_switch_lp_and_545_ssc_1
      , ActUnit_RunInst_switch_lp_and_547_ssc_1 , ActUnit_RunInst_switch_lp_and_551_ssc_1
      , ActUnit_RunInst_switch_lp_and_553_ssc_1});
  assign while_and_269_nl = while_while_mux1h_318_nl & (~ ActUnit_RunInst_switch_lp_and_549_ssc_1);
  assign while_while_mux1h_321_nl = MUX1HOT_s_1_6_2(act_regs_data_3_9_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[319]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_10_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_10_lpi_1_dfm_1_ftd, Silu_for_y_10_lpi_1_dfm_4_31_1, Gelu_for_y_10_lpi_1_dfm_4_31_1,
      {while_nand_112_ssc_1 , ActUnit_RunInst_switch_lp_and_801_ssc_1 , ActUnit_RunInst_switch_lp_and_545_ssc_1
      , ActUnit_RunInst_switch_lp_and_547_ssc_1 , ActUnit_RunInst_switch_lp_and_551_ssc_1
      , ActUnit_RunInst_switch_lp_and_553_ssc_1});
  assign while_and_270_nl = while_while_mux1h_321_nl & (~ ActUnit_RunInst_switch_lp_and_549_ssc_1);
  assign while_while_mux1h_324_nl = MUX1HOT_s_1_6_2(act_regs_data_3_10_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[351]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_11_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_11_lpi_1_dfm_1_ftd, Silu_for_y_11_lpi_1_dfm_4_31_1, Gelu_for_y_11_lpi_1_dfm_4_31_1,
      {while_nand_112_ssc_1 , ActUnit_RunInst_switch_lp_and_801_ssc_1 , ActUnit_RunInst_switch_lp_and_545_ssc_1
      , ActUnit_RunInst_switch_lp_and_547_ssc_1 , ActUnit_RunInst_switch_lp_and_551_ssc_1
      , ActUnit_RunInst_switch_lp_and_553_ssc_1});
  assign while_and_271_nl = while_while_mux1h_324_nl & (~ ActUnit_RunInst_switch_lp_and_549_ssc_1);
  assign while_while_mux1h_327_nl = MUX1HOT_s_1_6_2(act_regs_data_3_11_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[383]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_12_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_12_lpi_1_dfm_1_ftd, Silu_for_y_12_lpi_1_dfm_4_31_1, Gelu_for_y_12_lpi_1_dfm_4_31_1,
      {while_nand_112_ssc_1 , ActUnit_RunInst_switch_lp_and_801_ssc_1 , ActUnit_RunInst_switch_lp_and_545_ssc_1
      , ActUnit_RunInst_switch_lp_and_547_ssc_1 , ActUnit_RunInst_switch_lp_and_551_ssc_1
      , ActUnit_RunInst_switch_lp_and_553_ssc_1});
  assign while_and_272_nl = while_while_mux1h_327_nl & (~ ActUnit_RunInst_switch_lp_and_549_ssc_1);
  assign while_while_mux1h_330_nl = MUX1HOT_s_1_6_2(act_regs_data_3_12_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[415]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_13_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_13_lpi_1_dfm_1_ftd, Silu_for_y_13_lpi_1_dfm_4_31_1, Gelu_for_y_13_lpi_1_dfm_4_31_1,
      {while_nand_112_ssc_1 , ActUnit_RunInst_switch_lp_and_801_ssc_1 , ActUnit_RunInst_switch_lp_and_545_ssc_1
      , ActUnit_RunInst_switch_lp_and_547_ssc_1 , ActUnit_RunInst_switch_lp_and_551_ssc_1
      , ActUnit_RunInst_switch_lp_and_553_ssc_1});
  assign while_and_273_nl = while_while_mux1h_330_nl & (~ ActUnit_RunInst_switch_lp_and_549_ssc_1);
  assign while_while_mux1h_333_nl = MUX1HOT_s_1_6_2(act_regs_data_3_13_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[447]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_14_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_14_lpi_1_dfm_1_ftd, Silu_for_y_14_lpi_1_dfm_4_31_1, Gelu_for_y_14_lpi_1_dfm_4_31_1,
      {while_nand_112_ssc_1 , ActUnit_RunInst_switch_lp_and_801_ssc_1 , ActUnit_RunInst_switch_lp_and_545_ssc_1
      , ActUnit_RunInst_switch_lp_and_547_ssc_1 , ActUnit_RunInst_switch_lp_and_551_ssc_1
      , ActUnit_RunInst_switch_lp_and_553_ssc_1});
  assign while_and_274_nl = while_while_mux1h_333_nl & (~ ActUnit_RunInst_switch_lp_and_549_ssc_1);
  assign while_while_mux1h_336_nl = MUX1HOT_s_1_6_2(act_regs_data_3_14_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[479]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_15_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_15_lpi_1_dfm_1_ftd, Silu_for_y_15_lpi_1_dfm_4_31_1, Gelu_for_y_15_lpi_1_dfm_4_31_1,
      {while_nand_112_ssc_1 , ActUnit_RunInst_switch_lp_and_801_ssc_1 , ActUnit_RunInst_switch_lp_and_545_ssc_1
      , ActUnit_RunInst_switch_lp_and_547_ssc_1 , ActUnit_RunInst_switch_lp_and_551_ssc_1
      , ActUnit_RunInst_switch_lp_and_553_ssc_1});
  assign while_and_275_nl = while_while_mux1h_336_nl & (~ ActUnit_RunInst_switch_lp_and_549_ssc_1);
  assign while_while_mux1h_339_nl = MUX1HOT_s_1_6_2(act_regs_data_3_15_sva_31, (ActUnit_RunInst_case_3_act_port_reg_data_sva[511]),
      nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_16_nvhls_nv_scvector_spec_ActScalarType_16U_operator_4_for_slc_act_regs_data_32_31_0_1_ctmp_sva_31,
      reg_Tanh_for_y_25_0_lpi_1_dfm_1_ftd, Silu_for_y_lpi_1_dfm_4_31_1, Gelu_for_y_lpi_1_dfm_4_31_1,
      {while_nand_112_ssc_1 , ActUnit_RunInst_switch_lp_and_801_ssc_1 , ActUnit_RunInst_switch_lp_and_545_ssc_1
      , ActUnit_RunInst_switch_lp_and_547_ssc_1 , ActUnit_RunInst_switch_lp_and_551_ssc_1
      , ActUnit_RunInst_switch_lp_and_553_ssc_1});
  assign while_and_276_nl = while_while_mux1h_339_nl & (~ ActUnit_RunInst_switch_lp_and_549_ssc_1);
  assign act_config_InstIncr_if_act_config_InstIncr_if_and_nl = act_config_is_zero_first_sva_dfm_4
      & (~ act_config_InstIncr_if_act_config_InstIncr_if_if_nor_tmp);
  assign act_config_InstIncr_mux_2_nl = MUX_s_1_2_2(act_config_is_zero_first_sva_dfm_4,
      act_config_InstIncr_if_act_config_InstIncr_if_and_nl, act_config_InstIncr_act_config_InstIncr_if_and_svs_1);
  assign nor_1650_nl = ~((~ (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[0])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[8])
      | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[10]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[9])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0])));
  assign or_3343_nl = (rva_in_PopNB_mioi_data_data_rsc_z_mxwt[0]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[8])
      | (~ rva_in_PopNB_mioi_data_rw_rsc_z_mxwt) | (~ rva_in_PopNB_mioi_return_rsc_z_mxwt)
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[10]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[9])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[11])) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[7])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[6]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[5])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[3]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[2])
      | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[4]) | (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[1])
      | (~ (rva_in_PopNB_mioi_data_addr_rsc_z_mxwt[0]));
  assign mux_1474_nl = MUX_s_1_2_2(nor_1650_nl, or_3343_nl, act_config_is_valid_sva);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_122_nl = MUX_v_22_2_2(22'b0000000000000000000000,
      act_regs_data_0_0_sva_dfm_2_21_0, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_291);
  assign mux1h_11_nl = MUX1HOT_v_22_3_2((Silu_for_1_else_if_Silu_for_else_if_mul_cmp_6_z[44:23]),
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_21_0_mx0w1,
      act_regs_data_0_1_sva_dfm_2_21_0, {and_dcpl_1112 , and_dcpl_1393 , and_1720_cse});
  assign not_2658_nl = ~ or_dcpl_1012;
  assign and_1777_nl = MUX_v_22_2_2(22'b0000000000000000000000, mux1h_11_nl, not_2658_nl);
  assign and_1442_nl = and_dcpl_1235 & and_dcpl_1396 & and_dcpl_1395;
  assign mux1h_12_nl = MUX1HOT_v_22_3_2((Silu_for_1_else_if_Silu_for_else_if_mul_cmp_5_z[44:23]),
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_21_0_mx0w1,
      act_regs_data_0_10_sva_dfm_2_21_0, {and_dcpl_1112 , and_1442_nl , and_1720_cse});
  assign not_2660_nl = ~ or_dcpl_1012;
  assign and_1782_nl = MUX_v_22_2_2(22'b0000000000000000000000, mux1h_12_nl, not_2660_nl);
  assign and_1445_nl = and_dcpl_1235 & and_dcpl_1396 & and_2344_cse;
  assign mux1h_13_nl = MUX1HOT_v_22_3_2((Silu_for_1_else_if_Silu_for_else_if_mul_cmp_4_z[44:23]),
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_21_0_mx0w1,
      act_regs_data_0_11_sva_dfm_2_21_0, {and_dcpl_1112 , and_1445_nl , and_1720_cse});
  assign not_2662_nl = ~ or_dcpl_1012;
  assign and_1786_nl = MUX_v_22_2_2(22'b0000000000000000000000, mux1h_13_nl, not_2662_nl);
  assign and_1448_nl = and_dcpl_1235 & and_dcpl_1402 & nor_1553_cse;
  assign mux1h_14_nl = MUX1HOT_v_22_3_2((Silu_for_1_else_if_Silu_for_else_if_mul_cmp_3_z[44:23]),
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_21_0_mx0w1,
      act_regs_data_0_12_sva_dfm_2_21_0, {and_dcpl_1112 , and_1448_nl , and_1720_cse});
  assign not_2664_nl = ~ or_dcpl_1012;
  assign and_1790_nl = MUX_v_22_2_2(22'b0000000000000000000000, mux1h_14_nl, not_2664_nl);
  assign and_1450_nl = and_dcpl_1235 & and_dcpl_1402 & and_dcpl_1391;
  assign mux1h_15_nl = MUX1HOT_v_22_3_2((Silu_for_1_else_if_Silu_for_else_if_mul_cmp_2_z[44:23]),
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_21_0_mx0w1,
      act_regs_data_0_13_sva_dfm_2_21_0, {and_dcpl_1112 , and_1450_nl , and_1720_cse});
  assign not_2666_nl = ~ or_dcpl_1012;
  assign and_1794_nl = MUX_v_22_2_2(22'b0000000000000000000000, mux1h_15_nl, not_2666_nl);
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_6_nl = act_regs_data_0_0_sva_dfm_2_25_22_rsp_0
      & nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_291;
  assign nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_and_304_nl = MUX_v_3_2_2(3'b000,
      act_regs_data_0_0_sva_dfm_2_25_22_rsp_1, nvhls_nv_scvector_spec_ActScalarType_16U_operator_13_for_not_291);
  assign mux1h_nl = MUX1HOT_s_1_3_2((Silu_for_13_else_else_else_else_if_acc_sdt[3]),
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_25_22_mx0w2_3,
      act_regs_data_0_1_sva_dfm_2_25_22_rsp_0, {and_dcpl_331 , and_dcpl_1393 , and_1715_ssc});
  assign and_1711_nl = mux1h_nl & (~ or_1527_tmp);
  assign mux1h_16_nl = MUX1HOT_v_3_3_2((Silu_for_13_else_else_else_else_if_acc_sdt[2:0]),
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_25_22_mx0w2_2_0,
      act_regs_data_0_1_sva_dfm_2_25_22_rsp_1, {and_dcpl_331 , and_dcpl_1393 , and_1715_ssc});
  assign not_8904_nl = ~ or_1527_tmp;
  assign and_3505_nl = MUX_v_3_2_2(3'b000, mux1h_16_nl, not_8904_nl);
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_9_nl = MUX1HOT_s_1_3_2((Silu_for_14_else_else_else_else_if_acc_sdt[3]),
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_25_22_mx0w2_3,
      act_regs_data_0_10_sva_dfm_2_25_22_rsp_0, {and_dcpl_331 , and_dcpl_1235 , and_dcpl_1236});
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_191_nl = MUX1HOT_v_3_3_2((Silu_for_14_else_else_else_else_if_acc_sdt[2:0]),
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_25_22_mx0w2_2_0,
      act_regs_data_0_10_sva_dfm_2_25_22_rsp_1, {and_dcpl_331 , and_dcpl_1235 , and_dcpl_1236});
  assign not_8895_nl = ~ or_dcpl;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_14_nl = MUX1HOT_s_1_3_2((Silu_for_15_else_else_else_else_if_acc_sdt[3]),
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_25_22_mx0w2_3,
      act_regs_data_0_11_sva_dfm_2_25_22_rsp_0, {and_dcpl_331 , and_dcpl_1235 , and_dcpl_1236});
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_190_nl = MUX1HOT_v_3_3_2((Silu_for_15_else_else_else_else_if_acc_sdt[2:0]),
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_25_22_mx0w2_2_0,
      act_regs_data_0_11_sva_dfm_2_25_22_rsp_1, {and_dcpl_331 , and_dcpl_1235 , and_dcpl_1236});
  assign not_8894_nl = ~ or_dcpl;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_19_nl = MUX1HOT_s_1_3_2((Silu_for_16_else_else_else_else_if_acc_sdt[3]),
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_25_22_mx0w2_3,
      act_regs_data_0_12_sva_dfm_2_25_22_rsp_0, {and_dcpl_331 , and_dcpl_1235 , and_dcpl_1236});
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_189_nl = MUX1HOT_v_3_3_2((Silu_for_16_else_else_else_else_if_acc_sdt[2:0]),
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_25_22_mx0w2_2_0,
      act_regs_data_0_12_sva_dfm_2_25_22_rsp_1, {and_dcpl_331 , and_dcpl_1235 , and_dcpl_1236});
  assign not_8893_nl = ~ or_dcpl;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_24_nl = MUX1HOT_s_1_3_2((Silu_for_1_else_else_else_else_if_acc_sdt[3]),
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_25_22_mx0w2_3,
      act_regs_data_0_13_sva_dfm_2_25_22_rsp_0, {and_dcpl_331 , and_dcpl_1235 , and_dcpl_1236});
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_188_nl = MUX1HOT_v_3_3_2((Silu_for_1_else_else_else_else_if_acc_sdt[2:0]),
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_25_22_mx0w2_2_0,
      act_regs_data_0_13_sva_dfm_2_25_22_rsp_1, {and_dcpl_331 , and_dcpl_1235 , and_dcpl_1236});
  assign not_8892_nl = ~ or_dcpl;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_29_nl = MUX1HOT_s_1_3_2((Silu_for_2_else_else_else_else_if_acc_sdt[3]),
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_25_22_mx0w2_3,
      act_regs_data_0_14_sva_dfm_2_25_22_rsp_0, {and_dcpl_331 , and_dcpl_1235 , and_dcpl_1236});
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_187_nl = MUX1HOT_v_3_3_2((Silu_for_2_else_else_else_else_if_acc_sdt[2:0]),
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_25_22_mx0w2_2_0,
      act_regs_data_0_14_sva_dfm_2_25_22_rsp_1, {and_dcpl_331 , and_dcpl_1235 , and_dcpl_1236});
  assign not_8891_nl = ~ or_dcpl;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_34_nl = MUX1HOT_s_1_3_2((Silu_for_3_else_else_else_else_if_acc_sdt[3]),
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_25_22_mx0w2_3,
      act_regs_data_0_15_sva_dfm_2_25_22_rsp_0, {and_dcpl_331 , and_dcpl_1235 , and_dcpl_1236});
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_198_nl = MUX1HOT_v_3_3_2((Silu_for_3_else_else_else_else_if_acc_sdt[2:0]),
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_25_22_mx0w2_2_0,
      act_regs_data_0_15_sva_dfm_2_25_22_rsp_1, {and_dcpl_331 , and_dcpl_1235 , and_dcpl_1236});
  assign not_8903_nl = ~ or_dcpl;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_39_nl = MUX1HOT_s_1_3_2((Silu_for_4_else_else_else_else_if_acc_sdt[3]),
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_25_22_mx0w2_3,
      act_regs_data_0_2_sva_dfm_2_25_22_rsp_0, {and_dcpl_331 , and_dcpl_1235 , and_dcpl_1236});
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_197_nl = MUX1HOT_v_3_3_2((Silu_for_4_else_else_else_else_if_acc_sdt[2:0]),
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_25_22_mx0w2_2_0,
      act_regs_data_0_2_sva_dfm_2_25_22_rsp_1, {and_dcpl_331 , and_dcpl_1235 , and_dcpl_1236});
  assign not_8902_nl = ~ or_dcpl;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_44_nl = MUX1HOT_s_1_3_2((Silu_for_5_else_else_else_else_if_acc_sdt[3]),
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_25_22_mx0w2_3,
      act_regs_data_0_3_sva_dfm_2_25_22_rsp_0, {and_dcpl_331 , and_dcpl_1235 , and_dcpl_1236});
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_196_nl = MUX1HOT_v_3_3_2((Silu_for_5_else_else_else_else_if_acc_sdt[2:0]),
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_25_22_mx0w2_2_0,
      act_regs_data_0_3_sva_dfm_2_25_22_rsp_1, {and_dcpl_331 , and_dcpl_1235 , and_dcpl_1236});
  assign not_8901_nl = ~ or_dcpl;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_49_nl = MUX1HOT_s_1_3_2((Silu_for_6_else_else_else_else_if_acc_sdt[3]),
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_25_22_mx0w2_3,
      act_regs_data_0_4_sva_dfm_2_25_22_rsp_0, {and_dcpl_331 , and_dcpl_1235 , and_dcpl_1236});
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_195_nl = MUX1HOT_v_3_3_2((Silu_for_6_else_else_else_else_if_acc_sdt[2:0]),
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_25_22_mx0w2_2_0,
      act_regs_data_0_4_sva_dfm_2_25_22_rsp_1, {and_dcpl_331 , and_dcpl_1235 , and_dcpl_1236});
  assign not_8900_nl = ~ or_dcpl;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_54_nl = MUX1HOT_s_1_3_2((Silu_for_7_else_else_else_else_if_acc_sdt[3]),
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_25_22_mx0w2_3,
      act_regs_data_0_5_sva_dfm_2_25_22_rsp_0, {and_dcpl_331 , and_dcpl_1235 , and_dcpl_1236});
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_194_nl = MUX1HOT_v_3_3_2((Silu_for_7_else_else_else_else_if_acc_sdt[2:0]),
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_25_22_mx0w2_2_0,
      act_regs_data_0_5_sva_dfm_2_25_22_rsp_1, {and_dcpl_331 , and_dcpl_1235 , and_dcpl_1236});
  assign not_8899_nl = ~ or_dcpl;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_59_nl = MUX1HOT_s_1_3_2((Silu_for_8_else_else_else_else_if_acc_sdt[3]),
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_25_22_mx0w2_3,
      act_regs_data_0_6_sva_dfm_2_25_22_rsp_0, {and_dcpl_331 , and_dcpl_1235 , and_dcpl_1236});
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_193_nl = MUX1HOT_v_3_3_2((Silu_for_8_else_else_else_else_if_acc_sdt[2:0]),
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_25_22_mx0w2_2_0,
      act_regs_data_0_6_sva_dfm_2_25_22_rsp_1, {and_dcpl_331 , and_dcpl_1235 , and_dcpl_1236});
  assign not_8898_nl = ~ or_dcpl;
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_64_nl = MUX1HOT_s_1_3_2((Silu_for_9_else_else_else_else_if_acc_sdt[3]),
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_25_22_mx0w2_3,
      act_regs_data_0_7_sva_dfm_2_25_22_rsp_0, {and_dcpl_331 , and_dcpl_1235 , and_dcpl_1236});
  assign ActUnit_PushOutput_if_output_port_reg_data_data_mux1h_192_nl = MUX1HOT_v_3_3_2((Silu_for_9_else_else_else_else_if_acc_sdt[2:0]),
      ActUnit_PushOutput_if_for_slc_act_regs_data_32_31_0_2_ctmp_sva_25_22_mx0w2_2_0,
      act_regs_data_0_7_sva_dfm_2_25_22_rsp_1, {and_dcpl_331 , and_dcpl_1235 , and_dcpl_1236});
  assign not_8897_nl = ~ or_dcpl;
  assign Silu_for_else_else_else_else_if_mux_nl = MUX_v_4_2_2(({reg_nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_0
      , reg_nv_scvector_cctor_nv_scvector_5_for_10_nv_scvector_cctor_nv_scvector_5_for_slc_act_regs_data_32_31_0_1_ncse_1_ftd_rsp_1}),
      ActUnit_PushOutput_if_for_i_4_0_sva_3_0, not_tmp_646);
  assign nl_z_out = conv_u2u_4_5(Silu_for_else_else_else_else_if_mux_nl) + conv_s2u_2_5({(~
      not_tmp_646) , 1'b1});
  assign z_out = nl_z_out[4:0];

  function automatic  MUX1HOT_s_1_1_2;
    input  input_0;
    input  sel;
    reg  result;
  begin
    result = input_0 & sel;
    MUX1HOT_s_1_1_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_3_2;
    input  input_2;
    input  input_1;
    input  input_0;
    input [2:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_4_2;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [3:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_5_2;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [4:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    MUX1HOT_s_1_5_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_6_2;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [5:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    MUX1HOT_s_1_6_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_8_2;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [7:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    MUX1HOT_s_1_8_2 = result;
  end
  endfunction


  function automatic [19:0] MUX1HOT_v_20_4_2;
    input [19:0] input_3;
    input [19:0] input_2;
    input [19:0] input_1;
    input [19:0] input_0;
    input [3:0] sel;
    reg [19:0] result;
  begin
    result = input_0 & {20{sel[0]}};
    result = result | (input_1 & {20{sel[1]}});
    result = result | (input_2 & {20{sel[2]}});
    result = result | (input_3 & {20{sel[3]}});
    MUX1HOT_v_20_4_2 = result;
  end
  endfunction


  function automatic [21:0] MUX1HOT_v_22_3_2;
    input [21:0] input_2;
    input [21:0] input_1;
    input [21:0] input_0;
    input [2:0] sel;
    reg [21:0] result;
  begin
    result = input_0 & {22{sel[0]}};
    result = result | (input_1 & {22{sel[1]}});
    result = result | (input_2 & {22{sel[2]}});
    MUX1HOT_v_22_3_2 = result;
  end
  endfunction


  function automatic [21:0] MUX1HOT_v_22_4_2;
    input [21:0] input_3;
    input [21:0] input_2;
    input [21:0] input_1;
    input [21:0] input_0;
    input [3:0] sel;
    reg [21:0] result;
  begin
    result = input_0 & {22{sel[0]}};
    result = result | (input_1 & {22{sel[1]}});
    result = result | (input_2 & {22{sel[2]}});
    result = result | (input_3 & {22{sel[3]}});
    MUX1HOT_v_22_4_2 = result;
  end
  endfunction


  function automatic [21:0] MUX1HOT_v_22_8_2;
    input [21:0] input_7;
    input [21:0] input_6;
    input [21:0] input_5;
    input [21:0] input_4;
    input [21:0] input_3;
    input [21:0] input_2;
    input [21:0] input_1;
    input [21:0] input_0;
    input [7:0] sel;
    reg [21:0] result;
  begin
    result = input_0 & {22{sel[0]}};
    result = result | (input_1 & {22{sel[1]}});
    result = result | (input_2 & {22{sel[2]}});
    result = result | (input_3 & {22{sel[3]}});
    result = result | (input_4 & {22{sel[4]}});
    result = result | (input_5 & {22{sel[5]}});
    result = result | (input_6 & {22{sel[6]}});
    result = result | (input_7 & {22{sel[7]}});
    MUX1HOT_v_22_8_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_4_2;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [3:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    result = result | (input_3 & {2{sel[3]}});
    MUX1HOT_v_2_4_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_3_2;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [2:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | (input_1 & {3{sel[1]}});
    result = result | (input_2 & {3{sel[2]}});
    MUX1HOT_v_3_3_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_4_2;
    input [2:0] input_3;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [3:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | (input_1 & {3{sel[1]}});
    result = result | (input_2 & {3{sel[2]}});
    result = result | (input_3 & {3{sel[3]}});
    MUX1HOT_v_3_4_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_5_2;
    input [2:0] input_4;
    input [2:0] input_3;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [4:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | (input_1 & {3{sel[1]}});
    result = result | (input_2 & {3{sel[2]}});
    result = result | (input_3 & {3{sel[3]}});
    result = result | (input_4 & {3{sel[4]}});
    MUX1HOT_v_3_5_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_8_2;
    input [2:0] input_7;
    input [2:0] input_6;
    input [2:0] input_5;
    input [2:0] input_4;
    input [2:0] input_3;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [7:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | (input_1 & {3{sel[1]}});
    result = result | (input_2 & {3{sel[2]}});
    result = result | (input_3 & {3{sel[3]}});
    result = result | (input_4 & {3{sel[4]}});
    result = result | (input_5 & {3{sel[5]}});
    result = result | (input_6 & {3{sel[6]}});
    result = result | (input_7 & {3{sel[7]}});
    MUX1HOT_v_3_8_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_4_2;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [3:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    MUX1HOT_v_4_4_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_3_2;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [2:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    MUX1HOT_v_5_3_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_4_2;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [3:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    result = result | (input_3 & {5{sel[3]}});
    MUX1HOT_v_5_4_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_5_2;
    input [4:0] input_4;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [4:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    result = result | (input_3 & {5{sel[3]}});
    result = result | (input_4 & {5{sel[4]}});
    MUX1HOT_v_5_5_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_8_2;
    input [4:0] input_7;
    input [4:0] input_6;
    input [4:0] input_5;
    input [4:0] input_4;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [7:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    result = result | (input_3 & {5{sel[3]}});
    result = result | (input_4 & {5{sel[4]}});
    result = result | (input_5 & {5{sel[5]}});
    result = result | (input_6 & {5{sel[6]}});
    result = result | (input_7 & {5{sel[7]}});
    MUX1HOT_v_5_8_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_4_2;
    input  input_0;
    input  input_1;
    input  input_2;
    input  input_3;
    input [1:0] sel;
    reg  result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      2'b10 : begin
        result = input_2;
      end
      default : begin
        result = input_3;
      end
    endcase
    MUX_s_1_4_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_64_2;
    input  input_0;
    input  input_1;
    input  input_2;
    input  input_3;
    input  input_4;
    input  input_5;
    input  input_6;
    input  input_7;
    input  input_8;
    input  input_9;
    input  input_10;
    input  input_11;
    input  input_12;
    input  input_13;
    input  input_14;
    input  input_15;
    input  input_16;
    input  input_17;
    input  input_18;
    input  input_19;
    input  input_20;
    input  input_21;
    input  input_22;
    input  input_23;
    input  input_24;
    input  input_25;
    input  input_26;
    input  input_27;
    input  input_28;
    input  input_29;
    input  input_30;
    input  input_31;
    input  input_32;
    input  input_33;
    input  input_34;
    input  input_35;
    input  input_36;
    input  input_37;
    input  input_38;
    input  input_39;
    input  input_40;
    input  input_41;
    input  input_42;
    input  input_43;
    input  input_44;
    input  input_45;
    input  input_46;
    input  input_47;
    input  input_48;
    input  input_49;
    input  input_50;
    input  input_51;
    input  input_52;
    input  input_53;
    input  input_54;
    input  input_55;
    input  input_56;
    input  input_57;
    input  input_58;
    input  input_59;
    input  input_60;
    input  input_61;
    input  input_62;
    input  input_63;
    input [5:0] sel;
    reg  result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      6'b110111 : begin
        result = input_55;
      end
      6'b111000 : begin
        result = input_56;
      end
      6'b111001 : begin
        result = input_57;
      end
      6'b111010 : begin
        result = input_58;
      end
      6'b111011 : begin
        result = input_59;
      end
      6'b111100 : begin
        result = input_60;
      end
      6'b111101 : begin
        result = input_61;
      end
      6'b111110 : begin
        result = input_62;
      end
      default : begin
        result = input_63;
      end
    endcase
    MUX_s_1_64_2 = result;
  end
  endfunction


  function automatic [21:0] MUX_v_22_2_2;
    input [21:0] input_0;
    input [21:0] input_1;
    input  sel;
    reg [21:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_22_2_2 = result;
  end
  endfunction


  function automatic [21:0] MUX_v_22_4_2;
    input [21:0] input_0;
    input [21:0] input_1;
    input [21:0] input_2;
    input [21:0] input_3;
    input [1:0] sel;
    reg [21:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      2'b10 : begin
        result = input_2;
      end
      default : begin
        result = input_3;
      end
    endcase
    MUX_v_22_4_2 = result;
  end
  endfunction


  function automatic [21:0] MUX_v_22_64_2;
    input [21:0] input_0;
    input [21:0] input_1;
    input [21:0] input_2;
    input [21:0] input_3;
    input [21:0] input_4;
    input [21:0] input_5;
    input [21:0] input_6;
    input [21:0] input_7;
    input [21:0] input_8;
    input [21:0] input_9;
    input [21:0] input_10;
    input [21:0] input_11;
    input [21:0] input_12;
    input [21:0] input_13;
    input [21:0] input_14;
    input [21:0] input_15;
    input [21:0] input_16;
    input [21:0] input_17;
    input [21:0] input_18;
    input [21:0] input_19;
    input [21:0] input_20;
    input [21:0] input_21;
    input [21:0] input_22;
    input [21:0] input_23;
    input [21:0] input_24;
    input [21:0] input_25;
    input [21:0] input_26;
    input [21:0] input_27;
    input [21:0] input_28;
    input [21:0] input_29;
    input [21:0] input_30;
    input [21:0] input_31;
    input [21:0] input_32;
    input [21:0] input_33;
    input [21:0] input_34;
    input [21:0] input_35;
    input [21:0] input_36;
    input [21:0] input_37;
    input [21:0] input_38;
    input [21:0] input_39;
    input [21:0] input_40;
    input [21:0] input_41;
    input [21:0] input_42;
    input [21:0] input_43;
    input [21:0] input_44;
    input [21:0] input_45;
    input [21:0] input_46;
    input [21:0] input_47;
    input [21:0] input_48;
    input [21:0] input_49;
    input [21:0] input_50;
    input [21:0] input_51;
    input [21:0] input_52;
    input [21:0] input_53;
    input [21:0] input_54;
    input [21:0] input_55;
    input [21:0] input_56;
    input [21:0] input_57;
    input [21:0] input_58;
    input [21:0] input_59;
    input [21:0] input_60;
    input [21:0] input_61;
    input [21:0] input_62;
    input [21:0] input_63;
    input [5:0] sel;
    reg [21:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      6'b110111 : begin
        result = input_55;
      end
      6'b111000 : begin
        result = input_56;
      end
      6'b111001 : begin
        result = input_57;
      end
      6'b111010 : begin
        result = input_58;
      end
      6'b111011 : begin
        result = input_59;
      end
      6'b111100 : begin
        result = input_60;
      end
      6'b111101 : begin
        result = input_61;
      end
      6'b111110 : begin
        result = input_62;
      end
      default : begin
        result = input_63;
      end
    endcase
    MUX_v_22_64_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input  sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_32_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [1:0] input_2;
    input [1:0] input_3;
    input [1:0] input_4;
    input [1:0] input_5;
    input [1:0] input_6;
    input [1:0] input_7;
    input [1:0] input_8;
    input [1:0] input_9;
    input [1:0] input_10;
    input [1:0] input_11;
    input [1:0] input_12;
    input [1:0] input_13;
    input [1:0] input_14;
    input [1:0] input_15;
    input [1:0] input_16;
    input [1:0] input_17;
    input [1:0] input_18;
    input [1:0] input_19;
    input [1:0] input_20;
    input [1:0] input_21;
    input [1:0] input_22;
    input [1:0] input_23;
    input [1:0] input_24;
    input [1:0] input_25;
    input [1:0] input_26;
    input [1:0] input_27;
    input [1:0] input_28;
    input [1:0] input_29;
    input [1:0] input_30;
    input [1:0] input_31;
    input [4:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      5'b00000 : begin
        result = input_0;
      end
      5'b00001 : begin
        result = input_1;
      end
      5'b00010 : begin
        result = input_2;
      end
      5'b00011 : begin
        result = input_3;
      end
      5'b00100 : begin
        result = input_4;
      end
      5'b00101 : begin
        result = input_5;
      end
      5'b00110 : begin
        result = input_6;
      end
      5'b00111 : begin
        result = input_7;
      end
      5'b01000 : begin
        result = input_8;
      end
      5'b01001 : begin
        result = input_9;
      end
      5'b01010 : begin
        result = input_10;
      end
      5'b01011 : begin
        result = input_11;
      end
      5'b01100 : begin
        result = input_12;
      end
      5'b01101 : begin
        result = input_13;
      end
      5'b01110 : begin
        result = input_14;
      end
      5'b01111 : begin
        result = input_15;
      end
      5'b10000 : begin
        result = input_16;
      end
      5'b10001 : begin
        result = input_17;
      end
      5'b10010 : begin
        result = input_18;
      end
      5'b10011 : begin
        result = input_19;
      end
      5'b10100 : begin
        result = input_20;
      end
      5'b10101 : begin
        result = input_21;
      end
      5'b10110 : begin
        result = input_22;
      end
      5'b10111 : begin
        result = input_23;
      end
      5'b11000 : begin
        result = input_24;
      end
      5'b11001 : begin
        result = input_25;
      end
      5'b11010 : begin
        result = input_26;
      end
      5'b11011 : begin
        result = input_27;
      end
      5'b11100 : begin
        result = input_28;
      end
      5'b11101 : begin
        result = input_29;
      end
      5'b11110 : begin
        result = input_30;
      end
      default : begin
        result = input_31;
      end
    endcase
    MUX_v_2_32_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_16_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [31:0] input_3;
    input [31:0] input_4;
    input [31:0] input_5;
    input [31:0] input_6;
    input [31:0] input_7;
    input [31:0] input_8;
    input [31:0] input_9;
    input [31:0] input_10;
    input [31:0] input_11;
    input [31:0] input_12;
    input [31:0] input_13;
    input [31:0] input_14;
    input [31:0] input_15;
    input [3:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      4'b0000 : begin
        result = input_0;
      end
      4'b0001 : begin
        result = input_1;
      end
      4'b0010 : begin
        result = input_2;
      end
      4'b0011 : begin
        result = input_3;
      end
      4'b0100 : begin
        result = input_4;
      end
      4'b0101 : begin
        result = input_5;
      end
      4'b0110 : begin
        result = input_6;
      end
      4'b0111 : begin
        result = input_7;
      end
      4'b1000 : begin
        result = input_8;
      end
      4'b1001 : begin
        result = input_9;
      end
      4'b1010 : begin
        result = input_10;
      end
      4'b1011 : begin
        result = input_11;
      end
      4'b1100 : begin
        result = input_12;
      end
      4'b1101 : begin
        result = input_13;
      end
      4'b1110 : begin
        result = input_14;
      end
      default : begin
        result = input_15;
      end
    endcase
    MUX_v_32_16_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input  sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_32_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [31:0] input_3;
    input [31:0] input_4;
    input [31:0] input_5;
    input [31:0] input_6;
    input [31:0] input_7;
    input [31:0] input_8;
    input [31:0] input_9;
    input [31:0] input_10;
    input [31:0] input_11;
    input [31:0] input_12;
    input [31:0] input_13;
    input [31:0] input_14;
    input [31:0] input_15;
    input [31:0] input_16;
    input [31:0] input_17;
    input [31:0] input_18;
    input [31:0] input_19;
    input [31:0] input_20;
    input [31:0] input_21;
    input [31:0] input_22;
    input [31:0] input_23;
    input [31:0] input_24;
    input [31:0] input_25;
    input [31:0] input_26;
    input [31:0] input_27;
    input [31:0] input_28;
    input [31:0] input_29;
    input [31:0] input_30;
    input [31:0] input_31;
    input [4:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      5'b00000 : begin
        result = input_0;
      end
      5'b00001 : begin
        result = input_1;
      end
      5'b00010 : begin
        result = input_2;
      end
      5'b00011 : begin
        result = input_3;
      end
      5'b00100 : begin
        result = input_4;
      end
      5'b00101 : begin
        result = input_5;
      end
      5'b00110 : begin
        result = input_6;
      end
      5'b00111 : begin
        result = input_7;
      end
      5'b01000 : begin
        result = input_8;
      end
      5'b01001 : begin
        result = input_9;
      end
      5'b01010 : begin
        result = input_10;
      end
      5'b01011 : begin
        result = input_11;
      end
      5'b01100 : begin
        result = input_12;
      end
      5'b01101 : begin
        result = input_13;
      end
      5'b01110 : begin
        result = input_14;
      end
      5'b01111 : begin
        result = input_15;
      end
      5'b10000 : begin
        result = input_16;
      end
      5'b10001 : begin
        result = input_17;
      end
      5'b10010 : begin
        result = input_18;
      end
      5'b10011 : begin
        result = input_19;
      end
      5'b10100 : begin
        result = input_20;
      end
      5'b10101 : begin
        result = input_21;
      end
      5'b10110 : begin
        result = input_22;
      end
      5'b10111 : begin
        result = input_23;
      end
      5'b11000 : begin
        result = input_24;
      end
      5'b11001 : begin
        result = input_25;
      end
      5'b11010 : begin
        result = input_26;
      end
      5'b11011 : begin
        result = input_27;
      end
      5'b11100 : begin
        result = input_28;
      end
      5'b11101 : begin
        result = input_29;
      end
      5'b11110 : begin
        result = input_30;
      end
      default : begin
        result = input_31;
      end
    endcase
    MUX_v_32_32_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input  sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_4_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [2:0] input_2;
    input [2:0] input_3;
    input [1:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      2'b10 : begin
        result = input_2;
      end
      default : begin
        result = input_3;
      end
    endcase
    MUX_v_3_4_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_64_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [2:0] input_2;
    input [2:0] input_3;
    input [2:0] input_4;
    input [2:0] input_5;
    input [2:0] input_6;
    input [2:0] input_7;
    input [2:0] input_8;
    input [2:0] input_9;
    input [2:0] input_10;
    input [2:0] input_11;
    input [2:0] input_12;
    input [2:0] input_13;
    input [2:0] input_14;
    input [2:0] input_15;
    input [2:0] input_16;
    input [2:0] input_17;
    input [2:0] input_18;
    input [2:0] input_19;
    input [2:0] input_20;
    input [2:0] input_21;
    input [2:0] input_22;
    input [2:0] input_23;
    input [2:0] input_24;
    input [2:0] input_25;
    input [2:0] input_26;
    input [2:0] input_27;
    input [2:0] input_28;
    input [2:0] input_29;
    input [2:0] input_30;
    input [2:0] input_31;
    input [2:0] input_32;
    input [2:0] input_33;
    input [2:0] input_34;
    input [2:0] input_35;
    input [2:0] input_36;
    input [2:0] input_37;
    input [2:0] input_38;
    input [2:0] input_39;
    input [2:0] input_40;
    input [2:0] input_41;
    input [2:0] input_42;
    input [2:0] input_43;
    input [2:0] input_44;
    input [2:0] input_45;
    input [2:0] input_46;
    input [2:0] input_47;
    input [2:0] input_48;
    input [2:0] input_49;
    input [2:0] input_50;
    input [2:0] input_51;
    input [2:0] input_52;
    input [2:0] input_53;
    input [2:0] input_54;
    input [2:0] input_55;
    input [2:0] input_56;
    input [2:0] input_57;
    input [2:0] input_58;
    input [2:0] input_59;
    input [2:0] input_60;
    input [2:0] input_61;
    input [2:0] input_62;
    input [2:0] input_63;
    input [5:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      6'b110111 : begin
        result = input_55;
      end
      6'b111000 : begin
        result = input_56;
      end
      6'b111001 : begin
        result = input_57;
      end
      6'b111010 : begin
        result = input_58;
      end
      6'b111011 : begin
        result = input_59;
      end
      6'b111100 : begin
        result = input_60;
      end
      6'b111101 : begin
        result = input_61;
      end
      6'b111110 : begin
        result = input_62;
      end
      default : begin
        result = input_63;
      end
    endcase
    MUX_v_3_64_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input  sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input  sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_4_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [4:0] input_2;
    input [4:0] input_3;
    input [1:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      2'b10 : begin
        result = input_2;
      end
      default : begin
        result = input_3;
      end
    endcase
    MUX_v_5_4_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_64_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [4:0] input_2;
    input [4:0] input_3;
    input [4:0] input_4;
    input [4:0] input_5;
    input [4:0] input_6;
    input [4:0] input_7;
    input [4:0] input_8;
    input [4:0] input_9;
    input [4:0] input_10;
    input [4:0] input_11;
    input [4:0] input_12;
    input [4:0] input_13;
    input [4:0] input_14;
    input [4:0] input_15;
    input [4:0] input_16;
    input [4:0] input_17;
    input [4:0] input_18;
    input [4:0] input_19;
    input [4:0] input_20;
    input [4:0] input_21;
    input [4:0] input_22;
    input [4:0] input_23;
    input [4:0] input_24;
    input [4:0] input_25;
    input [4:0] input_26;
    input [4:0] input_27;
    input [4:0] input_28;
    input [4:0] input_29;
    input [4:0] input_30;
    input [4:0] input_31;
    input [4:0] input_32;
    input [4:0] input_33;
    input [4:0] input_34;
    input [4:0] input_35;
    input [4:0] input_36;
    input [4:0] input_37;
    input [4:0] input_38;
    input [4:0] input_39;
    input [4:0] input_40;
    input [4:0] input_41;
    input [4:0] input_42;
    input [4:0] input_43;
    input [4:0] input_44;
    input [4:0] input_45;
    input [4:0] input_46;
    input [4:0] input_47;
    input [4:0] input_48;
    input [4:0] input_49;
    input [4:0] input_50;
    input [4:0] input_51;
    input [4:0] input_52;
    input [4:0] input_53;
    input [4:0] input_54;
    input [4:0] input_55;
    input [4:0] input_56;
    input [4:0] input_57;
    input [4:0] input_58;
    input [4:0] input_59;
    input [4:0] input_60;
    input [4:0] input_61;
    input [4:0] input_62;
    input [4:0] input_63;
    input [5:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      6'b110111 : begin
        result = input_55;
      end
      6'b111000 : begin
        result = input_56;
      end
      6'b111001 : begin
        result = input_57;
      end
      6'b111010 : begin
        result = input_58;
      end
      6'b111011 : begin
        result = input_59;
      end
      6'b111100 : begin
        result = input_60;
      end
      6'b111101 : begin
        result = input_61;
      end
      6'b111110 : begin
        result = input_62;
      end
      default : begin
        result = input_63;
      end
    endcase
    MUX_v_5_64_2 = result;
  end
  endfunction


  function automatic [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input  sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input  sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_32_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [7:0] input_2;
    input [7:0] input_3;
    input [7:0] input_4;
    input [7:0] input_5;
    input [7:0] input_6;
    input [7:0] input_7;
    input [7:0] input_8;
    input [7:0] input_9;
    input [7:0] input_10;
    input [7:0] input_11;
    input [7:0] input_12;
    input [7:0] input_13;
    input [7:0] input_14;
    input [7:0] input_15;
    input [7:0] input_16;
    input [7:0] input_17;
    input [7:0] input_18;
    input [7:0] input_19;
    input [7:0] input_20;
    input [7:0] input_21;
    input [7:0] input_22;
    input [7:0] input_23;
    input [7:0] input_24;
    input [7:0] input_25;
    input [7:0] input_26;
    input [7:0] input_27;
    input [7:0] input_28;
    input [7:0] input_29;
    input [7:0] input_30;
    input [7:0] input_31;
    input [4:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      5'b00000 : begin
        result = input_0;
      end
      5'b00001 : begin
        result = input_1;
      end
      5'b00010 : begin
        result = input_2;
      end
      5'b00011 : begin
        result = input_3;
      end
      5'b00100 : begin
        result = input_4;
      end
      5'b00101 : begin
        result = input_5;
      end
      5'b00110 : begin
        result = input_6;
      end
      5'b00111 : begin
        result = input_7;
      end
      5'b01000 : begin
        result = input_8;
      end
      5'b01001 : begin
        result = input_9;
      end
      5'b01010 : begin
        result = input_10;
      end
      5'b01011 : begin
        result = input_11;
      end
      5'b01100 : begin
        result = input_12;
      end
      5'b01101 : begin
        result = input_13;
      end
      5'b01110 : begin
        result = input_14;
      end
      5'b01111 : begin
        result = input_15;
      end
      5'b10000 : begin
        result = input_16;
      end
      5'b10001 : begin
        result = input_17;
      end
      5'b10010 : begin
        result = input_18;
      end
      5'b10011 : begin
        result = input_19;
      end
      5'b10100 : begin
        result = input_20;
      end
      5'b10101 : begin
        result = input_21;
      end
      5'b10110 : begin
        result = input_22;
      end
      5'b10111 : begin
        result = input_23;
      end
      5'b11000 : begin
        result = input_24;
      end
      5'b11001 : begin
        result = input_25;
      end
      5'b11010 : begin
        result = input_26;
      end
      5'b11011 : begin
        result = input_27;
      end
      5'b11100 : begin
        result = input_28;
      end
      5'b11101 : begin
        result = input_29;
      end
      5'b11110 : begin
        result = input_30;
      end
      default : begin
        result = input_31;
      end
    endcase
    MUX_v_8_32_2 = result;
  end
  endfunction


  function automatic [24:0] readslicef_26_25_1;
    input [25:0] vector;
    reg [25:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_26_25_1 = tmp[24:0];
  end
  endfunction


  function automatic [31:0] signext_32_1;
    input  vector;
  begin
    signext_32_1= {{31{vector}}, vector};
  end
  endfunction


  function automatic [2:0] signext_3_1;
    input  vector;
  begin
    signext_3_1= {{2{vector}}, vector};
  end
  endfunction


  function automatic [3:0] signext_4_3;
    input [2:0] vector;
  begin
    signext_4_3= {{1{vector[2]}}, vector};
  end
  endfunction


  function automatic [4:0] signext_5_1;
    input  vector;
  begin
    signext_5_1= {{4{vector}}, vector};
  end
  endfunction


  function automatic [4:0] signext_5_2;
    input [1:0] vector;
  begin
    signext_5_2= {{3{vector[1]}}, vector};
  end
  endfunction


  function automatic [4:0] conv_s2u_2_5 ;
    input [1:0]  vector ;
  begin
    conv_s2u_2_5 = {{3{vector[1]}}, vector};
  end
  endfunction


  function automatic [3:0] conv_u2s_3_4 ;
    input [2:0]  vector ;
  begin
    conv_u2s_3_4 =  {1'b0, vector};
  end
  endfunction


  function automatic [5:0] conv_u2s_5_6 ;
    input [4:0]  vector ;
  begin
    conv_u2s_5_6 =  {1'b0, vector};
  end
  endfunction


  function automatic [6:0] conv_u2s_6_7 ;
    input [5:0]  vector ;
  begin
    conv_u2s_6_7 =  {1'b0, vector};
  end
  endfunction


  function automatic [8:0] conv_u2s_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2s_8_9 =  {1'b0, vector};
  end
  endfunction


  function automatic [4:0] conv_u2u_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2u_4_5 = {1'b0, vector};
  end
  endfunction


  function automatic [25:0] conv_u2u_25_26 ;
    input [24:0]  vector ;
  begin
    conv_u2u_25_26 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ActUnit
// ------------------------------------------------------------------


module ActUnit (
  clk, rst, start_vld, start_rdy, start_dat, act_port_vld, act_port_rdy, act_port_dat,
      rva_in_vld, rva_in_rdy, rva_in_dat, rva_out_vld, rva_out_rdy, rva_out_dat,
      output_port_vld, output_port_rdy, output_port_dat, done_vld, done_rdy, done_dat
);
  input clk;
  input rst;
  input start_vld;
  output start_rdy;
  input start_dat;
  input act_port_vld;
  output act_port_rdy;
  input [511:0] act_port_dat;
  input rva_in_vld;
  output rva_in_rdy;
  input [600:0] rva_in_dat;
  output rva_out_vld;
  input rva_out_rdy;
  output [511:0] rva_out_dat;
  output output_port_vld;
  input output_port_rdy;
  output [521:0] output_port_dat;
  output done_vld;
  input done_rdy;
  output done_dat;



  // Interconnect Declarations for Component Instantiations 
  ActUnit_ActUnit_ActUnitRun ActUnit_ActUnitRun_inst (
      .clk(clk),
      .rst(rst),
      .start_vld(start_vld),
      .start_rdy(start_rdy),
      .start_dat(start_dat),
      .act_port_vld(act_port_vld),
      .act_port_rdy(act_port_rdy),
      .act_port_dat(act_port_dat),
      .rva_in_vld(rva_in_vld),
      .rva_in_rdy(rva_in_rdy),
      .rva_in_dat(rva_in_dat),
      .rva_out_vld(rva_out_vld),
      .rva_out_rdy(rva_out_rdy),
      .rva_out_dat(rva_out_dat),
      .output_port_vld(output_port_vld),
      .output_port_rdy(output_port_rdy),
      .output_port_dat(output_port_dat),
      .done_vld(done_vld),
      .done_rdy(done_rdy),
      .done_dat(done_dat)
    );
endmodule



