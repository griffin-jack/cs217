
//------> ./counter_top_Connections_InBlockingless_NVUINT32comma_Connections_SYN_PORTgreater_Pop_mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module counter_top_Connections_InBlockingless_NVUINT32comma_Connections_SYN_PORTgreater_Pop_mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ./counter_top_Connections_InBlockingless_NVUINT32comma_Connections_SYN_PORTgreater_Pop_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module counter_top_Connections_InBlockingless_NVUINT32comma_Connections_SYN_PORTgreater_Pop_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./counter_top_Connections_InBlockingless_NVUINT32comma_Connections_SYN_PORTgreater_Pop_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module counter_top_Connections_InBlockingless_NVUINT32comma_Connections_SYN_PORTgreater_Pop_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./counter_top_Connections_InBlockingless_NVUINT32comma_Connections_SYN_PORTgreater_Pop.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   code@rice-02
//  Generated date: Sat Jan 10 19:43:05 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlockingless_NVUINT32comma_Connections_SYN_PORTgreater_Pop_Connections_InBlocking_NVUINT32_Connections_SYN_PORT_Pop_core
// ------------------------------------------------------------------


module counter_top_Connections_InBlockingless_NVUINT32comma_Connections_SYN_PORTgreater_Pop_Connections_InBlocking_NVUINT32_Connections_SYN_PORT_Pop_core
    (
  this_vld, this_rdy, this_dat, return_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  reg this_rdy;
  input [31:0] this_dat;
  output [31:0] return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_3_cse;
  wire this_rdy_mx0c1;


  // Interconnect Declarations for Component Instantiations
  wire  nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_vld;
  counter_top_Connections_InBlockingless_NVUINT32comma_Connections_SYN_PORTgreater_Pop_mgc_out_dreg_v2
      #(.rscid(32'sd3),
  .width(32'sd32)) return_rsci (
      .d(this_dat),
      .z(return_rsc_z)
    );
  counter_top_Connections_InBlockingless_NVUINT32comma_Connections_SYN_PORTgreater_Pop_ccs_in_v1
      #(.rscid(32'sd13),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  counter_top_Connections_InBlockingless_NVUINT32comma_Connections_SYN_PORTgreater_Pop_ccs_sync_out_vld_v1
      #(.rscid(32'sd17)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld)
    );
  assign or_3_cse = ccs_ccore_start_rsci_idat | (io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & (~ this_vld));
  assign this_rdy_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_vld
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( or_3_cse | this_rdy_mx0c1 ) begin
      this_rdy <= ~ this_rdy_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_3_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_NVUINT32_Connections_SYN_PORT_Pop
// ------------------------------------------------------------------


module counter_top_Connections_InBlocking_NVUINT32_Connections_SYN_PORT_Pop (
  this_vld, this_rdy, this_dat, return_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  input [31:0] this_dat;
  output [31:0] return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  counter_top_Connections_InBlockingless_NVUINT32comma_Connections_SYN_PORTgreater_Pop_Connections_InBlocking_NVUINT32_Connections_SYN_PORT_Pop_core
      Connections_InBlocking_NVUINT32_Connections_SYN_PORT_Pop_core_inst (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./counter_top_Connections_OutBlockingless_NVUINT32comma_Connections_SYN_PORTgreater_Push_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module counter_top_Connections_OutBlockingless_NVUINT32comma_Connections_SYN_PORTgreater_Push_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./counter_top_Connections_OutBlockingless_NVUINT32comma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module counter_top_Connections_OutBlockingless_NVUINT32comma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./counter_top_Connections_OutBlockingless_NVUINT32comma_Connections_SYN_PORTgreater_Push.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   code@rice-02
//  Generated date: Sat Jan 10 19:43:03 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlockingless_NVUINT32comma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_NVUINT32_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module counter_top_Connections_OutBlockingless_NVUINT32comma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_NVUINT32_Connections_SYN_PORT_Push_core
    (
  this_vld, this_rdy, this_dat, m_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  reg this_vld;
  input this_rdy;
  output [31:0] this_dat;
  reg [31:0] this_dat;
  input [31:0] m_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire [31:0] m_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  wire and_dcpl;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_4_cse;
  wire this_vld_mx0c1;


  // Interconnect Declarations for Component Instantiations
  wire  nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  counter_top_Connections_OutBlockingless_NVUINT32comma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd1),
  .width(32'sd32)) m_rsci (
      .dat(m_rsc_dat),
      .idat(m_rsci_idat)
    );
  counter_top_Connections_OutBlockingless_NVUINT32comma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd14),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  counter_top_Connections_OutBlockingless_NVUINT32comma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1
      #(.rscid(32'sd18)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld)
    );
  assign or_4_cse = ccs_ccore_start_rsci_idat | and_dcpl;
  assign and_dcpl = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_rdy);
  assign this_vld_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_vld <= 1'b0;
    end
    else if ( or_4_cse | this_vld_mx0c1 ) begin
      this_vld <= ~ this_vld_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_dat <= 32'b00000000000000000000000000000000;
    end
    else if ( ~(and_dcpl | (~ ccs_ccore_start_rsci_idat)) ) begin
      this_dat <= m_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_4_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_NVUINT32_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module counter_top_Connections_OutBlocking_NVUINT32_Connections_SYN_PORT_Push (
  this_vld, this_rdy, this_dat, m_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  input this_rdy;
  output [31:0] this_dat;
  input [31:0] m_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  counter_top_Connections_OutBlockingless_NVUINT32comma_Connections_SYN_PORTgreater_Push_Connections_OutBlocking_NVUINT32_Connections_SYN_PORT_Push_core
      Connections_OutBlocking_NVUINT32_Connections_SYN_PORT_Push_core_inst (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .m_rsc_dat(m_rsc_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./counter_top_Connections_Combinationalless_NVUINT32comma_Connections_SYN_PORTgreater_Pop_mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module counter_top_Connections_Combinationalless_NVUINT32comma_Connections_SYN_PORTgreater_Pop_mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ./counter_top_Connections_Combinationalless_NVUINT32comma_Connections_SYN_PORTgreater_Pop_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module counter_top_Connections_Combinationalless_NVUINT32comma_Connections_SYN_PORTgreater_Pop_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./counter_top_Connections_Combinationalless_NVUINT32comma_Connections_SYN_PORTgreater_Pop_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module counter_top_Connections_Combinationalless_NVUINT32comma_Connections_SYN_PORTgreater_Pop_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./counter_top_Connections_Combinationalless_NVUINT32comma_Connections_SYN_PORTgreater_Pop.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   code@rice-02
//  Generated date: Sat Jan 10 19:43:01 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_Combinationalless_NVUINT32comma_Connections_SYN_PORTgreater_Pop_Connections_Combinational_NVUINT32_Connections_SYN_PORT_Pop_core
// ------------------------------------------------------------------


module counter_top_Connections_Combinationalless_NVUINT32comma_Connections_SYN_PORTgreater_Pop_Connections_Combinational_NVUINT32_Connections_SYN_PORT_Pop_core
    (
  this_vld, this_rdy, this_dat, return_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  reg this_rdy;
  input [31:0] this_dat;
  output [31:0] return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_3_cse;
  wire this_rdy_mx0c1;


  // Interconnect Declarations for Component Instantiations
  wire  nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_vld;
  counter_top_Connections_Combinationalless_NVUINT32comma_Connections_SYN_PORTgreater_Pop_mgc_out_dreg_v2
      #(.rscid(32'sd6),
  .width(32'sd32)) return_rsci (
      .d(this_dat),
      .z(return_rsc_z)
    );
  counter_top_Connections_Combinationalless_NVUINT32comma_Connections_SYN_PORTgreater_Pop_ccs_in_v1
      #(.rscid(32'sd12),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  counter_top_Connections_Combinationalless_NVUINT32comma_Connections_SYN_PORTgreater_Pop_ccs_sync_out_vld_v1
      #(.rscid(32'sd16)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld)
    );
  assign or_3_cse = ccs_ccore_start_rsci_idat | (io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & (~ this_vld));
  assign this_rdy_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_vld
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( or_3_cse | this_rdy_mx0c1 ) begin
      this_rdy <= ~ this_rdy_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_3_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_Combinational_NVUINT32_Connections_SYN_PORT_Pop
// ------------------------------------------------------------------


module counter_top_Connections_Combinational_NVUINT32_Connections_SYN_PORT_Pop (
  this_vld, this_rdy, this_dat, return_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_vld;
  output this_rdy;
  input [31:0] this_dat;
  output [31:0] return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  counter_top_Connections_Combinationalless_NVUINT32comma_Connections_SYN_PORTgreater_Pop_Connections_Combinational_NVUINT32_Connections_SYN_PORT_Pop_core
      Connections_Combinational_NVUINT32_Connections_SYN_PORT_Pop_core_inst (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./counter_top_Connections_Combinationalless_NVUINT32comma_Connections_SYN_PORTgreater_Push_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module counter_top_Connections_Combinationalless_NVUINT32comma_Connections_SYN_PORTgreater_Push_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./counter_top_Connections_Combinationalless_NVUINT32comma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module counter_top_Connections_Combinationalless_NVUINT32comma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./counter_top_Connections_Combinationalless_NVUINT32comma_Connections_SYN_PORTgreater_Push.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
//
//  Generated by:   code@rice-02
//  Generated date: Sat Jan 10 19:42:59 2026
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    Connections_Combinationalless_NVUINT32comma_Connections_SYN_PORTgreater_Push_Connections_Combinational_NVUINT32_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module counter_top_Connections_Combinationalless_NVUINT32comma_Connections_SYN_PORTgreater_Push_Connections_Combinational_NVUINT32_Connections_SYN_PORT_Push_core
    (
  this_vld, this_rdy, this_dat, m_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  reg this_vld;
  input this_rdy;
  output [31:0] this_dat;
  reg [31:0] this_dat;
  input [31:0] m_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire [31:0] m_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  wire and_dcpl;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_4_cse;
  wire this_vld_mx0c1;


  // Interconnect Declarations for Component Instantiations
  wire  nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  counter_top_Connections_Combinationalless_NVUINT32comma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd7),
  .width(32'sd32)) m_rsci (
      .dat(m_rsc_dat),
      .idat(m_rsci_idat)
    );
  counter_top_Connections_Combinationalless_NVUINT32comma_Connections_SYN_PORTgreater_Push_ccs_in_v1
      #(.rscid(32'sd11),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  counter_top_Connections_Combinationalless_NVUINT32comma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1
      #(.rscid(32'sd15)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld)
    );
  assign or_4_cse = ccs_ccore_start_rsci_idat | and_dcpl;
  assign and_dcpl = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_rdy);
  assign this_vld_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_vld <= 1'b0;
    end
    else if ( or_4_cse | this_vld_mx0c1 ) begin
      this_vld <= ~ this_vld_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_dat <= 32'b00000000000000000000000000000000;
    end
    else if ( ~(and_dcpl | (~ ccs_ccore_start_rsci_idat)) ) begin
      this_dat <= m_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_4_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_Combinational_NVUINT32_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module counter_top_Connections_Combinational_NVUINT32_Connections_SYN_PORT_Push (
  this_vld, this_rdy, this_dat, m_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_vld;
  input this_rdy;
  output [31:0] this_dat;
  input [31:0] m_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations
  counter_top_Connections_Combinationalless_NVUINT32comma_Connections_SYN_PORTgreater_Push_Connections_Combinational_NVUINT32_Connections_SYN_PORT_Push_core
      Connections_Combinational_NVUINT32_Connections_SYN_PORT_Push_core_inst (
      .this_vld(this_vld),
      .this_rdy(this_rdy),
      .this_dat(this_dat),
      .m_rsc_dat(m_rsc_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./counter_top.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.2_1/1143609 Production Release
//  HLS Date:       Wed Nov 13 18:57:31 PST 2024
// 
//  Generated by:   code@rice-01
//  Generated date: Sun Jan 11 13:03:22 2026
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    counter_top_counter_top_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module counter_top_counter_top_run_run_fsm (
  clk, rst, run_wen, fsm_output
);
  input clk;
  input rst;
  input run_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for counter_top_counter_top_run_run_fsm_1
  parameter
    run_rlp_C_0 = 2'd0,
    while_C_0 = 2'd1,
    while_C_1 = 2'd2,
    while_C_2 = 2'd3;

  reg [1:0] state_var;
  reg [1:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : counter_top_counter_top_run_run_fsm_1
    case (state_var)
      while_C_0 : begin
        fsm_output = 2'b01;
        state_var_NS = while_C_1;
      end
      while_C_1 : begin
        fsm_output = 2'b10;
        state_var_NS = while_C_2;
      end
      while_C_2 : begin
        fsm_output = 2'b11;
        state_var_NS = while_C_0;
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 2'b00;
        state_var_NS = while_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    counter_top_counter_top_run_staller
// ------------------------------------------------------------------


module counter_top_counter_top_run_staller (
  run_wen, counter_module_out_Pop_mioi_wen_comp, counter_in_Push_mioi_wen_comp, add_to_top_Pop_mioi_wen_comp
);
  output run_wen;
  input counter_module_out_Pop_mioi_wen_comp;
  input counter_in_Push_mioi_wen_comp;
  input add_to_top_Pop_mioi_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = counter_module_out_Pop_mioi_wen_comp & counter_in_Push_mioi_wen_comp
      & add_to_top_Pop_mioi_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    counter_top_counter_top_run_add_to_top_Pop_mioi_add_to_top_Pop_mio_wait_dp
// ------------------------------------------------------------------


module counter_top_counter_top_run_add_to_top_Pop_mioi_add_to_top_Pop_mio_wait_dp
    (
  clk, rst, add_to_top_Pop_mioi_oswt, add_to_top_Pop_mioi_wen_comp, add_to_top_Pop_mioi_return_rsc_z_mxwt,
      add_to_top_Pop_mioi_biwt, add_to_top_Pop_mioi_bdwt, add_to_top_Pop_mioi_bcwt,
      add_to_top_Pop_mioi_return_rsc_z
);
  input clk;
  input rst;
  input add_to_top_Pop_mioi_oswt;
  output add_to_top_Pop_mioi_wen_comp;
  output [31:0] add_to_top_Pop_mioi_return_rsc_z_mxwt;
  input add_to_top_Pop_mioi_biwt;
  input add_to_top_Pop_mioi_bdwt;
  output add_to_top_Pop_mioi_bcwt;
  reg add_to_top_Pop_mioi_bcwt;
  input [31:0] add_to_top_Pop_mioi_return_rsc_z;


  // Interconnect Declarations
  reg [31:0] add_to_top_Pop_mioi_return_rsc_z_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign add_to_top_Pop_mioi_wen_comp = (~ add_to_top_Pop_mioi_oswt) | add_to_top_Pop_mioi_biwt
      | add_to_top_Pop_mioi_bcwt;
  assign add_to_top_Pop_mioi_return_rsc_z_mxwt = MUX_v_32_2_2(add_to_top_Pop_mioi_return_rsc_z,
      add_to_top_Pop_mioi_return_rsc_z_bfwt, add_to_top_Pop_mioi_bcwt);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      add_to_top_Pop_mioi_bcwt <= 1'b0;
    end
    else begin
      add_to_top_Pop_mioi_bcwt <= ~((~(add_to_top_Pop_mioi_bcwt | add_to_top_Pop_mioi_biwt))
          | add_to_top_Pop_mioi_bdwt);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      add_to_top_Pop_mioi_return_rsc_z_bfwt <= 32'b00000000000000000000000000000000;
    end
    else if ( add_to_top_Pop_mioi_biwt ) begin
      add_to_top_Pop_mioi_return_rsc_z_bfwt <= add_to_top_Pop_mioi_return_rsc_z;
    end
  end

  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input  sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    counter_top_counter_top_run_add_to_top_Pop_mioi_add_to_top_Pop_mio_wait_ctrl
// ------------------------------------------------------------------


module counter_top_counter_top_run_add_to_top_Pop_mioi_add_to_top_Pop_mio_wait_ctrl
    (
  run_wen, add_to_top_Pop_mioi_oswt, add_to_top_Pop_mioi_biwt, add_to_top_Pop_mioi_bdwt,
      add_to_top_Pop_mioi_bcwt, add_to_top_Pop_mioi_ccs_ccore_start_rsc_dat_run_sct,
      add_to_top_Pop_mioi_ccs_ccore_done_sync_vld, add_to_top_Pop_mioi_oswt_pff
);
  input run_wen;
  input add_to_top_Pop_mioi_oswt;
  output add_to_top_Pop_mioi_biwt;
  output add_to_top_Pop_mioi_bdwt;
  input add_to_top_Pop_mioi_bcwt;
  output add_to_top_Pop_mioi_ccs_ccore_start_rsc_dat_run_sct;
  input add_to_top_Pop_mioi_ccs_ccore_done_sync_vld;
  input add_to_top_Pop_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign add_to_top_Pop_mioi_bdwt = add_to_top_Pop_mioi_oswt & run_wen;
  assign add_to_top_Pop_mioi_biwt = add_to_top_Pop_mioi_oswt & (~ add_to_top_Pop_mioi_bcwt)
      & add_to_top_Pop_mioi_ccs_ccore_done_sync_vld;
  assign add_to_top_Pop_mioi_ccs_ccore_start_rsc_dat_run_sct = run_wen & add_to_top_Pop_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    counter_top_counter_top_run_counter_in_Push_mioi_counter_in_Push_mio_wait_dp
// ------------------------------------------------------------------


module counter_top_counter_top_run_counter_in_Push_mioi_counter_in_Push_mio_wait_dp
    (
  clk, rst, counter_in_Push_mioi_oswt, counter_in_Push_mioi_wen_comp, counter_in_Push_mioi_biwt,
      counter_in_Push_mioi_bdwt, counter_in_Push_mioi_bcwt
);
  input clk;
  input rst;
  input counter_in_Push_mioi_oswt;
  output counter_in_Push_mioi_wen_comp;
  input counter_in_Push_mioi_biwt;
  input counter_in_Push_mioi_bdwt;
  output counter_in_Push_mioi_bcwt;
  reg counter_in_Push_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign counter_in_Push_mioi_wen_comp = (~ counter_in_Push_mioi_oswt) | counter_in_Push_mioi_biwt
      | counter_in_Push_mioi_bcwt;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      counter_in_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      counter_in_Push_mioi_bcwt <= ~((~(counter_in_Push_mioi_bcwt | counter_in_Push_mioi_biwt))
          | counter_in_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    counter_top_counter_top_run_counter_in_Push_mioi_counter_in_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module counter_top_counter_top_run_counter_in_Push_mioi_counter_in_Push_mio_wait_ctrl
    (
  run_wen, counter_in_Push_mioi_oswt, counter_in_Push_mioi_biwt, counter_in_Push_mioi_bdwt,
      counter_in_Push_mioi_bcwt, counter_in_Push_mioi_ccs_ccore_start_rsc_dat_run_sct,
      counter_in_Push_mioi_ccs_ccore_done_sync_vld, counter_in_Push_mioi_oswt_pff
);
  input run_wen;
  input counter_in_Push_mioi_oswt;
  output counter_in_Push_mioi_biwt;
  output counter_in_Push_mioi_bdwt;
  input counter_in_Push_mioi_bcwt;
  output counter_in_Push_mioi_ccs_ccore_start_rsc_dat_run_sct;
  input counter_in_Push_mioi_ccs_ccore_done_sync_vld;
  input counter_in_Push_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign counter_in_Push_mioi_bdwt = counter_in_Push_mioi_oswt & run_wen;
  assign counter_in_Push_mioi_biwt = counter_in_Push_mioi_oswt & (~ counter_in_Push_mioi_bcwt)
      & counter_in_Push_mioi_ccs_ccore_done_sync_vld;
  assign counter_in_Push_mioi_ccs_ccore_start_rsc_dat_run_sct = run_wen & counter_in_Push_mioi_oswt_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    counter_top_counter_top_run_counter_module_out_Pop_mioi_counter_module_out_Pop_mio_wait_ctrl
// ------------------------------------------------------------------


module counter_top_counter_top_run_counter_module_out_Pop_mioi_counter_module_out_Pop_mio_wait_ctrl
    (
  run_wten, counter_module_out_Pop_mioi_iswt0, counter_module_out_Pop_mioi_biwt,
      counter_module_out_Pop_mioi_ccs_ccore_start_rsc_dat_run_sct, counter_module_out_Pop_mioi_ccs_ccore_done_sync_vld,
      counter_module_out_Pop_mioi_iswt0_pff
);
  input run_wten;
  input counter_module_out_Pop_mioi_iswt0;
  output counter_module_out_Pop_mioi_biwt;
  output counter_module_out_Pop_mioi_ccs_ccore_start_rsc_dat_run_sct;
  input counter_module_out_Pop_mioi_ccs_ccore_done_sync_vld;
  input counter_module_out_Pop_mioi_iswt0_pff;



  // Interconnect Declarations for Component Instantiations 
  assign counter_module_out_Pop_mioi_biwt = counter_module_out_Pop_mioi_iswt0 & counter_module_out_Pop_mioi_ccs_ccore_done_sync_vld;
  assign counter_module_out_Pop_mioi_ccs_ccore_start_rsc_dat_run_sct = (~ run_wten)
      & counter_module_out_Pop_mioi_iswt0_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    counter_top_counter_module_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module counter_top_counter_module_run_run_fsm (
  clk, rst, counter_out_Push_mioi_wen_comp, fsm_output
);
  input clk;
  input rst;
  input counter_out_Push_mioi_wen_comp;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for counter_top_counter_module_run_run_fsm_1
  parameter
    run_rlp_C_0 = 2'd0,
    while_C_0 = 2'd1,
    while_C_1 = 2'd2;

  reg [1:0] state_var;
  reg [1:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : counter_top_counter_module_run_run_fsm_1
    case (state_var)
      while_C_0 : begin
        fsm_output = 2'b01;
        state_var_NS = while_C_1;
      end
      while_C_1 : begin
        fsm_output = 2'b10;
        state_var_NS = while_C_0;
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 2'b00;
        state_var_NS = while_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( counter_out_Push_mioi_wen_comp ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    counter_top_counter_module_run_staller
// ------------------------------------------------------------------


module counter_top_counter_module_run_staller (
  run_wten, counter_out_Push_mioi_wen_comp
);
  output run_wten;
  input counter_out_Push_mioi_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wten = ~ counter_out_Push_mioi_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    counter_top_counter_module_run_counter_out_Push_mioi_counter_out_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module counter_top_counter_module_run_counter_out_Push_mioi_counter_out_Push_mio_wait_ctrl
    (
  run_wten, counter_out_Push_mioi_iswt0, counter_out_Push_mioi_biwt, counter_out_Push_mioi_ccs_ccore_start_rsc_dat_run_sct,
      counter_out_Push_mioi_ccs_ccore_done_sync_vld, counter_out_Push_mioi_iswt0_pff
);
  input run_wten;
  input counter_out_Push_mioi_iswt0;
  output counter_out_Push_mioi_biwt;
  output counter_out_Push_mioi_ccs_ccore_start_rsc_dat_run_sct;
  input counter_out_Push_mioi_ccs_ccore_done_sync_vld;
  input counter_out_Push_mioi_iswt0_pff;



  // Interconnect Declarations for Component Instantiations 
  assign counter_out_Push_mioi_biwt = counter_out_Push_mioi_iswt0 & counter_out_Push_mioi_ccs_ccore_done_sync_vld;
  assign counter_out_Push_mioi_ccs_ccore_start_rsc_dat_run_sct = (~ run_wten) & counter_out_Push_mioi_iswt0_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    counter_top_add_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module counter_top_add_run_run_fsm (
  clk, rst, run_wen, fsm_output
);
  input clk;
  input rst;
  input run_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for counter_top_add_run_run_fsm_1
  parameter
    run_rlp_C_0 = 2'd0,
    while_C_0 = 2'd1,
    while_C_1 = 2'd2,
    while_C_2 = 2'd3;

  reg [1:0] state_var;
  reg [1:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : counter_top_add_run_run_fsm_1
    case (state_var)
      while_C_0 : begin
        fsm_output = 2'b01;
        state_var_NS = while_C_1;
      end
      while_C_1 : begin
        fsm_output = 2'b10;
        state_var_NS = while_C_2;
      end
      while_C_2 : begin
        fsm_output = 2'b11;
        state_var_NS = while_C_0;
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 2'b00;
        state_var_NS = while_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    counter_top_add_run_staller
// ------------------------------------------------------------------


module counter_top_add_run_staller (
  run_wen, counter_in_Pop_mioi_wen_comp, add_out_Push_mioi_wen_comp
);
  output run_wen;
  input counter_in_Pop_mioi_wen_comp;
  input add_out_Push_mioi_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = counter_in_Pop_mioi_wen_comp & add_out_Push_mioi_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    counter_top_add_run_add_out_Push_mioi_add_out_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module counter_top_add_run_add_out_Push_mioi_add_out_Push_mio_wait_ctrl (
  run_wten, add_out_Push_mioi_iswt0, add_out_Push_mioi_biwt, add_out_Push_mioi_ccs_ccore_start_rsc_dat_run_sct,
      add_out_Push_mioi_ccs_ccore_done_sync_vld, add_out_Push_mioi_iswt0_pff
);
  input run_wten;
  input add_out_Push_mioi_iswt0;
  output add_out_Push_mioi_biwt;
  output add_out_Push_mioi_ccs_ccore_start_rsc_dat_run_sct;
  input add_out_Push_mioi_ccs_ccore_done_sync_vld;
  input add_out_Push_mioi_iswt0_pff;



  // Interconnect Declarations for Component Instantiations 
  assign add_out_Push_mioi_biwt = add_out_Push_mioi_iswt0 & add_out_Push_mioi_ccs_ccore_done_sync_vld;
  assign add_out_Push_mioi_ccs_ccore_start_rsc_dat_run_sct = (~ run_wten) & add_out_Push_mioi_iswt0_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    counter_top_add_run_counter_in_Pop_mioi_counter_in_Pop_mio_wait_ctrl
// ------------------------------------------------------------------


module counter_top_add_run_counter_in_Pop_mioi_counter_in_Pop_mio_wait_ctrl (
  run_wten, counter_in_Pop_mioi_iswt0, counter_in_Pop_mioi_biwt, counter_in_Pop_mioi_ccs_ccore_start_rsc_dat_run_sct,
      counter_in_Pop_mioi_ccs_ccore_done_sync_vld, counter_in_Pop_mioi_iswt0_pff
);
  input run_wten;
  input counter_in_Pop_mioi_iswt0;
  output counter_in_Pop_mioi_biwt;
  output counter_in_Pop_mioi_ccs_ccore_start_rsc_dat_run_sct;
  input counter_in_Pop_mioi_ccs_ccore_done_sync_vld;
  input counter_in_Pop_mioi_iswt0_pff;



  // Interconnect Declarations for Component Instantiations 
  assign counter_in_Pop_mioi_biwt = counter_in_Pop_mioi_iswt0 & counter_in_Pop_mioi_ccs_ccore_done_sync_vld;
  assign counter_in_Pop_mioi_ccs_ccore_start_rsc_dat_run_sct = (~ run_wten) & counter_in_Pop_mioi_iswt0_pff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    counter_top_counter_top_run_add_to_top_Pop_mioi
// ------------------------------------------------------------------


module counter_top_counter_top_run_add_to_top_Pop_mioi (
  clk, rst, add_to_top_vld, add_to_top_rdy, add_to_top_dat, run_wen, add_to_top_Pop_mioi_oswt,
      add_to_top_Pop_mioi_wen_comp, add_to_top_Pop_mioi_return_rsc_z_mxwt, add_to_top_Pop_mioi_oswt_pff
);
  input clk;
  input rst;
  input add_to_top_vld;
  output add_to_top_rdy;
  input [31:0] add_to_top_dat;
  input run_wen;
  input add_to_top_Pop_mioi_oswt;
  output add_to_top_Pop_mioi_wen_comp;
  output [31:0] add_to_top_Pop_mioi_return_rsc_z_mxwt;
  input add_to_top_Pop_mioi_oswt_pff;


  // Interconnect Declarations
  wire add_to_top_Pop_mioi_biwt;
  wire add_to_top_Pop_mioi_bdwt;
  wire add_to_top_Pop_mioi_bcwt;
  wire [31:0] add_to_top_Pop_mioi_return_rsc_z;
  wire add_to_top_Pop_mioi_ccs_ccore_start_rsc_dat_run_sct;
  wire add_to_top_Pop_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  counter_top_Connections_Combinational_NVUINT32_Connections_SYN_PORT_Pop  add_to_top_Pop_mioi
      (
      .this_vld(add_to_top_vld),
      .this_rdy(add_to_top_rdy),
      .this_dat(add_to_top_dat),
      .return_rsc_z(add_to_top_Pop_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(add_to_top_Pop_mioi_ccs_ccore_start_rsc_dat_run_sct),
      .ccs_ccore_done_sync_vld(add_to_top_Pop_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  counter_top_counter_top_run_add_to_top_Pop_mioi_add_to_top_Pop_mio_wait_ctrl counter_top_run_add_to_top_Pop_mioi_add_to_top_Pop_mio_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .add_to_top_Pop_mioi_oswt(add_to_top_Pop_mioi_oswt),
      .add_to_top_Pop_mioi_biwt(add_to_top_Pop_mioi_biwt),
      .add_to_top_Pop_mioi_bdwt(add_to_top_Pop_mioi_bdwt),
      .add_to_top_Pop_mioi_bcwt(add_to_top_Pop_mioi_bcwt),
      .add_to_top_Pop_mioi_ccs_ccore_start_rsc_dat_run_sct(add_to_top_Pop_mioi_ccs_ccore_start_rsc_dat_run_sct),
      .add_to_top_Pop_mioi_ccs_ccore_done_sync_vld(add_to_top_Pop_mioi_ccs_ccore_done_sync_vld),
      .add_to_top_Pop_mioi_oswt_pff(add_to_top_Pop_mioi_oswt_pff)
    );
  counter_top_counter_top_run_add_to_top_Pop_mioi_add_to_top_Pop_mio_wait_dp counter_top_run_add_to_top_Pop_mioi_add_to_top_Pop_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .add_to_top_Pop_mioi_oswt(add_to_top_Pop_mioi_oswt),
      .add_to_top_Pop_mioi_wen_comp(add_to_top_Pop_mioi_wen_comp),
      .add_to_top_Pop_mioi_return_rsc_z_mxwt(add_to_top_Pop_mioi_return_rsc_z_mxwt),
      .add_to_top_Pop_mioi_biwt(add_to_top_Pop_mioi_biwt),
      .add_to_top_Pop_mioi_bdwt(add_to_top_Pop_mioi_bdwt),
      .add_to_top_Pop_mioi_bcwt(add_to_top_Pop_mioi_bcwt),
      .add_to_top_Pop_mioi_return_rsc_z(add_to_top_Pop_mioi_return_rsc_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    counter_top_counter_top_run_counter_in_Push_mioi
// ------------------------------------------------------------------


module counter_top_counter_top_run_counter_in_Push_mioi (
  clk, rst, counter_in_vld, counter_in_rdy, counter_in_dat, run_wen, counter_in_Push_mioi_oswt,
      counter_in_Push_mioi_wen_comp, counter_in_Push_mioi_m_rsc_dat_run, counter_in_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output counter_in_vld;
  input counter_in_rdy;
  output [31:0] counter_in_dat;
  input run_wen;
  input counter_in_Push_mioi_oswt;
  output counter_in_Push_mioi_wen_comp;
  input [31:0] counter_in_Push_mioi_m_rsc_dat_run;
  input counter_in_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire counter_in_Push_mioi_biwt;
  wire counter_in_Push_mioi_bdwt;
  wire counter_in_Push_mioi_bcwt;
  wire counter_in_Push_mioi_ccs_ccore_start_rsc_dat_run_sct;
  wire counter_in_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  counter_top_Connections_Combinational_NVUINT32_Connections_SYN_PORT_Push  counter_in_Push_mioi
      (
      .this_vld(counter_in_vld),
      .this_rdy(counter_in_rdy),
      .this_dat(counter_in_dat),
      .m_rsc_dat(counter_in_Push_mioi_m_rsc_dat_run),
      .ccs_ccore_start_rsc_dat(counter_in_Push_mioi_ccs_ccore_start_rsc_dat_run_sct),
      .ccs_ccore_done_sync_vld(counter_in_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  counter_top_counter_top_run_counter_in_Push_mioi_counter_in_Push_mio_wait_ctrl
      counter_top_run_counter_in_Push_mioi_counter_in_Push_mio_wait_ctrl_inst (
      .run_wen(run_wen),
      .counter_in_Push_mioi_oswt(counter_in_Push_mioi_oswt),
      .counter_in_Push_mioi_biwt(counter_in_Push_mioi_biwt),
      .counter_in_Push_mioi_bdwt(counter_in_Push_mioi_bdwt),
      .counter_in_Push_mioi_bcwt(counter_in_Push_mioi_bcwt),
      .counter_in_Push_mioi_ccs_ccore_start_rsc_dat_run_sct(counter_in_Push_mioi_ccs_ccore_start_rsc_dat_run_sct),
      .counter_in_Push_mioi_ccs_ccore_done_sync_vld(counter_in_Push_mioi_ccs_ccore_done_sync_vld),
      .counter_in_Push_mioi_oswt_pff(counter_in_Push_mioi_oswt_pff)
    );
  counter_top_counter_top_run_counter_in_Push_mioi_counter_in_Push_mio_wait_dp counter_top_run_counter_in_Push_mioi_counter_in_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .counter_in_Push_mioi_oswt(counter_in_Push_mioi_oswt),
      .counter_in_Push_mioi_wen_comp(counter_in_Push_mioi_wen_comp),
      .counter_in_Push_mioi_biwt(counter_in_Push_mioi_biwt),
      .counter_in_Push_mioi_bdwt(counter_in_Push_mioi_bdwt),
      .counter_in_Push_mioi_bcwt(counter_in_Push_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    counter_top_counter_top_run_counter_module_out_Pop_mioi
// ------------------------------------------------------------------


module counter_top_counter_top_run_counter_module_out_Pop_mioi (
  clk, rst, counter_module_out_vld, counter_module_out_rdy, counter_module_out_dat,
      run_wten, counter_module_out_Pop_mioi_oswt, counter_module_out_Pop_mioi_wen_comp,
      counter_module_out_Pop_mioi_return_rsc_z_mxwt, counter_module_out_Pop_mioi_oswt_pff
);
  input clk;
  input rst;
  input counter_module_out_vld;
  output counter_module_out_rdy;
  input [31:0] counter_module_out_dat;
  input run_wten;
  input counter_module_out_Pop_mioi_oswt;
  output counter_module_out_Pop_mioi_wen_comp;
  output [31:0] counter_module_out_Pop_mioi_return_rsc_z_mxwt;
  input counter_module_out_Pop_mioi_oswt_pff;


  // Interconnect Declarations
  wire counter_module_out_Pop_mioi_biwt;
  wire [31:0] counter_module_out_Pop_mioi_return_rsc_z;
  wire counter_module_out_Pop_mioi_ccs_ccore_start_rsc_dat_run_sct;
  wire counter_module_out_Pop_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  counter_top_Connections_Combinational_NVUINT32_Connections_SYN_PORT_Pop  counter_module_out_Pop_mioi
      (
      .this_vld(counter_module_out_vld),
      .this_rdy(counter_module_out_rdy),
      .this_dat(counter_module_out_dat),
      .return_rsc_z(counter_module_out_Pop_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(counter_module_out_Pop_mioi_ccs_ccore_start_rsc_dat_run_sct),
      .ccs_ccore_done_sync_vld(counter_module_out_Pop_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  counter_top_counter_top_run_counter_module_out_Pop_mioi_counter_module_out_Pop_mio_wait_ctrl
      counter_top_run_counter_module_out_Pop_mioi_counter_module_out_Pop_mio_wait_ctrl_inst
      (
      .run_wten(run_wten),
      .counter_module_out_Pop_mioi_iswt0(counter_module_out_Pop_mioi_oswt),
      .counter_module_out_Pop_mioi_biwt(counter_module_out_Pop_mioi_biwt),
      .counter_module_out_Pop_mioi_ccs_ccore_start_rsc_dat_run_sct(counter_module_out_Pop_mioi_ccs_ccore_start_rsc_dat_run_sct),
      .counter_module_out_Pop_mioi_ccs_ccore_done_sync_vld(counter_module_out_Pop_mioi_ccs_ccore_done_sync_vld),
      .counter_module_out_Pop_mioi_iswt0_pff(counter_module_out_Pop_mioi_oswt_pff)
    );
  assign counter_module_out_Pop_mioi_return_rsc_z_mxwt = counter_module_out_Pop_mioi_return_rsc_z;
  assign counter_module_out_Pop_mioi_wen_comp = (~ counter_module_out_Pop_mioi_oswt)
      | counter_module_out_Pop_mioi_biwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    counter_top_counter_module_run_counter_out_Push_mioi
// ------------------------------------------------------------------


module counter_top_counter_module_run_counter_out_Push_mioi (
  clk, rst, counter_out_vld, counter_out_rdy, counter_out_dat, run_wten, counter_out_Push_mioi_oswt,
      counter_out_Push_mioi_wen_comp, counter_out_Push_mioi_m_rsc_dat_run, counter_out_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output counter_out_vld;
  input counter_out_rdy;
  output [31:0] counter_out_dat;
  input run_wten;
  input counter_out_Push_mioi_oswt;
  output counter_out_Push_mioi_wen_comp;
  input [31:0] counter_out_Push_mioi_m_rsc_dat_run;
  input counter_out_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire counter_out_Push_mioi_biwt;
  wire counter_out_Push_mioi_ccs_ccore_start_rsc_dat_run_sct;
  wire counter_out_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  counter_top_Connections_OutBlocking_NVUINT32_Connections_SYN_PORT_Push  counter_out_Push_mioi
      (
      .this_vld(counter_out_vld),
      .this_rdy(counter_out_rdy),
      .this_dat(counter_out_dat),
      .m_rsc_dat(counter_out_Push_mioi_m_rsc_dat_run),
      .ccs_ccore_start_rsc_dat(counter_out_Push_mioi_ccs_ccore_start_rsc_dat_run_sct),
      .ccs_ccore_done_sync_vld(counter_out_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  counter_top_counter_module_run_counter_out_Push_mioi_counter_out_Push_mio_wait_ctrl
      counter_module_run_counter_out_Push_mioi_counter_out_Push_mio_wait_ctrl_inst
      (
      .run_wten(run_wten),
      .counter_out_Push_mioi_iswt0(counter_out_Push_mioi_oswt),
      .counter_out_Push_mioi_biwt(counter_out_Push_mioi_biwt),
      .counter_out_Push_mioi_ccs_ccore_start_rsc_dat_run_sct(counter_out_Push_mioi_ccs_ccore_start_rsc_dat_run_sct),
      .counter_out_Push_mioi_ccs_ccore_done_sync_vld(counter_out_Push_mioi_ccs_ccore_done_sync_vld),
      .counter_out_Push_mioi_iswt0_pff(counter_out_Push_mioi_oswt_pff)
    );
  assign counter_out_Push_mioi_wen_comp = (~ counter_out_Push_mioi_oswt) | counter_out_Push_mioi_biwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    counter_top_add_run_add_out_Push_mioi
// ------------------------------------------------------------------


module counter_top_add_run_add_out_Push_mioi (
  clk, rst, add_out_vld, add_out_rdy, add_out_dat, run_wten, add_out_Push_mioi_oswt,
      add_out_Push_mioi_wen_comp, add_out_Push_mioi_m_rsc_dat_run, add_out_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output add_out_vld;
  input add_out_rdy;
  output [31:0] add_out_dat;
  input run_wten;
  input add_out_Push_mioi_oswt;
  output add_out_Push_mioi_wen_comp;
  input [31:0] add_out_Push_mioi_m_rsc_dat_run;
  input add_out_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire add_out_Push_mioi_biwt;
  wire add_out_Push_mioi_ccs_ccore_start_rsc_dat_run_sct;
  wire add_out_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  counter_top_Connections_OutBlocking_NVUINT32_Connections_SYN_PORT_Push  add_out_Push_mioi
      (
      .this_vld(add_out_vld),
      .this_rdy(add_out_rdy),
      .this_dat(add_out_dat),
      .m_rsc_dat(add_out_Push_mioi_m_rsc_dat_run),
      .ccs_ccore_start_rsc_dat(add_out_Push_mioi_ccs_ccore_start_rsc_dat_run_sct),
      .ccs_ccore_done_sync_vld(add_out_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  counter_top_add_run_add_out_Push_mioi_add_out_Push_mio_wait_ctrl add_run_add_out_Push_mioi_add_out_Push_mio_wait_ctrl_inst
      (
      .run_wten(run_wten),
      .add_out_Push_mioi_iswt0(add_out_Push_mioi_oswt),
      .add_out_Push_mioi_biwt(add_out_Push_mioi_biwt),
      .add_out_Push_mioi_ccs_ccore_start_rsc_dat_run_sct(add_out_Push_mioi_ccs_ccore_start_rsc_dat_run_sct),
      .add_out_Push_mioi_ccs_ccore_done_sync_vld(add_out_Push_mioi_ccs_ccore_done_sync_vld),
      .add_out_Push_mioi_iswt0_pff(add_out_Push_mioi_oswt_pff)
    );
  assign add_out_Push_mioi_wen_comp = (~ add_out_Push_mioi_oswt) | add_out_Push_mioi_biwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    counter_top_add_run_counter_in_Pop_mioi
// ------------------------------------------------------------------


module counter_top_add_run_counter_in_Pop_mioi (
  clk, rst, counter_in_vld, counter_in_rdy, counter_in_dat, run_wten, counter_in_Pop_mioi_oswt,
      counter_in_Pop_mioi_wen_comp, counter_in_Pop_mioi_return_rsc_z_mxwt, counter_in_Pop_mioi_oswt_pff
);
  input clk;
  input rst;
  input counter_in_vld;
  output counter_in_rdy;
  input [31:0] counter_in_dat;
  input run_wten;
  input counter_in_Pop_mioi_oswt;
  output counter_in_Pop_mioi_wen_comp;
  output [31:0] counter_in_Pop_mioi_return_rsc_z_mxwt;
  input counter_in_Pop_mioi_oswt_pff;


  // Interconnect Declarations
  wire counter_in_Pop_mioi_biwt;
  wire [31:0] counter_in_Pop_mioi_return_rsc_z;
  wire counter_in_Pop_mioi_ccs_ccore_start_rsc_dat_run_sct;
  wire counter_in_Pop_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  counter_top_Connections_InBlocking_NVUINT32_Connections_SYN_PORT_Pop  counter_in_Pop_mioi
      (
      .this_vld(counter_in_vld),
      .this_rdy(counter_in_rdy),
      .this_dat(counter_in_dat),
      .return_rsc_z(counter_in_Pop_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(counter_in_Pop_mioi_ccs_ccore_start_rsc_dat_run_sct),
      .ccs_ccore_done_sync_vld(counter_in_Pop_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst)
    );
  counter_top_add_run_counter_in_Pop_mioi_counter_in_Pop_mio_wait_ctrl add_run_counter_in_Pop_mioi_counter_in_Pop_mio_wait_ctrl_inst
      (
      .run_wten(run_wten),
      .counter_in_Pop_mioi_iswt0(counter_in_Pop_mioi_oswt),
      .counter_in_Pop_mioi_biwt(counter_in_Pop_mioi_biwt),
      .counter_in_Pop_mioi_ccs_ccore_start_rsc_dat_run_sct(counter_in_Pop_mioi_ccs_ccore_start_rsc_dat_run_sct),
      .counter_in_Pop_mioi_ccs_ccore_done_sync_vld(counter_in_Pop_mioi_ccs_ccore_done_sync_vld),
      .counter_in_Pop_mioi_iswt0_pff(counter_in_Pop_mioi_oswt_pff)
    );
  assign counter_in_Pop_mioi_return_rsc_z_mxwt = counter_in_Pop_mioi_return_rsc_z;
  assign counter_in_Pop_mioi_wen_comp = (~ counter_in_Pop_mioi_oswt) | counter_in_Pop_mioi_biwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    counter_top_counter_top_run
// ------------------------------------------------------------------


module counter_top_counter_top_run (
  clk, rst, counter_out, add_out, counter_module_out_vld, counter_module_out_rdy,
      counter_module_out_dat, counter_in_vld, counter_in_rdy, counter_in_dat, add_to_top_vld,
      add_to_top_rdy, add_to_top_dat
);
  input clk;
  input rst;
  output [31:0] counter_out;
  reg [31:0] counter_out;
  output [31:0] add_out;
  reg [31:0] add_out;
  input counter_module_out_vld;
  output counter_module_out_rdy;
  input [31:0] counter_module_out_dat;
  output counter_in_vld;
  input counter_in_rdy;
  output [31:0] counter_in_dat;
  input add_to_top_vld;
  output add_to_top_rdy;
  input [31:0] add_to_top_dat;


  // Interconnect Declarations
  wire run_wen;
  wire counter_module_out_Pop_mioi_wen_comp;
  wire [31:0] counter_module_out_Pop_mioi_return_rsc_z_mxwt;
  wire counter_in_Push_mioi_wen_comp;
  reg [31:0] counter_in_Push_mioi_m_rsc_dat_run;
  wire add_to_top_Pop_mioi_wen_comp;
  wire [31:0] add_to_top_Pop_mioi_return_rsc_z_mxwt;
  wire [1:0] fsm_output;
  reg reg_add_to_top_Pop_mioi_iswt0_cse;
  reg reg_counter_module_out_Pop_mioi_iswt0_cse;
  wire add_out_and_cse;
  wire and_1_rmff;
  wire and_rmff;
  reg reg_counter_in_Push_mioi_m_rsc_dat_run_enexo;
  wire counter_out_and_enex5;


  // Interconnect Declarations for Component Instantiations 
  wire  nl_counter_top_run_counter_module_out_Pop_mioi_inst_run_wten;
  assign nl_counter_top_run_counter_module_out_Pop_mioi_inst_run_wten = ~ run_wen;
  counter_top_counter_top_run_counter_module_out_Pop_mioi counter_top_run_counter_module_out_Pop_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .counter_module_out_vld(counter_module_out_vld),
      .counter_module_out_rdy(counter_module_out_rdy),
      .counter_module_out_dat(counter_module_out_dat),
      .run_wten(nl_counter_top_run_counter_module_out_Pop_mioi_inst_run_wten),
      .counter_module_out_Pop_mioi_oswt(reg_counter_module_out_Pop_mioi_iswt0_cse),
      .counter_module_out_Pop_mioi_wen_comp(counter_module_out_Pop_mioi_wen_comp),
      .counter_module_out_Pop_mioi_return_rsc_z_mxwt(counter_module_out_Pop_mioi_return_rsc_z_mxwt),
      .counter_module_out_Pop_mioi_oswt_pff(and_1_rmff)
    );
  counter_top_counter_top_run_counter_in_Push_mioi counter_top_run_counter_in_Push_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .counter_in_vld(counter_in_vld),
      .counter_in_rdy(counter_in_rdy),
      .counter_in_dat(counter_in_dat),
      .run_wen(run_wen),
      .counter_in_Push_mioi_oswt(reg_add_to_top_Pop_mioi_iswt0_cse),
      .counter_in_Push_mioi_wen_comp(counter_in_Push_mioi_wen_comp),
      .counter_in_Push_mioi_m_rsc_dat_run(counter_module_out_Pop_mioi_return_rsc_z_mxwt),
      .counter_in_Push_mioi_oswt_pff(and_rmff)
    );
  counter_top_counter_top_run_add_to_top_Pop_mioi counter_top_run_add_to_top_Pop_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .add_to_top_vld(add_to_top_vld),
      .add_to_top_rdy(add_to_top_rdy),
      .add_to_top_dat(add_to_top_dat),
      .run_wen(run_wen),
      .add_to_top_Pop_mioi_oswt(reg_add_to_top_Pop_mioi_iswt0_cse),
      .add_to_top_Pop_mioi_wen_comp(add_to_top_Pop_mioi_wen_comp),
      .add_to_top_Pop_mioi_return_rsc_z_mxwt(add_to_top_Pop_mioi_return_rsc_z_mxwt),
      .add_to_top_Pop_mioi_oswt_pff(and_rmff)
    );
  counter_top_counter_top_run_staller counter_top_run_staller_inst (
      .run_wen(run_wen),
      .counter_module_out_Pop_mioi_wen_comp(counter_module_out_Pop_mioi_wen_comp),
      .counter_in_Push_mioi_wen_comp(counter_in_Push_mioi_wen_comp),
      .add_to_top_Pop_mioi_wen_comp(add_to_top_Pop_mioi_wen_comp)
    );
  counter_top_counter_top_run_run_fsm counter_top_run_run_fsm_inst (
      .clk(clk),
      .rst(rst),
      .run_wen(run_wen),
      .fsm_output(fsm_output)
    );
  assign and_rmff = (fsm_output==2'b10);
  assign and_1_rmff = (fsm_output==2'b01);
  assign add_out_and_cse = run_wen & (fsm_output==2'b11);
  assign counter_out_and_enex5 = add_out_and_cse & reg_counter_in_Push_mioi_m_rsc_dat_run_enexo;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_add_to_top_Pop_mioi_iswt0_cse <= 1'b0;
      counter_in_Push_mioi_m_rsc_dat_run <= 32'b00000000000000000000000000000000;
      reg_counter_module_out_Pop_mioi_iswt0_cse <= 1'b0;
    end
    else if ( run_wen ) begin
      reg_add_to_top_Pop_mioi_iswt0_cse <= and_rmff;
      counter_in_Push_mioi_m_rsc_dat_run <= counter_module_out_Pop_mioi_return_rsc_z_mxwt;
      reg_counter_module_out_Pop_mioi_iswt0_cse <= and_1_rmff;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      add_out <= 32'b00000000000000000000000000000000;
    end
    else if ( add_out_and_cse ) begin
      add_out <= add_to_top_Pop_mioi_return_rsc_z_mxwt;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      counter_out <= 32'b00000000000000000000000000000000;
    end
    else if ( counter_out_and_enex5 ) begin
      counter_out <= counter_in_Push_mioi_m_rsc_dat_run;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_counter_in_Push_mioi_m_rsc_dat_run_enexo <= 1'b1;
    end
    else if ( run_wen | counter_out_and_enex5 ) begin
      reg_counter_in_Push_mioi_m_rsc_dat_run_enexo <= run_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    counter_top_counter_module_run
// ------------------------------------------------------------------


module counter_top_counter_module_run (
  clk, rst, counter_out_vld, counter_out_rdy, counter_out_dat
);
  input clk;
  input rst;
  output counter_out_vld;
  input counter_out_rdy;
  output [31:0] counter_out_dat;


  // Interconnect Declarations
  wire run_wten;
  wire counter_out_Push_mioi_wen_comp;
  wire [1:0] fsm_output;
  reg reg_counter_out_Push_mioi_iswt0_cse;
  wire and_rmff;
  wire [31:0] while_ac_int_cctor_sva_1;
  wire [32:0] nl_while_ac_int_cctor_sva_1;
  reg [31:0] counter_out_sig_sva;


  // Interconnect Declarations for Component Instantiations 
  counter_top_counter_module_run_counter_out_Push_mioi counter_module_run_counter_out_Push_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .counter_out_vld(counter_out_vld),
      .counter_out_rdy(counter_out_rdy),
      .counter_out_dat(counter_out_dat),
      .run_wten(run_wten),
      .counter_out_Push_mioi_oswt(reg_counter_out_Push_mioi_iswt0_cse),
      .counter_out_Push_mioi_wen_comp(counter_out_Push_mioi_wen_comp),
      .counter_out_Push_mioi_m_rsc_dat_run(while_ac_int_cctor_sva_1),
      .counter_out_Push_mioi_oswt_pff(and_rmff)
    );
  counter_top_counter_module_run_staller counter_module_run_staller_inst (
      .run_wten(run_wten),
      .counter_out_Push_mioi_wen_comp(counter_out_Push_mioi_wen_comp)
    );
  counter_top_counter_module_run_run_fsm counter_module_run_run_fsm_inst (
      .clk(clk),
      .rst(rst),
      .counter_out_Push_mioi_wen_comp(counter_out_Push_mioi_wen_comp),
      .fsm_output(fsm_output)
    );
  assign and_rmff = (fsm_output==2'b01);
  assign nl_while_ac_int_cctor_sva_1 = counter_out_sig_sva + 32'b00000000000000000000000000000001;
  assign while_ac_int_cctor_sva_1 = nl_while_ac_int_cctor_sva_1[31:0];
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_counter_out_Push_mioi_iswt0_cse <= 1'b0;
    end
    else if ( counter_out_Push_mioi_wen_comp ) begin
      reg_counter_out_Push_mioi_iswt0_cse <= and_rmff;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      counter_out_sig_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( counter_out_Push_mioi_wen_comp & (~((fsm_output!=2'b01))) ) begin
      counter_out_sig_sva <= while_ac_int_cctor_sva_1;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    counter_top_add_run
// ------------------------------------------------------------------


module counter_top_add_run (
  clk, rst, counter_in_vld, counter_in_rdy, counter_in_dat, add_out_vld, add_out_rdy,
      add_out_dat
);
  input clk;
  input rst;
  input counter_in_vld;
  output counter_in_rdy;
  input [31:0] counter_in_dat;
  output add_out_vld;
  input add_out_rdy;
  output [31:0] add_out_dat;


  // Interconnect Declarations
  wire run_wen;
  wire counter_in_Pop_mioi_wen_comp;
  wire [31:0] counter_in_Pop_mioi_return_rsc_z_mxwt;
  wire add_out_Push_mioi_wen_comp;
  wire [1:0] fsm_output;
  reg reg_add_out_Push_mioi_iswt0_cse;
  reg reg_counter_in_Pop_mioi_iswt0_cse;
  wire and_1_rmff;
  wire and_rmff;


  // Interconnect Declarations for Component Instantiations 
  wire  nl_add_run_counter_in_Pop_mioi_inst_run_wten;
  assign nl_add_run_counter_in_Pop_mioi_inst_run_wten = ~ run_wen;
  wire  nl_add_run_add_out_Push_mioi_inst_run_wten;
  assign nl_add_run_add_out_Push_mioi_inst_run_wten = ~ run_wen;
  wire [32:0] nl_add_run_add_out_Push_mioi_inst_add_out_Push_mioi_m_rsc_dat_run;
  assign nl_add_run_add_out_Push_mioi_inst_add_out_Push_mioi_m_rsc_dat_run = counter_in_Pop_mioi_return_rsc_z_mxwt
      + 32'b00000000000000000000000000000101;
  counter_top_add_run_counter_in_Pop_mioi add_run_counter_in_Pop_mioi_inst (
      .clk(clk),
      .rst(rst),
      .counter_in_vld(counter_in_vld),
      .counter_in_rdy(counter_in_rdy),
      .counter_in_dat(counter_in_dat),
      .run_wten(nl_add_run_counter_in_Pop_mioi_inst_run_wten),
      .counter_in_Pop_mioi_oswt(reg_counter_in_Pop_mioi_iswt0_cse),
      .counter_in_Pop_mioi_wen_comp(counter_in_Pop_mioi_wen_comp),
      .counter_in_Pop_mioi_return_rsc_z_mxwt(counter_in_Pop_mioi_return_rsc_z_mxwt),
      .counter_in_Pop_mioi_oswt_pff(and_1_rmff)
    );
  counter_top_add_run_add_out_Push_mioi add_run_add_out_Push_mioi_inst (
      .clk(clk),
      .rst(rst),
      .add_out_vld(add_out_vld),
      .add_out_rdy(add_out_rdy),
      .add_out_dat(add_out_dat),
      .run_wten(nl_add_run_add_out_Push_mioi_inst_run_wten),
      .add_out_Push_mioi_oswt(reg_add_out_Push_mioi_iswt0_cse),
      .add_out_Push_mioi_wen_comp(add_out_Push_mioi_wen_comp),
      .add_out_Push_mioi_m_rsc_dat_run(nl_add_run_add_out_Push_mioi_inst_add_out_Push_mioi_m_rsc_dat_run[31:0]),
      .add_out_Push_mioi_oswt_pff(and_rmff)
    );
  counter_top_add_run_staller add_run_staller_inst (
      .run_wen(run_wen),
      .counter_in_Pop_mioi_wen_comp(counter_in_Pop_mioi_wen_comp),
      .add_out_Push_mioi_wen_comp(add_out_Push_mioi_wen_comp)
    );
  counter_top_add_run_run_fsm add_run_run_fsm_inst (
      .clk(clk),
      .rst(rst),
      .run_wen(run_wen),
      .fsm_output(fsm_output)
    );
  assign and_rmff = (fsm_output==2'b10);
  assign and_1_rmff = (fsm_output==2'b01);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_add_out_Push_mioi_iswt0_cse <= 1'b0;
      reg_counter_in_Pop_mioi_iswt0_cse <= 1'b0;
    end
    else if ( run_wen ) begin
      reg_add_out_Push_mioi_iswt0_cse <= and_rmff;
      reg_counter_in_Pop_mioi_iswt0_cse <= and_1_rmff;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    counter_top_counter_module
// ------------------------------------------------------------------


module counter_top_counter_module (
  clk, rst, counter_out_vld, counter_out_rdy, counter_out_dat
);
  input clk;
  input rst;
  output counter_out_vld;
  input counter_out_rdy;
  output [31:0] counter_out_dat;



  // Interconnect Declarations for Component Instantiations 
  counter_top_counter_module_run counter_module_run_inst (
      .clk(clk),
      .rst(rst),
      .counter_out_vld(counter_out_vld),
      .counter_out_rdy(counter_out_rdy),
      .counter_out_dat(counter_out_dat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    counter_top_add
// ------------------------------------------------------------------


module counter_top_add (
  clk, rst, counter_in_vld, counter_in_rdy, counter_in_dat, add_out_vld, add_out_rdy,
      add_out_dat
);
  input clk;
  input rst;
  input counter_in_vld;
  output counter_in_rdy;
  input [31:0] counter_in_dat;
  output add_out_vld;
  input add_out_rdy;
  output [31:0] add_out_dat;



  // Interconnect Declarations for Component Instantiations 
  counter_top_add_run add_run_inst (
      .clk(clk),
      .rst(rst),
      .counter_in_vld(counter_in_vld),
      .counter_in_rdy(counter_in_rdy),
      .counter_in_dat(counter_in_dat),
      .add_out_vld(add_out_vld),
      .add_out_rdy(add_out_rdy),
      .add_out_dat(add_out_dat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    counter_top
// ------------------------------------------------------------------


module counter_top (
  clk, rst, counter_out, add_out
);
  input clk;
  input rst;
  output [31:0] counter_out;
  output [31:0] add_out;


  // Interconnect Declarations
  wire counter_module_out_vld;
  wire counter_module_out_rdy;
  wire [31:0] counter_module_out_dat;
  wire counter_in_vld;
  wire counter_in_rdy;
  wire [31:0] counter_in_dat;
  wire add_to_top_vld;
  wire add_to_top_rdy;
  wire [31:0] add_to_top_dat;


  // Interconnect Declarations for Component Instantiations 
  counter_top_counter_module counter_inst (
      .clk(clk),
      .rst(rst),
      .counter_out_vld(counter_module_out_vld),
      .counter_out_rdy(counter_module_out_rdy),
      .counter_out_dat(counter_module_out_dat)
    );
  counter_top_add add_inst (
      .clk(clk),
      .rst(rst),
      .counter_in_vld(counter_in_vld),
      .counter_in_rdy(counter_in_rdy),
      .counter_in_dat(counter_in_dat),
      .add_out_vld(add_to_top_vld),
      .add_out_rdy(add_to_top_rdy),
      .add_out_dat(add_to_top_dat)
    );
  counter_top_counter_top_run counter_top_run_inst (
      .clk(clk),
      .rst(rst),
      .counter_out(counter_out),
      .add_out(add_out),
      .counter_module_out_vld(counter_module_out_vld),
      .counter_module_out_rdy(counter_module_out_rdy),
      .counter_module_out_dat(counter_module_out_dat),
      .counter_in_vld(counter_in_vld),
      .counter_in_rdy(counter_in_rdy),
      .counter_in_dat(counter_in_dat),
      .add_to_top_vld(add_to_top_vld),
      .add_to_top_rdy(add_to_top_rdy),
      .add_to_top_dat(add_to_top_dat)
    );
endmodule



